module tt_um_flummer_ltc (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire \ltc.bit_clk ;
 wire \ltc.bit_counter[0] ;
 wire \ltc.bit_counter[10] ;
 wire \ltc.bit_counter[11] ;
 wire \ltc.bit_counter[1] ;
 wire \ltc.bit_counter[2] ;
 wire \ltc.bit_counter[3] ;
 wire \ltc.bit_counter[4] ;
 wire \ltc.bit_counter[5] ;
 wire \ltc.bit_counter[6] ;
 wire \ltc.bit_counter[7] ;
 wire \ltc.bit_counter[8] ;
 wire \ltc.bit_counter[9] ;
 wire \ltc.frm_counter[0] ;
 wire \ltc.frm_counter[10] ;
 wire \ltc.frm_counter[11] ;
 wire \ltc.frm_counter[12] ;
 wire \ltc.frm_counter[13] ;
 wire \ltc.frm_counter[14] ;
 wire \ltc.frm_counter[15] ;
 wire \ltc.frm_counter[16] ;
 wire \ltc.frm_counter[17] ;
 wire \ltc.frm_counter[18] ;
 wire \ltc.frm_counter[19] ;
 wire \ltc.frm_counter[1] ;
 wire \ltc.frm_counter[20] ;
 wire \ltc.frm_counter[21] ;
 wire \ltc.frm_counter[22] ;
 wire \ltc.frm_counter[23] ;
 wire \ltc.frm_counter[2] ;
 wire \ltc.frm_counter[3] ;
 wire \ltc.frm_counter[4] ;
 wire \ltc.frm_counter[5] ;
 wire \ltc.frm_counter[6] ;
 wire \ltc.frm_counter[7] ;
 wire \ltc.frm_counter[8] ;
 wire \ltc.frm_counter[9] ;
 wire \ltc.frm_d[0] ;
 wire \ltc.frm_d[1] ;
 wire \ltc.frm_u[0] ;
 wire \ltc.frm_u[1] ;
 wire \ltc.frm_u[2] ;
 wire \ltc.frm_u[3] ;
 wire \ltc.hrs_d[0] ;
 wire \ltc.hrs_d[1] ;
 wire \ltc.hrs_u[0] ;
 wire \ltc.hrs_u[1] ;
 wire \ltc.hrs_u[2] ;
 wire \ltc.hrs_u[3] ;
 wire \ltc.min_d[0] ;
 wire \ltc.min_d[1] ;
 wire \ltc.min_d[2] ;
 wire \ltc.min_u[0] ;
 wire \ltc.min_u[1] ;
 wire \ltc.min_u[2] ;
 wire \ltc.min_u[3] ;
 wire \ltc.output_buffer[0] ;
 wire \ltc.output_buffer[10] ;
 wire \ltc.output_buffer[11] ;
 wire \ltc.output_buffer[12] ;
 wire \ltc.output_buffer[13] ;
 wire \ltc.output_buffer[14] ;
 wire \ltc.output_buffer[15] ;
 wire \ltc.output_buffer[16] ;
 wire \ltc.output_buffer[17] ;
 wire \ltc.output_buffer[18] ;
 wire \ltc.output_buffer[19] ;
 wire \ltc.output_buffer[1] ;
 wire \ltc.output_buffer[20] ;
 wire \ltc.output_buffer[21] ;
 wire \ltc.output_buffer[22] ;
 wire \ltc.output_buffer[23] ;
 wire \ltc.output_buffer[24] ;
 wire \ltc.output_buffer[25] ;
 wire \ltc.output_buffer[26] ;
 wire \ltc.output_buffer[27] ;
 wire \ltc.output_buffer[28] ;
 wire \ltc.output_buffer[29] ;
 wire \ltc.output_buffer[2] ;
 wire \ltc.output_buffer[30] ;
 wire \ltc.output_buffer[31] ;
 wire \ltc.output_buffer[32] ;
 wire \ltc.output_buffer[33] ;
 wire \ltc.output_buffer[34] ;
 wire \ltc.output_buffer[35] ;
 wire \ltc.output_buffer[36] ;
 wire \ltc.output_buffer[37] ;
 wire \ltc.output_buffer[38] ;
 wire \ltc.output_buffer[39] ;
 wire \ltc.output_buffer[3] ;
 wire \ltc.output_buffer[40] ;
 wire \ltc.output_buffer[41] ;
 wire \ltc.output_buffer[42] ;
 wire \ltc.output_buffer[43] ;
 wire \ltc.output_buffer[44] ;
 wire \ltc.output_buffer[45] ;
 wire \ltc.output_buffer[46] ;
 wire \ltc.output_buffer[47] ;
 wire \ltc.output_buffer[48] ;
 wire \ltc.output_buffer[49] ;
 wire \ltc.output_buffer[4] ;
 wire \ltc.output_buffer[50] ;
 wire \ltc.output_buffer[51] ;
 wire \ltc.output_buffer[52] ;
 wire \ltc.output_buffer[53] ;
 wire \ltc.output_buffer[54] ;
 wire \ltc.output_buffer[55] ;
 wire \ltc.output_buffer[56] ;
 wire \ltc.output_buffer[57] ;
 wire \ltc.output_buffer[58] ;
 wire \ltc.output_buffer[59] ;
 wire \ltc.output_buffer[5] ;
 wire \ltc.output_buffer[60] ;
 wire \ltc.output_buffer[61] ;
 wire \ltc.output_buffer[62] ;
 wire \ltc.output_buffer[63] ;
 wire \ltc.output_buffer[64] ;
 wire \ltc.output_buffer[65] ;
 wire \ltc.output_buffer[66] ;
 wire \ltc.output_buffer[67] ;
 wire \ltc.output_buffer[68] ;
 wire \ltc.output_buffer[69] ;
 wire \ltc.output_buffer[6] ;
 wire \ltc.output_buffer[70] ;
 wire \ltc.output_buffer[71] ;
 wire \ltc.output_buffer[72] ;
 wire \ltc.output_buffer[73] ;
 wire \ltc.output_buffer[74] ;
 wire \ltc.output_buffer[75] ;
 wire \ltc.output_buffer[76] ;
 wire \ltc.output_buffer[77] ;
 wire \ltc.output_buffer[78] ;
 wire \ltc.output_buffer[79] ;
 wire \ltc.output_buffer[7] ;
 wire \ltc.output_buffer[8] ;
 wire \ltc.output_buffer[9] ;
 wire \ltc.sec_d[0] ;
 wire \ltc.sec_d[1] ;
 wire \ltc.sec_d[2] ;
 wire \ltc.sec_u[0] ;
 wire \ltc.sec_u[1] ;
 wire \ltc.sec_u[2] ;
 wire \ltc.sec_u[3] ;
 wire \ltc.timecode ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;

 sg13g2_inv_1 _0714_ (.Y(_0144_),
    .A(net445));
 sg13g2_inv_1 _0715_ (.Y(_0145_),
    .A(net413));
 sg13g2_inv_1 _0716_ (.Y(_0146_),
    .A(\ltc.frm_u[0] ));
 sg13g2_inv_1 _0717_ (.Y(_0147_),
    .A(net469));
 sg13g2_inv_1 _0718_ (.Y(_0148_),
    .A(net464));
 sg13g2_inv_1 _0719_ (.Y(_0149_),
    .A(net452));
 sg13g2_inv_1 _0720_ (.Y(_0150_),
    .A(net409));
 sg13g2_inv_1 _0721_ (.Y(_0151_),
    .A(net426));
 sg13g2_inv_1 _0722_ (.Y(_0152_),
    .A(\ltc.frm_counter[12] ));
 sg13g2_inv_1 _0723_ (.Y(_0153_),
    .A(net473));
 sg13g2_inv_1 _0724_ (.Y(_0154_),
    .A(\ltc.bit_counter[6] ));
 sg13g2_inv_1 _0725_ (.Y(_0155_),
    .A(net177));
 sg13g2_inv_1 _0726_ (.Y(_0156_),
    .A(net251));
 sg13g2_inv_1 _0727_ (.Y(_0157_),
    .A(net260));
 sg13g2_inv_1 _0728_ (.Y(_0158_),
    .A(net264));
 sg13g2_inv_1 _0729_ (.Y(_0159_),
    .A(net247));
 sg13g2_inv_1 _0730_ (.Y(_0160_),
    .A(net250));
 sg13g2_inv_1 _0731_ (.Y(_0161_),
    .A(net233));
 sg13g2_inv_1 _0732_ (.Y(_0162_),
    .A(net242));
 sg13g2_inv_1 _0733_ (.Y(_0163_),
    .A(net237));
 sg13g2_inv_1 _0734_ (.Y(_0164_),
    .A(net255));
 sg13g2_inv_1 _0735_ (.Y(_0165_),
    .A(net245));
 sg13g2_inv_1 _0736_ (.Y(_0166_),
    .A(net243));
 sg13g2_inv_1 _0737_ (.Y(_0167_),
    .A(net256));
 sg13g2_inv_1 _0738_ (.Y(_0168_),
    .A(net253));
 sg13g2_nand2_1 _0739_ (.Y(_0169_),
    .A(net7),
    .B(net8));
 sg13g2_nand4_1 _0740_ (.B(net5),
    .C(net2),
    .A(net6),
    .Y(_0170_),
    .D(net1));
 sg13g2_nor2_1 _0741_ (.A(_0169_),
    .B(_0170_),
    .Y(uo_out[0]));
 sg13g2_nor2_1 _0742_ (.A(net361),
    .B(net227),
    .Y(_0171_));
 sg13g2_nor3_1 _0743_ (.A(\ltc.bit_counter[2] ),
    .B(\ltc.bit_counter[10] ),
    .C(\ltc.bit_counter[11] ),
    .Y(_0172_));
 sg13g2_nor2_1 _0744_ (.A(\ltc.bit_counter[5] ),
    .B(\ltc.bit_counter[4] ),
    .Y(_0173_));
 sg13g2_nor2_1 _0745_ (.A(\ltc.bit_counter[8] ),
    .B(\ltc.bit_counter[9] ),
    .Y(_0174_));
 sg13g2_nor4_1 _0746_ (.A(\ltc.bit_counter[1] ),
    .B(net227),
    .C(\ltc.bit_counter[6] ),
    .D(\ltc.bit_counter[7] ),
    .Y(_0175_));
 sg13g2_nor3_1 _0747_ (.A(\ltc.bit_counter[5] ),
    .B(\ltc.bit_counter[4] ),
    .C(\ltc.bit_counter[3] ),
    .Y(_0176_));
 sg13g2_nand4_1 _0748_ (.B(_0174_),
    .C(_0175_),
    .A(_0172_),
    .Y(_0177_),
    .D(_0176_));
 sg13g2_nor2_1 _0749_ (.A(net231),
    .B(_0177_),
    .Y(_0178_));
 sg13g2_nor2_2 _0750_ (.A(net173),
    .B(net163),
    .Y(_0179_));
 sg13g2_nor3_1 _0751_ (.A(\ltc.frm_counter[16] ),
    .B(\ltc.frm_counter[17] ),
    .C(\ltc.frm_counter[18] ),
    .Y(_0180_));
 sg13g2_nor4_1 _0752_ (.A(\ltc.frm_counter[10] ),
    .B(\ltc.frm_counter[11] ),
    .C(\ltc.frm_counter[12] ),
    .D(\ltc.frm_counter[13] ),
    .Y(_0181_));
 sg13g2_nor4_1 _0753_ (.A(\ltc.frm_counter[3] ),
    .B(\ltc.frm_counter[2] ),
    .C(\ltc.frm_counter[6] ),
    .D(\ltc.frm_counter[7] ),
    .Y(_0182_));
 sg13g2_nand3_1 _0754_ (.B(_0181_),
    .C(_0182_),
    .A(_0180_),
    .Y(_0183_));
 sg13g2_nor2_1 _0755_ (.A(\ltc.frm_counter[19] ),
    .B(\ltc.frm_counter[20] ),
    .Y(_0184_));
 sg13g2_nor3_1 _0756_ (.A(\ltc.frm_counter[21] ),
    .B(\ltc.frm_counter[22] ),
    .C(\ltc.frm_counter[23] ),
    .Y(_0185_));
 sg13g2_nand2_1 _0757_ (.Y(_0186_),
    .A(_0184_),
    .B(_0185_));
 sg13g2_nor2_1 _0758_ (.A(\ltc.frm_counter[14] ),
    .B(\ltc.frm_counter[15] ),
    .Y(_0187_));
 sg13g2_nor2_1 _0759_ (.A(net466),
    .B(net463),
    .Y(_0188_));
 sg13g2_nor2_1 _0760_ (.A(\ltc.frm_counter[5] ),
    .B(\ltc.frm_counter[4] ),
    .Y(_0189_));
 sg13g2_nand3_1 _0761_ (.B(_0188_),
    .C(_0189_),
    .A(_0187_),
    .Y(_0190_));
 sg13g2_nor3_2 _0762_ (.A(_0183_),
    .B(_0186_),
    .C(_0190_),
    .Y(_0191_));
 sg13g2_nor2b_2 _0763_ (.A(net450),
    .B_N(net230),
    .Y(_0192_));
 sg13g2_and2_1 _0764_ (.A(_0191_),
    .B(_0192_),
    .X(_0193_));
 sg13g2_nand2_2 _0765_ (.Y(_0194_),
    .A(_0191_),
    .B(_0192_));
 sg13g2_o21ai_1 _0766_ (.B1(net147),
    .Y(_0195_),
    .A1(net415),
    .A2(net142));
 sg13g2_inv_1 _0767_ (.Y(_0000_),
    .A(_0195_));
 sg13g2_nor2_1 _0768_ (.A(net155),
    .B(net143),
    .Y(_0196_));
 sg13g2_a22oi_1 _0769_ (.Y(_0197_),
    .B1(net132),
    .B2(net251),
    .A2(net155),
    .A1(\ltc.output_buffer[0] ));
 sg13g2_nor2_1 _0770_ (.A(net169),
    .B(net252),
    .Y(_0001_));
 sg13g2_a221oi_1 _0771_ (.B2(_0157_),
    .C1(net169),
    .B1(net133),
    .A1(_0156_),
    .Y(_0002_),
    .A2(net155));
 sg13g2_a221oi_1 _0772_ (.B2(_0158_),
    .C1(net169),
    .B1(net133),
    .A1(_0157_),
    .Y(_0003_),
    .A2(net157));
 sg13g2_a221oi_1 _0773_ (.B2(_0159_),
    .C1(net169),
    .B1(net133),
    .A1(_0158_),
    .Y(_0004_),
    .A2(net155));
 sg13g2_a221oi_1 _0774_ (.B2(_0160_),
    .C1(net167),
    .B1(net133),
    .A1(_0159_),
    .Y(_0005_),
    .A2(net155));
 sg13g2_a221oi_1 _0775_ (.B2(_0161_),
    .C1(net167),
    .B1(net132),
    .A1(_0160_),
    .Y(_0006_),
    .A2(net154));
 sg13g2_a221oi_1 _0776_ (.B2(_0162_),
    .C1(net167),
    .B1(net131),
    .A1(_0161_),
    .Y(_0007_),
    .A2(net154));
 sg13g2_a221oi_1 _0777_ (.B2(_0163_),
    .C1(net166),
    .B1(net131),
    .A1(_0162_),
    .Y(_0008_),
    .A2(net152));
 sg13g2_a221oi_1 _0778_ (.B2(_0164_),
    .C1(net166),
    .B1(net131),
    .A1(_0163_),
    .Y(_0009_),
    .A2(net153));
 sg13g2_a221oi_1 _0779_ (.B2(_0165_),
    .C1(net166),
    .B1(net132),
    .A1(_0164_),
    .Y(_0010_),
    .A2(net152));
 sg13g2_a221oi_1 _0780_ (.B2(_0166_),
    .C1(net167),
    .B1(net132),
    .A1(_0165_),
    .Y(_0011_),
    .A2(net152));
 sg13g2_a221oi_1 _0781_ (.B2(_0167_),
    .C1(net166),
    .B1(net131),
    .A1(_0166_),
    .Y(_0012_),
    .A2(net152));
 sg13g2_a221oi_1 _0782_ (.B2(_0168_),
    .C1(net166),
    .B1(net132),
    .A1(_0167_),
    .Y(_0013_),
    .A2(net152));
 sg13g2_a22oi_1 _0783_ (.Y(_0198_),
    .B1(net131),
    .B2(net235),
    .A2(net152),
    .A1(\ltc.output_buffer[13] ));
 sg13g2_nor2_1 _0784_ (.A(net166),
    .B(net236),
    .Y(_0014_));
 sg13g2_a22oi_1 _0785_ (.Y(_0199_),
    .B1(net131),
    .B2(net249),
    .A2(net152),
    .A1(net235));
 sg13g2_nor2_1 _0786_ (.A(net166),
    .B(_0199_),
    .Y(_0015_));
 sg13g2_a22oi_1 _0787_ (.Y(_0200_),
    .B1(net131),
    .B2(net288),
    .A2(net152),
    .A1(net249));
 sg13g2_nor2_1 _0788_ (.A(net166),
    .B(_0200_),
    .Y(_0016_));
 sg13g2_a22oi_1 _0789_ (.Y(_0201_),
    .B1(net131),
    .B2(net360),
    .A2(net154),
    .A1(net288));
 sg13g2_nor2_1 _0790_ (.A(net167),
    .B(_0201_),
    .Y(_0017_));
 sg13g2_a22oi_1 _0791_ (.Y(_0202_),
    .B1(net132),
    .B2(net326),
    .A2(net154),
    .A1(\ltc.output_buffer[17] ));
 sg13g2_nor2_1 _0792_ (.A(net167),
    .B(net327),
    .Y(_0018_));
 sg13g2_a22oi_1 _0793_ (.Y(_0203_),
    .B1(net132),
    .B2(net282),
    .A2(net155),
    .A1(net326));
 sg13g2_nor2_1 _0794_ (.A(net169),
    .B(_0203_),
    .Y(_0019_));
 sg13g2_nand2_1 _0795_ (.Y(_0204_),
    .A(net282),
    .B(net155));
 sg13g2_nor2b_1 _0796_ (.A(net230),
    .B_N(net450),
    .Y(_0205_));
 sg13g2_and2_1 _0797_ (.A(_0191_),
    .B(_0205_),
    .X(_0206_));
 sg13g2_nor2b_2 _0798_ (.A(net4),
    .B_N(net3),
    .Y(_0207_));
 sg13g2_nand2_2 _0799_ (.Y(_0208_),
    .A(_0206_),
    .B(_0207_));
 sg13g2_xor2_1 _0800_ (.B(\ltc.output_buffer[66] ),
    .A(\ltc.output_buffer[67] ),
    .X(_0209_));
 sg13g2_xor2_1 _0801_ (.B(\ltc.output_buffer[64] ),
    .A(\ltc.output_buffer[65] ),
    .X(_0210_));
 sg13g2_xnor2_1 _0802_ (.Y(_0211_),
    .A(_0209_),
    .B(_0210_));
 sg13g2_xnor2_1 _0803_ (.Y(_0212_),
    .A(\ltc.output_buffer[71] ),
    .B(\ltc.output_buffer[70] ));
 sg13g2_xor2_1 _0804_ (.B(\ltc.output_buffer[68] ),
    .A(\ltc.output_buffer[69] ),
    .X(_0213_));
 sg13g2_xnor2_1 _0805_ (.Y(_0214_),
    .A(_0212_),
    .B(_0213_));
 sg13g2_xnor2_1 _0806_ (.Y(_0215_),
    .A(_0211_),
    .B(_0214_));
 sg13g2_xnor2_1 _0807_ (.Y(_0216_),
    .A(\ltc.output_buffer[51] ),
    .B(\ltc.output_buffer[50] ));
 sg13g2_xor2_1 _0808_ (.B(\ltc.output_buffer[48] ),
    .A(\ltc.output_buffer[49] ),
    .X(_0217_));
 sg13g2_xnor2_1 _0809_ (.Y(_0218_),
    .A(_0216_),
    .B(_0217_));
 sg13g2_xnor2_1 _0810_ (.Y(_0219_),
    .A(\ltc.output_buffer[55] ),
    .B(\ltc.output_buffer[54] ));
 sg13g2_xor2_1 _0811_ (.B(\ltc.output_buffer[53] ),
    .A(\ltc.output_buffer[52] ),
    .X(_0220_));
 sg13g2_xnor2_1 _0812_ (.Y(_0221_),
    .A(_0219_),
    .B(_0220_));
 sg13g2_xnor2_1 _0813_ (.Y(_0222_),
    .A(_0218_),
    .B(_0221_));
 sg13g2_xnor2_1 _0814_ (.Y(_0223_),
    .A(_0215_),
    .B(_0222_));
 sg13g2_xnor2_1 _0815_ (.Y(_0224_),
    .A(\ltc.output_buffer[63] ),
    .B(\ltc.output_buffer[62] ));
 sg13g2_xor2_1 _0816_ (.B(\ltc.output_buffer[60] ),
    .A(\ltc.output_buffer[61] ),
    .X(_0225_));
 sg13g2_xnor2_1 _0817_ (.Y(_0226_),
    .A(_0224_),
    .B(_0225_));
 sg13g2_xnor2_1 _0818_ (.Y(_0227_),
    .A(\ltc.output_buffer[76] ),
    .B(\ltc.output_buffer[78] ));
 sg13g2_xor2_1 _0819_ (.B(\ltc.output_buffer[77] ),
    .A(\ltc.output_buffer[79] ),
    .X(_0228_));
 sg13g2_xnor2_1 _0820_ (.Y(_0229_),
    .A(_0227_),
    .B(_0228_));
 sg13g2_xnor2_1 _0821_ (.Y(_0230_),
    .A(_0226_),
    .B(_0229_));
 sg13g2_xnor2_1 _0822_ (.Y(_0231_),
    .A(\ltc.output_buffer[59] ),
    .B(\ltc.output_buffer[58] ));
 sg13g2_xnor2_1 _0823_ (.Y(_0232_),
    .A(\ltc.output_buffer[73] ),
    .B(\ltc.output_buffer[72] ));
 sg13g2_xnor2_1 _0824_ (.Y(_0233_),
    .A(_0231_),
    .B(_0232_));
 sg13g2_xor2_1 _0825_ (.B(\ltc.output_buffer[56] ),
    .A(\ltc.output_buffer[57] ),
    .X(_0234_));
 sg13g2_xnor2_1 _0826_ (.Y(_0235_),
    .A(\ltc.output_buffer[75] ),
    .B(\ltc.output_buffer[74] ));
 sg13g2_xnor2_1 _0827_ (.Y(_0236_),
    .A(_0234_),
    .B(_0235_));
 sg13g2_xnor2_1 _0828_ (.Y(_0237_),
    .A(_0233_),
    .B(_0236_));
 sg13g2_xnor2_1 _0829_ (.Y(_0238_),
    .A(_0230_),
    .B(_0237_));
 sg13g2_xnor2_1 _0830_ (.Y(_0239_),
    .A(_0223_),
    .B(_0238_));
 sg13g2_xnor2_1 _0831_ (.Y(_0240_),
    .A(\ltc.output_buffer[19] ),
    .B(\ltc.output_buffer[18] ));
 sg13g2_xor2_1 _0832_ (.B(\ltc.output_buffer[16] ),
    .A(\ltc.output_buffer[17] ),
    .X(_0241_));
 sg13g2_xnor2_1 _0833_ (.Y(_0242_),
    .A(_0240_),
    .B(_0241_));
 sg13g2_xnor2_1 _0834_ (.Y(_0243_),
    .A(\ltc.output_buffer[23] ),
    .B(\ltc.output_buffer[22] ));
 sg13g2_xor2_1 _0835_ (.B(\ltc.output_buffer[20] ),
    .A(\ltc.output_buffer[21] ),
    .X(_0244_));
 sg13g2_xnor2_1 _0836_ (.Y(_0245_),
    .A(_0243_),
    .B(_0244_));
 sg13g2_xnor2_1 _0837_ (.Y(_0246_),
    .A(_0242_),
    .B(_0245_));
 sg13g2_xor2_1 _0838_ (.B(\ltc.output_buffer[34] ),
    .A(\ltc.output_buffer[35] ),
    .X(_0247_));
 sg13g2_xnor2_1 _0839_ (.Y(_0248_),
    .A(\ltc.output_buffer[37] ),
    .B(\ltc.output_buffer[36] ));
 sg13g2_xnor2_1 _0840_ (.Y(_0249_),
    .A(_0247_),
    .B(_0248_));
 sg13g2_xor2_1 _0841_ (.B(\ltc.output_buffer[32] ),
    .A(\ltc.output_buffer[33] ),
    .X(_0250_));
 sg13g2_xnor2_1 _0842_ (.Y(_0251_),
    .A(\ltc.output_buffer[39] ),
    .B(\ltc.output_buffer[38] ));
 sg13g2_xnor2_1 _0843_ (.Y(_0252_),
    .A(_0250_),
    .B(_0251_));
 sg13g2_xnor2_1 _0844_ (.Y(_0253_),
    .A(_0249_),
    .B(_0252_));
 sg13g2_xnor2_1 _0845_ (.Y(_0254_),
    .A(_0246_),
    .B(_0253_));
 sg13g2_xor2_1 _0846_ (.B(\ltc.output_buffer[30] ),
    .A(\ltc.output_buffer[31] ),
    .X(_0255_));
 sg13g2_xor2_1 _0847_ (.B(\ltc.output_buffer[28] ),
    .A(\ltc.output_buffer[29] ),
    .X(_0256_));
 sg13g2_xnor2_1 _0848_ (.Y(_0257_),
    .A(_0255_),
    .B(_0256_));
 sg13g2_xnor2_1 _0849_ (.Y(_0258_),
    .A(\ltc.output_buffer[47] ),
    .B(\ltc.output_buffer[46] ));
 sg13g2_xor2_1 _0850_ (.B(\ltc.output_buffer[44] ),
    .A(\ltc.output_buffer[45] ),
    .X(_0259_));
 sg13g2_xnor2_1 _0851_ (.Y(_0260_),
    .A(_0258_),
    .B(_0259_));
 sg13g2_xnor2_1 _0852_ (.Y(_0261_),
    .A(_0257_),
    .B(_0260_));
 sg13g2_xnor2_1 _0853_ (.Y(_0262_),
    .A(\ltc.output_buffer[27] ),
    .B(\ltc.output_buffer[26] ));
 sg13g2_xnor2_1 _0854_ (.Y(_0263_),
    .A(\ltc.output_buffer[41] ),
    .B(\ltc.output_buffer[40] ));
 sg13g2_xnor2_1 _0855_ (.Y(_0264_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_xor2_1 _0856_ (.B(\ltc.output_buffer[24] ),
    .A(\ltc.output_buffer[25] ),
    .X(_0265_));
 sg13g2_xnor2_1 _0857_ (.Y(_0266_),
    .A(\ltc.output_buffer[43] ),
    .B(\ltc.output_buffer[42] ));
 sg13g2_xnor2_1 _0858_ (.Y(_0267_),
    .A(_0265_),
    .B(_0266_));
 sg13g2_xnor2_1 _0859_ (.Y(_0268_),
    .A(_0264_),
    .B(_0267_));
 sg13g2_xnor2_1 _0860_ (.Y(_0269_),
    .A(_0261_),
    .B(_0268_));
 sg13g2_xnor2_1 _0861_ (.Y(_0270_),
    .A(_0254_),
    .B(_0269_));
 sg13g2_xnor2_1 _0862_ (.Y(_0271_),
    .A(_0239_),
    .B(_0270_));
 sg13g2_nand2_1 _0863_ (.Y(_0272_),
    .A(\ltc.output_buffer[20] ),
    .B(net139));
 sg13g2_a21oi_1 _0864_ (.A1(_0208_),
    .A2(_0272_),
    .Y(_0273_),
    .B1(net156));
 sg13g2_o21ai_1 _0865_ (.B1(_0273_),
    .Y(_0274_),
    .A1(_0208_),
    .A2(_0271_));
 sg13g2_a21oi_1 _0866_ (.A1(_0204_),
    .A2(_0274_),
    .Y(_0020_),
    .B1(net169));
 sg13g2_a22oi_1 _0867_ (.Y(_0275_),
    .B1(net134),
    .B2(net368),
    .A2(net155),
    .A1(\ltc.output_buffer[20] ));
 sg13g2_nor2_1 _0868_ (.A(net170),
    .B(net369),
    .Y(_0021_));
 sg13g2_nand3_1 _0869_ (.B(net368),
    .C(net156),
    .A(net177),
    .Y(_0276_));
 sg13g2_nor2_1 _0870_ (.A(net409),
    .B(net138),
    .Y(_0277_));
 sg13g2_o21ai_1 _0871_ (.B1(net146),
    .Y(_0278_),
    .A1(net295),
    .A2(net143));
 sg13g2_o21ai_1 _0872_ (.B1(_0276_),
    .Y(_0022_),
    .A1(_0277_),
    .A2(_0278_));
 sg13g2_nor2_1 _0873_ (.A(\ltc.hrs_d[0] ),
    .B(net139),
    .Y(_0279_));
 sg13g2_o21ai_1 _0874_ (.B1(net147),
    .Y(_0280_),
    .A1(\ltc.output_buffer[23] ),
    .A2(net143));
 sg13g2_nand3_1 _0875_ (.B(net295),
    .C(net150),
    .A(net176),
    .Y(_0281_));
 sg13g2_o21ai_1 _0876_ (.B1(_0281_),
    .Y(_0023_),
    .A1(_0279_),
    .A2(_0280_));
 sg13g2_a22oi_1 _0877_ (.Y(_0282_),
    .B1(net129),
    .B2(net353),
    .A2(net154),
    .A1(\ltc.output_buffer[23] ));
 sg13g2_nor2_1 _0878_ (.A(net168),
    .B(net354),
    .Y(_0024_));
 sg13g2_a22oi_1 _0879_ (.Y(_0283_),
    .B1(net130),
    .B2(net371),
    .A2(net153),
    .A1(net353));
 sg13g2_nor2_1 _0880_ (.A(net165),
    .B(_0283_),
    .Y(_0025_));
 sg13g2_a22oi_1 _0881_ (.Y(_0284_),
    .B1(net130),
    .B2(net309),
    .A2(net153),
    .A1(\ltc.output_buffer[25] ));
 sg13g2_nor2_1 _0882_ (.A(net165),
    .B(net310),
    .Y(_0026_));
 sg13g2_a22oi_1 _0883_ (.Y(_0285_),
    .B1(net129),
    .B2(net289),
    .A2(net150),
    .A1(net309));
 sg13g2_nor2_1 _0884_ (.A(net165),
    .B(_0285_),
    .Y(_0027_));
 sg13g2_nand3_1 _0885_ (.B(net289),
    .C(net151),
    .A(net176),
    .Y(_0286_));
 sg13g2_nor2_1 _0886_ (.A(\ltc.hrs_u[3] ),
    .B(net138),
    .Y(_0287_));
 sg13g2_o21ai_1 _0887_ (.B1(net146),
    .Y(_0288_),
    .A1(\ltc.output_buffer[28] ),
    .A2(net142));
 sg13g2_o21ai_1 _0888_ (.B1(_0286_),
    .Y(_0028_),
    .A1(_0287_),
    .A2(_0288_));
 sg13g2_nor2_1 _0889_ (.A(\ltc.hrs_u[2] ),
    .B(net138),
    .Y(_0289_));
 sg13g2_o21ai_1 _0890_ (.B1(net146),
    .Y(_0290_),
    .A1(\ltc.output_buffer[29] ),
    .A2(net142));
 sg13g2_nand3_1 _0891_ (.B(net293),
    .C(net156),
    .A(net175),
    .Y(_0291_));
 sg13g2_o21ai_1 _0892_ (.B1(_0291_),
    .Y(_0029_),
    .A1(_0289_),
    .A2(_0290_));
 sg13g2_nor2_1 _0893_ (.A(\ltc.hrs_u[1] ),
    .B(net138),
    .Y(_0292_));
 sg13g2_o21ai_1 _0894_ (.B1(net146),
    .Y(_0293_),
    .A1(net331),
    .A2(net142));
 sg13g2_nand3_1 _0895_ (.B(net335),
    .C(net156),
    .A(net175),
    .Y(_0294_));
 sg13g2_o21ai_1 _0896_ (.B1(_0294_),
    .Y(_0030_),
    .A1(_0292_),
    .A2(_0293_));
 sg13g2_nor2_1 _0897_ (.A(\ltc.output_buffer[31] ),
    .B(net142),
    .Y(_0295_));
 sg13g2_o21ai_1 _0898_ (.B1(net146),
    .Y(_0296_),
    .A1(\ltc.hrs_u[0] ),
    .A2(net138));
 sg13g2_nand3_1 _0899_ (.B(net331),
    .C(net151),
    .A(net175),
    .Y(_0297_));
 sg13g2_o21ai_1 _0900_ (.B1(_0297_),
    .Y(_0031_),
    .A1(_0295_),
    .A2(_0296_));
 sg13g2_a22oi_1 _0901_ (.Y(_0298_),
    .B1(net129),
    .B2(net333),
    .A2(net150),
    .A1(\ltc.output_buffer[31] ));
 sg13g2_nor2_1 _0902_ (.A(net165),
    .B(net334),
    .Y(_0032_));
 sg13g2_a22oi_1 _0903_ (.Y(_0299_),
    .B1(net129),
    .B2(net392),
    .A2(net150),
    .A1(net333));
 sg13g2_nor2_1 _0904_ (.A(net165),
    .B(_0299_),
    .Y(_0033_));
 sg13g2_a22oi_1 _0905_ (.Y(_0300_),
    .B1(net129),
    .B2(net324),
    .A2(net150),
    .A1(\ltc.output_buffer[33] ));
 sg13g2_nor2_1 _0906_ (.A(net165),
    .B(net325),
    .Y(_0034_));
 sg13g2_a22oi_1 _0907_ (.Y(_0301_),
    .B1(net129),
    .B2(net341),
    .A2(net150),
    .A1(net324));
 sg13g2_nor2_1 _0908_ (.A(net165),
    .B(_0301_),
    .Y(_0035_));
 sg13g2_a22oi_1 _0909_ (.Y(_0302_),
    .B1(net129),
    .B2(net291),
    .A2(net150),
    .A1(net341));
 sg13g2_nor2_1 _0910_ (.A(net165),
    .B(_0302_),
    .Y(_0036_));
 sg13g2_nand3_1 _0911_ (.B(net291),
    .C(net150),
    .A(net175),
    .Y(_0303_));
 sg13g2_nor2_1 _0912_ (.A(\ltc.output_buffer[37] ),
    .B(net142),
    .Y(_0304_));
 sg13g2_o21ai_1 _0913_ (.B1(net146),
    .Y(_0305_),
    .A1(\ltc.min_d[2] ),
    .A2(net138));
 sg13g2_o21ai_1 _0914_ (.B1(_0303_),
    .Y(_0037_),
    .A1(_0304_),
    .A2(_0305_));
 sg13g2_nor2_1 _0915_ (.A(\ltc.min_d[1] ),
    .B(net138),
    .Y(_0306_));
 sg13g2_o21ai_1 _0916_ (.B1(net146),
    .Y(_0307_),
    .A1(\ltc.output_buffer[38] ),
    .A2(net142));
 sg13g2_nand3_1 _0917_ (.B(net301),
    .C(net151),
    .A(net175),
    .Y(_0308_));
 sg13g2_o21ai_1 _0918_ (.B1(_0308_),
    .Y(_0038_),
    .A1(_0306_),
    .A2(_0307_));
 sg13g2_nor2_1 _0919_ (.A(\ltc.min_d[0] ),
    .B(net138),
    .Y(_0309_));
 sg13g2_o21ai_1 _0920_ (.B1(net146),
    .Y(_0310_),
    .A1(\ltc.output_buffer[39] ),
    .A2(net142));
 sg13g2_nand3_1 _0921_ (.B(net307),
    .C(net151),
    .A(net176),
    .Y(_0311_));
 sg13g2_o21ai_1 _0922_ (.B1(_0311_),
    .Y(_0039_),
    .A1(_0309_),
    .A2(_0310_));
 sg13g2_a22oi_1 _0923_ (.Y(_0312_),
    .B1(net129),
    .B2(net364),
    .A2(net151),
    .A1(\ltc.output_buffer[39] ));
 sg13g2_nor2_1 _0924_ (.A(net168),
    .B(net365),
    .Y(_0040_));
 sg13g2_a22oi_1 _0925_ (.Y(_0313_),
    .B1(net130),
    .B2(net388),
    .A2(net151),
    .A1(net364));
 sg13g2_nor2_1 _0926_ (.A(net168),
    .B(_0313_),
    .Y(_0041_));
 sg13g2_a22oi_1 _0927_ (.Y(_0314_),
    .B1(net130),
    .B2(net311),
    .A2(net156),
    .A1(\ltc.output_buffer[41] ));
 sg13g2_nor2_1 _0928_ (.A(net170),
    .B(net312),
    .Y(_0042_));
 sg13g2_a22oi_1 _0929_ (.Y(_0315_),
    .B1(net130),
    .B2(net372),
    .A2(net156),
    .A1(net311));
 sg13g2_nor2_1 _0930_ (.A(net170),
    .B(_0315_),
    .Y(_0043_));
 sg13g2_nand3_1 _0931_ (.B(net372),
    .C(net156),
    .A(net177),
    .Y(_0316_));
 sg13g2_nor2_1 _0932_ (.A(\ltc.min_u[3] ),
    .B(net139),
    .Y(_0317_));
 sg13g2_o21ai_1 _0933_ (.B1(net147),
    .Y(_0318_),
    .A1(net351),
    .A2(net143));
 sg13g2_o21ai_1 _0934_ (.B1(_0316_),
    .Y(_0044_),
    .A1(_0317_),
    .A2(_0318_));
 sg13g2_nor2_1 _0935_ (.A(\ltc.min_u[2] ),
    .B(net139),
    .Y(_0319_));
 sg13g2_o21ai_1 _0936_ (.B1(net147),
    .Y(_0320_),
    .A1(net299),
    .A2(net143));
 sg13g2_nand3_1 _0937_ (.B(net351),
    .C(net156),
    .A(net176),
    .Y(_0321_));
 sg13g2_o21ai_1 _0938_ (.B1(_0321_),
    .Y(_0045_),
    .A1(_0319_),
    .A2(_0320_));
 sg13g2_nor2_1 _0939_ (.A(\ltc.min_u[1] ),
    .B(net139),
    .Y(_0322_));
 sg13g2_o21ai_1 _0940_ (.B1(net147),
    .Y(_0323_),
    .A1(net286),
    .A2(net143));
 sg13g2_nand3_1 _0941_ (.B(net299),
    .C(net158),
    .A(net176),
    .Y(_0324_));
 sg13g2_o21ai_1 _0942_ (.B1(_0324_),
    .Y(_0046_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_nor2_1 _0943_ (.A(\ltc.min_u[0] ),
    .B(net139),
    .Y(_0325_));
 sg13g2_o21ai_1 _0944_ (.B1(net147),
    .Y(_0326_),
    .A1(\ltc.output_buffer[47] ),
    .A2(net143));
 sg13g2_nand3_1 _0945_ (.B(net286),
    .C(net158),
    .A(net176),
    .Y(_0327_));
 sg13g2_o21ai_1 _0946_ (.B1(_0327_),
    .Y(_0047_),
    .A1(_0325_),
    .A2(_0326_));
 sg13g2_a22oi_1 _0947_ (.Y(_0328_),
    .B1(net134),
    .B2(net383),
    .A2(net158),
    .A1(\ltc.output_buffer[47] ));
 sg13g2_nor2_1 _0948_ (.A(net170),
    .B(net384),
    .Y(_0048_));
 sg13g2_a22oi_1 _0949_ (.Y(_0329_),
    .B1(net134),
    .B2(net342),
    .A2(net158),
    .A1(\ltc.output_buffer[48] ));
 sg13g2_nor2_1 _0950_ (.A(net170),
    .B(net343),
    .Y(_0049_));
 sg13g2_a22oi_1 _0951_ (.Y(_0330_),
    .B1(net134),
    .B2(net370),
    .A2(net158),
    .A1(net342));
 sg13g2_nor2_1 _0952_ (.A(net170),
    .B(_0330_),
    .Y(_0050_));
 sg13g2_a22oi_1 _0953_ (.Y(_0331_),
    .B1(net134),
    .B2(net270),
    .A2(net158),
    .A1(net370));
 sg13g2_nor2_1 _0954_ (.A(net170),
    .B(_0331_),
    .Y(_0051_));
 sg13g2_nand2_1 _0955_ (.Y(_0332_),
    .A(net270),
    .B(net158));
 sg13g2_nor2_2 _0956_ (.A(net4),
    .B(net3),
    .Y(_0333_));
 sg13g2_and2_1 _0957_ (.A(net4),
    .B(net3),
    .X(_0334_));
 sg13g2_o21ai_1 _0958_ (.B1(_0206_),
    .Y(_0335_),
    .A1(_0333_),
    .A2(_0334_));
 sg13g2_nand2_1 _0959_ (.Y(_0336_),
    .A(\ltc.output_buffer[52] ),
    .B(net141));
 sg13g2_a21oi_1 _0960_ (.A1(_0335_),
    .A2(_0336_),
    .Y(_0337_),
    .B1(net158));
 sg13g2_o21ai_1 _0961_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0271_),
    .A2(_0335_));
 sg13g2_a21oi_1 _0962_ (.A1(_0332_),
    .A2(_0338_),
    .Y(_0052_),
    .B1(net171));
 sg13g2_nor2_1 _0963_ (.A(\ltc.sec_d[2] ),
    .B(net141),
    .Y(_0339_));
 sg13g2_o21ai_1 _0964_ (.B1(net149),
    .Y(_0340_),
    .A1(net272),
    .A2(net145));
 sg13g2_nand3_1 _0965_ (.B(net303),
    .C(net159),
    .A(net178),
    .Y(_0341_));
 sg13g2_o21ai_1 _0966_ (.B1(_0341_),
    .Y(_0053_),
    .A1(_0339_),
    .A2(_0340_));
 sg13g2_nor2_1 _0967_ (.A(\ltc.sec_d[1] ),
    .B(net141),
    .Y(_0342_));
 sg13g2_o21ai_1 _0968_ (.B1(net149),
    .Y(_0343_),
    .A1(net265),
    .A2(net145));
 sg13g2_nand3_1 _0969_ (.B(net272),
    .C(net159),
    .A(net178),
    .Y(_0344_));
 sg13g2_o21ai_1 _0970_ (.B1(_0344_),
    .Y(_0054_),
    .A1(_0342_),
    .A2(_0343_));
 sg13g2_nor2_1 _0971_ (.A(\ltc.sec_d[0] ),
    .B(net141),
    .Y(_0345_));
 sg13g2_o21ai_1 _0972_ (.B1(net149),
    .Y(_0346_),
    .A1(\ltc.output_buffer[55] ),
    .A2(net145));
 sg13g2_nand3_1 _0973_ (.B(net265),
    .C(net159),
    .A(net178),
    .Y(_0347_));
 sg13g2_o21ai_1 _0974_ (.B1(_0347_),
    .Y(_0055_),
    .A1(_0345_),
    .A2(_0346_));
 sg13g2_a22oi_1 _0975_ (.Y(_0348_),
    .B1(net134),
    .B2(net337),
    .A2(net159),
    .A1(\ltc.output_buffer[55] ));
 sg13g2_nor2_1 _0976_ (.A(net171),
    .B(net338),
    .Y(_0056_));
 sg13g2_a22oi_1 _0977_ (.Y(_0349_),
    .B1(net134),
    .B2(net344),
    .A2(net159),
    .A1(net337));
 sg13g2_nor2_1 _0978_ (.A(net171),
    .B(_0349_),
    .Y(_0057_));
 sg13g2_a22oi_1 _0979_ (.Y(_0350_),
    .B1(net134),
    .B2(net345),
    .A2(net160),
    .A1(net344));
 sg13g2_nor2_1 _0980_ (.A(net171),
    .B(_0350_),
    .Y(_0058_));
 sg13g2_a22oi_1 _0981_ (.Y(_0351_),
    .B1(net136),
    .B2(net366),
    .A2(net161),
    .A1(net345));
 sg13g2_nor2_1 _0982_ (.A(net171),
    .B(_0351_),
    .Y(_0059_));
 sg13g2_nand3_1 _0983_ (.B(net366),
    .C(net159),
    .A(net179),
    .Y(_0352_));
 sg13g2_nor2_1 _0984_ (.A(\ltc.sec_u[3] ),
    .B(net141),
    .Y(_0353_));
 sg13g2_o21ai_1 _0985_ (.B1(net149),
    .Y(_0354_),
    .A1(net280),
    .A2(net144));
 sg13g2_o21ai_1 _0986_ (.B1(_0352_),
    .Y(_0060_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_nor2_1 _0987_ (.A(\ltc.output_buffer[61] ),
    .B(net144),
    .Y(_0355_));
 sg13g2_o21ai_1 _0988_ (.B1(net148),
    .Y(_0356_),
    .A1(\ltc.sec_u[2] ),
    .A2(net140));
 sg13g2_nand3_1 _0989_ (.B(net280),
    .C(net163),
    .A(net178),
    .Y(_0357_));
 sg13g2_o21ai_1 _0990_ (.B1(_0357_),
    .Y(_0061_),
    .A1(_0355_),
    .A2(_0356_));
 sg13g2_nor2_1 _0991_ (.A(\ltc.sec_u[1] ),
    .B(net140),
    .Y(_0358_));
 sg13g2_o21ai_1 _0992_ (.B1(net148),
    .Y(_0359_),
    .A1(net284),
    .A2(net145));
 sg13g2_nand3_1 _0993_ (.B(net305),
    .C(net163),
    .A(net178),
    .Y(_0360_));
 sg13g2_o21ai_1 _0994_ (.B1(_0360_),
    .Y(_0062_),
    .A1(_0358_),
    .A2(_0359_));
 sg13g2_nor2_1 _0995_ (.A(\ltc.output_buffer[63] ),
    .B(net144),
    .Y(_0361_));
 sg13g2_o21ai_1 _0996_ (.B1(net148),
    .Y(_0362_),
    .A1(\ltc.sec_u[0] ),
    .A2(net140));
 sg13g2_nand3_1 _0997_ (.B(net284),
    .C(net163),
    .A(net179),
    .Y(_0363_));
 sg13g2_o21ai_1 _0998_ (.B1(_0363_),
    .Y(_0063_),
    .A1(_0361_),
    .A2(_0362_));
 sg13g2_a22oi_1 _0999_ (.Y(_0364_),
    .B1(net136),
    .B2(net320),
    .A2(net160),
    .A1(\ltc.output_buffer[63] ));
 sg13g2_nor2_1 _1000_ (.A(net171),
    .B(net321),
    .Y(_0064_));
 sg13g2_a22oi_1 _1001_ (.Y(_0365_),
    .B1(net135),
    .B2(net376),
    .A2(net160),
    .A1(net320));
 sg13g2_nor2_1 _1002_ (.A(net169),
    .B(_0365_),
    .Y(_0065_));
 sg13g2_a22oi_1 _1003_ (.Y(_0366_),
    .B1(net135),
    .B2(net315),
    .A2(net160),
    .A1(\ltc.output_buffer[65] ));
 sg13g2_nor2_1 _1004_ (.A(net169),
    .B(net316),
    .Y(_0066_));
 sg13g2_a22oi_1 _1005_ (.Y(_0367_),
    .B1(net135),
    .B2(net377),
    .A2(net160),
    .A1(net315));
 sg13g2_nor2_1 _1006_ (.A(net174),
    .B(_0367_),
    .Y(_0067_));
 sg13g2_a22oi_1 _1007_ (.Y(_0368_),
    .B1(net135),
    .B2(net349),
    .A2(net160),
    .A1(\ltc.output_buffer[67] ));
 sg13g2_nor2_1 _1008_ (.A(net172),
    .B(net350),
    .Y(_0068_));
 sg13g2_a22oi_1 _1009_ (.Y(_0369_),
    .B1(net135),
    .B2(net322),
    .A2(net160),
    .A1(net349));
 sg13g2_nor2_1 _1010_ (.A(net171),
    .B(_0369_),
    .Y(_0069_));
 sg13g2_nand3_1 _1011_ (.B(net322),
    .C(net160),
    .A(net179),
    .Y(_0370_));
 sg13g2_nor2_1 _1012_ (.A(\ltc.frm_d[1] ),
    .B(net140),
    .Y(_0371_));
 sg13g2_o21ai_1 _1013_ (.B1(net148),
    .Y(_0372_),
    .A1(\ltc.output_buffer[70] ),
    .A2(net144));
 sg13g2_o21ai_1 _1014_ (.B1(_0370_),
    .Y(_0070_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_nor2_1 _1015_ (.A(\ltc.frm_d[0] ),
    .B(net140),
    .Y(_0373_));
 sg13g2_o21ai_1 _1016_ (.B1(net149),
    .Y(_0374_),
    .A1(\ltc.output_buffer[71] ),
    .A2(net144));
 sg13g2_nand3_1 _1017_ (.B(net362),
    .C(net163),
    .A(net179),
    .Y(_0375_));
 sg13g2_o21ai_1 _1018_ (.B1(_0375_),
    .Y(_0071_),
    .A1(_0373_),
    .A2(_0374_));
 sg13g2_a22oi_1 _1019_ (.Y(_0376_),
    .B1(net135),
    .B2(net329),
    .A2(net161),
    .A1(\ltc.output_buffer[71] ));
 sg13g2_nor2_1 _1020_ (.A(net171),
    .B(net330),
    .Y(_0072_));
 sg13g2_a22oi_1 _1021_ (.Y(_0377_),
    .B1(net136),
    .B2(net389),
    .A2(net161),
    .A1(net329));
 sg13g2_nor2_1 _1022_ (.A(net172),
    .B(_0377_),
    .Y(_0073_));
 sg13g2_a22oi_1 _1023_ (.Y(_0378_),
    .B1(net135),
    .B2(net339),
    .A2(net161),
    .A1(\ltc.output_buffer[73] ));
 sg13g2_nor2_1 _1024_ (.A(net172),
    .B(net340),
    .Y(_0074_));
 sg13g2_a22oi_1 _1025_ (.Y(_0379_),
    .B1(net135),
    .B2(net297),
    .A2(net161),
    .A1(net339));
 sg13g2_nor2_1 _1026_ (.A(net172),
    .B(_0379_),
    .Y(_0075_));
 sg13g2_nand3_1 _1027_ (.B(net297),
    .C(net164),
    .A(net179),
    .Y(_0380_));
 sg13g2_nor2_1 _1028_ (.A(\ltc.frm_u[3] ),
    .B(net140),
    .Y(_0381_));
 sg13g2_o21ai_1 _1029_ (.B1(net148),
    .Y(_0382_),
    .A1(\ltc.output_buffer[76] ),
    .A2(net144));
 sg13g2_o21ai_1 _1030_ (.B1(_0380_),
    .Y(_0076_),
    .A1(_0381_),
    .A2(_0382_));
 sg13g2_nor2_1 _1031_ (.A(net313),
    .B(net144),
    .Y(_0383_));
 sg13g2_o21ai_1 _1032_ (.B1(net148),
    .Y(_0384_),
    .A1(\ltc.frm_u[2] ),
    .A2(net140));
 sg13g2_nand3_1 _1033_ (.B(net378),
    .C(net163),
    .A(net179),
    .Y(_0385_));
 sg13g2_o21ai_1 _1034_ (.B1(_0385_),
    .Y(_0077_),
    .A1(_0383_),
    .A2(_0384_));
 sg13g2_nor2_1 _1035_ (.A(\ltc.frm_u[1] ),
    .B(net140),
    .Y(_0386_));
 sg13g2_o21ai_1 _1036_ (.B1(net148),
    .Y(_0387_),
    .A1(\ltc.output_buffer[78] ),
    .A2(net145));
 sg13g2_nand3_1 _1037_ (.B(net313),
    .C(net163),
    .A(net180),
    .Y(_0388_));
 sg13g2_o21ai_1 _1038_ (.B1(_0388_),
    .Y(_0078_),
    .A1(_0386_),
    .A2(_0387_));
 sg13g2_nor2_1 _1039_ (.A(net328),
    .B(net141),
    .Y(_0389_));
 sg13g2_o21ai_1 _1040_ (.B1(net148),
    .Y(_0390_),
    .A1(\ltc.output_buffer[79] ),
    .A2(net144));
 sg13g2_nand3_1 _1041_ (.B(net358),
    .C(net163),
    .A(net180),
    .Y(_0391_));
 sg13g2_o21ai_1 _1042_ (.B1(_0391_),
    .Y(_0079_),
    .A1(_0389_),
    .A2(_0390_));
 sg13g2_nand3b_1 _1043_ (.B(net400),
    .C(net380),
    .Y(_0392_),
    .A_N(net317));
 sg13g2_nor2_1 _1044_ (.A(_0151_),
    .B(_0392_),
    .Y(_0393_));
 sg13g2_nor4_1 _1045_ (.A(net393),
    .B(_0150_),
    .C(net429),
    .D(net426),
    .Y(_0394_));
 sg13g2_nand3b_1 _1046_ (.B(net434),
    .C(_0394_),
    .Y(_0395_),
    .A_N(net439));
 sg13g2_nand2_1 _1047_ (.Y(_0396_),
    .A(net439),
    .B(net393));
 sg13g2_nor3_2 _1048_ (.A(net434),
    .B(net426),
    .C(_0396_),
    .Y(_0397_));
 sg13g2_nor2_1 _1049_ (.A(_0392_),
    .B(_0397_),
    .Y(_0398_));
 sg13g2_a21oi_1 _1050_ (.A1(_0395_),
    .A2(_0398_),
    .Y(_0399_),
    .B1(net426));
 sg13g2_o21ai_1 _1051_ (.B1(net175),
    .Y(_0080_),
    .A1(_0393_),
    .A2(net427));
 sg13g2_and4_1 _1052_ (.A(\ltc.frm_counter[3] ),
    .B(net274),
    .C(net230),
    .D(\ltc.frm_counter[1] ),
    .X(_0400_));
 sg13g2_nand4_1 _1053_ (.B(net274),
    .C(net230),
    .A(net443),
    .Y(_0401_),
    .D(\ltc.frm_counter[1] ));
 sg13g2_nand2_1 _1054_ (.Y(_0402_),
    .A(\ltc.frm_counter[6] ),
    .B(\ltc.frm_counter[7] ));
 sg13g2_and4_1 _1055_ (.A(\ltc.frm_counter[5] ),
    .B(\ltc.frm_counter[4] ),
    .C(\ltc.frm_counter[6] ),
    .D(\ltc.frm_counter[7] ),
    .X(_0403_));
 sg13g2_nand4_1 _1056_ (.B(\ltc.frm_counter[4] ),
    .C(\ltc.frm_counter[6] ),
    .A(\ltc.frm_counter[5] ),
    .Y(_0404_),
    .D(\ltc.frm_counter[7] ));
 sg13g2_nor2_1 _1057_ (.A(_0401_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_nand2_1 _1058_ (.Y(_0406_),
    .A(_0400_),
    .B(_0403_));
 sg13g2_nand4_1 _1059_ (.B(\ltc.frm_counter[8] ),
    .C(\ltc.frm_counter[10] ),
    .A(\ltc.frm_counter[9] ),
    .Y(_0407_),
    .D(net419));
 sg13g2_nor3_1 _1060_ (.A(_0401_),
    .B(_0404_),
    .C(_0407_),
    .Y(_0408_));
 sg13g2_nor4_2 _1061_ (.A(_0152_),
    .B(_0401_),
    .C(_0404_),
    .Y(_0409_),
    .D(_0407_));
 sg13g2_nand2_1 _1062_ (.Y(_0410_),
    .A(net460),
    .B(_0409_));
 sg13g2_nand3_1 _1063_ (.B(net472),
    .C(_0409_),
    .A(net460),
    .Y(_0411_));
 sg13g2_and4_1 _1064_ (.A(\ltc.frm_counter[13] ),
    .B(\ltc.frm_counter[14] ),
    .C(net455),
    .D(_0409_),
    .X(_0412_));
 sg13g2_and2_1 _1065_ (.A(net458),
    .B(_0412_),
    .X(_0413_));
 sg13g2_nand3_1 _1066_ (.B(\ltc.frm_counter[17] ),
    .C(_0412_),
    .A(\ltc.frm_counter[16] ),
    .Y(_0414_));
 sg13g2_nand3_1 _1067_ (.B(\ltc.frm_counter[18] ),
    .C(_0413_),
    .A(\ltc.frm_counter[17] ),
    .Y(_0415_));
 sg13g2_xor2_1 _1068_ (.B(_0414_),
    .A(net448),
    .X(_0416_));
 sg13g2_or2_1 _1069_ (.X(_0417_),
    .B(_0416_),
    .A(_0186_));
 sg13g2_xnor2_1 _1070_ (.Y(_0418_),
    .A(_0153_),
    .B(_0413_));
 sg13g2_xnor2_1 _1071_ (.Y(_0419_),
    .A(net458),
    .B(_0412_));
 sg13g2_xnor2_1 _1072_ (.Y(_0420_),
    .A(net468),
    .B(_0408_));
 sg13g2_or2_1 _1073_ (.X(_0421_),
    .B(_0409_),
    .A(net460));
 sg13g2_nor2_1 _1074_ (.A(net474),
    .B(_0420_),
    .Y(_0422_));
 sg13g2_and3_1 _1075_ (.X(_0423_),
    .A(net416),
    .B(net422),
    .C(_0400_));
 sg13g2_and4_1 _1076_ (.A(net416),
    .B(net422),
    .C(net451),
    .D(_0400_),
    .X(_0424_));
 sg13g2_nor2b_1 _1077_ (.A(\ltc.frm_counter[8] ),
    .B_N(\ltc.frm_counter[9] ),
    .Y(_0425_));
 sg13g2_nand2_1 _1078_ (.Y(_0426_),
    .A(\ltc.frm_counter[11] ),
    .B(_0425_));
 sg13g2_nand3_1 _1079_ (.B(_0334_),
    .C(_0402_),
    .A(_0187_),
    .Y(_0427_));
 sg13g2_nor3_1 _1080_ (.A(\ltc.frm_counter[10] ),
    .B(_0426_),
    .C(_0427_),
    .Y(_0428_));
 sg13g2_and2_1 _1081_ (.A(_0424_),
    .B(_0428_),
    .X(_0429_));
 sg13g2_nand4_1 _1082_ (.B(_0419_),
    .C(_0422_),
    .A(_0418_),
    .Y(_0430_),
    .D(_0429_));
 sg13g2_and4_1 _1083_ (.A(\ltc.frm_counter[9] ),
    .B(\ltc.frm_counter[8] ),
    .C(_0400_),
    .D(_0403_),
    .X(_0431_));
 sg13g2_a21oi_1 _1084_ (.A1(\ltc.frm_counter[10] ),
    .A2(_0431_),
    .Y(_0432_),
    .B1(net419));
 sg13g2_xnor2_1 _1085_ (.Y(_0433_),
    .A(net453),
    .B(_0431_));
 sg13g2_o21ai_1 _1086_ (.B1(_0433_),
    .Y(_0434_),
    .A1(_0408_),
    .A2(_0432_));
 sg13g2_nor3_1 _1087_ (.A(_0153_),
    .B(_0419_),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_xor2_1 _1088_ (.B(_0411_),
    .A(net455),
    .X(_0436_));
 sg13g2_a21oi_1 _1089_ (.A1(_0400_),
    .A2(_0403_),
    .Y(_0437_),
    .B1(net466));
 sg13g2_or3_1 _1090_ (.A(_0188_),
    .B(_0431_),
    .C(net467),
    .X(_0438_));
 sg13g2_o21ai_1 _1091_ (.B1(_0406_),
    .Y(_0439_),
    .A1(net465),
    .A2(_0424_));
 sg13g2_nand4_1 _1092_ (.B(_0421_),
    .C(_0438_),
    .A(_0420_),
    .Y(_0440_),
    .D(_0439_));
 sg13g2_xnor2_1 _1093_ (.Y(_0441_),
    .A(net451),
    .B(_0423_));
 sg13g2_and2_1 _1094_ (.A(net422),
    .B(_0400_),
    .X(_0442_));
 sg13g2_nor3_1 _1095_ (.A(\ltc.frm_counter[5] ),
    .B(net4),
    .C(net3),
    .Y(_0443_));
 sg13g2_xnor2_1 _1096_ (.Y(_0444_),
    .A(net463),
    .B(_0406_));
 sg13g2_nand4_1 _1097_ (.B(_0442_),
    .C(_0443_),
    .A(_0441_),
    .Y(_0445_),
    .D(_0444_));
 sg13g2_a21o_1 _1098_ (.A2(_0409_),
    .A1(net460),
    .B1(net472),
    .X(_0446_));
 sg13g2_nor4_1 _1099_ (.A(_0436_),
    .B(_0440_),
    .C(_0445_),
    .D(_0446_),
    .Y(_0447_));
 sg13g2_nand4_1 _1100_ (.B(_0405_),
    .C(_0425_),
    .A(_0207_),
    .Y(_0448_),
    .D(_0446_));
 sg13g2_nor4_1 _1101_ (.A(\ltc.frm_counter[13] ),
    .B(\ltc.frm_counter[15] ),
    .C(_0420_),
    .D(_0448_),
    .Y(_0449_));
 sg13g2_o21ai_1 _1102_ (.B1(_0435_),
    .Y(_0450_),
    .A1(_0447_),
    .A2(_0449_));
 sg13g2_a21oi_2 _1103_ (.B1(_0417_),
    .Y(_0451_),
    .A2(_0450_),
    .A1(_0430_));
 sg13g2_a21o_2 _1104_ (.A2(_0450_),
    .A1(_0430_),
    .B1(_0417_),
    .X(_0452_));
 sg13g2_nand2_1 _1105_ (.Y(_0453_),
    .A(net179),
    .B(_0452_));
 sg13g2_nor2_1 _1106_ (.A(net230),
    .B(net125),
    .Y(_0081_));
 sg13g2_nor2_1 _1107_ (.A(_0192_),
    .B(_0205_),
    .Y(_0454_));
 sg13g2_nor2_1 _1108_ (.A(net125),
    .B(_0454_),
    .Y(_0082_));
 sg13g2_and3_1 _1109_ (.X(_0455_),
    .A(net274),
    .B(net230),
    .C(\ltc.frm_counter[1] ));
 sg13g2_a21oi_1 _1110_ (.A1(net230),
    .A2(\ltc.frm_counter[1] ),
    .Y(_0456_),
    .B1(net274));
 sg13g2_nor3_1 _1111_ (.A(net125),
    .B(_0455_),
    .C(net275),
    .Y(_0083_));
 sg13g2_o21ai_1 _1112_ (.B1(_0401_),
    .Y(_0457_),
    .A1(net443),
    .A2(_0455_));
 sg13g2_nor2_1 _1113_ (.A(net125),
    .B(net444),
    .Y(_0084_));
 sg13g2_nor2_1 _1114_ (.A(net422),
    .B(_0400_),
    .Y(_0458_));
 sg13g2_nor3_1 _1115_ (.A(_0442_),
    .B(net126),
    .C(net423),
    .Y(_0085_));
 sg13g2_nor2_1 _1116_ (.A(net416),
    .B(_0442_),
    .Y(_0459_));
 sg13g2_nor3_1 _1117_ (.A(_0423_),
    .B(net126),
    .C(net417),
    .Y(_0086_));
 sg13g2_nor2_1 _1118_ (.A(_0441_),
    .B(net126),
    .Y(_0087_));
 sg13g2_nor2_1 _1119_ (.A(_0439_),
    .B(net126),
    .Y(_0088_));
 sg13g2_nor2b_1 _1120_ (.A(net126),
    .B_N(_0444_),
    .Y(_0089_));
 sg13g2_nor2_1 _1121_ (.A(_0438_),
    .B(net127),
    .Y(_0090_));
 sg13g2_nor2_1 _1122_ (.A(net454),
    .B(net127),
    .Y(_0091_));
 sg13g2_nor3_1 _1123_ (.A(_0408_),
    .B(net420),
    .C(net127),
    .Y(_0092_));
 sg13g2_nor2_1 _1124_ (.A(_0420_),
    .B(net126),
    .Y(_0093_));
 sg13g2_and4_1 _1125_ (.A(net180),
    .B(_0410_),
    .C(_0421_),
    .D(net128),
    .X(_0094_));
 sg13g2_and4_1 _1126_ (.A(net180),
    .B(_0411_),
    .C(_0446_),
    .D(net128),
    .X(_0095_));
 sg13g2_nor2_1 _1127_ (.A(net456),
    .B(net126),
    .Y(_0096_));
 sg13g2_nor2_1 _1128_ (.A(net459),
    .B(net126),
    .Y(_0097_));
 sg13g2_and3_1 _1129_ (.X(_0098_),
    .A(net180),
    .B(_0418_),
    .C(net128));
 sg13g2_nor2_1 _1130_ (.A(net449),
    .B(net125),
    .Y(_0099_));
 sg13g2_and4_1 _1131_ (.A(\ltc.frm_counter[17] ),
    .B(\ltc.frm_counter[18] ),
    .C(net257),
    .D(_0413_),
    .X(_0460_));
 sg13g2_nor2b_1 _1132_ (.A(net257),
    .B_N(_0415_),
    .Y(_0461_));
 sg13g2_nor3_1 _1133_ (.A(net125),
    .B(_0460_),
    .C(net258),
    .Y(_0100_));
 sg13g2_xnor2_1 _1134_ (.Y(_0462_),
    .A(net390),
    .B(_0460_));
 sg13g2_nor2_1 _1135_ (.A(net125),
    .B(net391),
    .Y(_0101_));
 sg13g2_and3_1 _1136_ (.X(_0463_),
    .A(\ltc.frm_counter[20] ),
    .B(net239),
    .C(_0460_));
 sg13g2_a21oi_1 _1137_ (.A1(\ltc.frm_counter[20] ),
    .A2(_0460_),
    .Y(_0464_),
    .B1(net239));
 sg13g2_nor3_1 _1138_ (.A(net125),
    .B(_0463_),
    .C(net240),
    .Y(_0102_));
 sg13g2_nor2_1 _1139_ (.A(net355),
    .B(_0463_),
    .Y(_0465_));
 sg13g2_and2_1 _1140_ (.A(net355),
    .B(_0463_),
    .X(_0466_));
 sg13g2_nor3_1 _1141_ (.A(net127),
    .B(net356),
    .C(_0466_),
    .Y(_0103_));
 sg13g2_nor2_1 _1142_ (.A(net374),
    .B(_0466_),
    .Y(_0467_));
 sg13g2_and2_1 _1143_ (.A(net374),
    .B(_0466_),
    .X(_0468_));
 sg13g2_nor3_1 _1144_ (.A(net127),
    .B(net375),
    .C(_0468_),
    .Y(_0104_));
 sg13g2_nand2_1 _1145_ (.Y(_0469_),
    .A(net175),
    .B(_0395_));
 sg13g2_nand2_1 _1146_ (.Y(_0470_),
    .A(net429),
    .B(_0397_));
 sg13g2_xnor2_1 _1147_ (.Y(_0471_),
    .A(net429),
    .B(_0397_));
 sg13g2_nor2_1 _1148_ (.A(_0469_),
    .B(net430),
    .Y(_0105_));
 sg13g2_xnor2_1 _1149_ (.Y(_0472_),
    .A(_0150_),
    .B(_0470_));
 sg13g2_nor2_1 _1150_ (.A(_0469_),
    .B(_0472_),
    .Y(_0106_));
 sg13g2_or2_1 _1151_ (.X(_0473_),
    .B(_0469_),
    .A(_0397_));
 sg13g2_and2_1 _1152_ (.A(net393),
    .B(_0393_),
    .X(_0474_));
 sg13g2_nor2_1 _1153_ (.A(net393),
    .B(_0393_),
    .Y(_0475_));
 sg13g2_nor3_1 _1154_ (.A(_0473_),
    .B(_0474_),
    .C(net394),
    .Y(_0107_));
 sg13g2_nand2_1 _1155_ (.Y(_0476_),
    .A(net434),
    .B(_0474_));
 sg13g2_xnor2_1 _1156_ (.Y(_0477_),
    .A(net434),
    .B(_0474_));
 sg13g2_nor2_1 _1157_ (.A(_0473_),
    .B(_0477_),
    .Y(_0108_));
 sg13g2_xor2_1 _1158_ (.B(_0476_),
    .A(net439),
    .X(_0478_));
 sg13g2_nor2_1 _1159_ (.A(_0473_),
    .B(_0478_),
    .Y(_0109_));
 sg13g2_nand2_1 _1160_ (.Y(_0479_),
    .A(\ltc.min_u[3] ),
    .B(net398));
 sg13g2_nor3_1 _1161_ (.A(net404),
    .B(\ltc.min_u[0] ),
    .C(_0479_),
    .Y(_0480_));
 sg13g2_and2_1 _1162_ (.A(net317),
    .B(_0480_),
    .X(_0481_));
 sg13g2_nand2_1 _1163_ (.Y(_0482_),
    .A(net175),
    .B(_0392_));
 sg13g2_nor2_1 _1164_ (.A(net317),
    .B(_0480_),
    .Y(_0483_));
 sg13g2_nor3_1 _1165_ (.A(_0481_),
    .B(_0482_),
    .C(net318),
    .Y(_0110_));
 sg13g2_nor2_1 _1166_ (.A(net400),
    .B(_0481_),
    .Y(_0484_));
 sg13g2_and2_1 _1167_ (.A(net400),
    .B(_0481_),
    .X(_0485_));
 sg13g2_nor3_1 _1168_ (.A(_0482_),
    .B(net401),
    .C(_0485_),
    .Y(_0111_));
 sg13g2_xnor2_1 _1169_ (.Y(_0486_),
    .A(net380),
    .B(_0485_));
 sg13g2_nor2_1 _1170_ (.A(_0482_),
    .B(net381),
    .Y(_0112_));
 sg13g2_nand3b_1 _1171_ (.B(net402),
    .C(net395),
    .Y(_0487_),
    .A_N(net346));
 sg13g2_nor2_1 _1172_ (.A(_0149_),
    .B(_0487_),
    .Y(_0488_));
 sg13g2_nand2b_2 _1173_ (.Y(_0489_),
    .B(net176),
    .A_N(_0480_));
 sg13g2_and2_1 _1174_ (.A(_0149_),
    .B(_0487_),
    .X(_0490_));
 sg13g2_nor3_1 _1175_ (.A(_0488_),
    .B(_0489_),
    .C(_0490_),
    .Y(_0113_));
 sg13g2_and2_1 _1176_ (.A(net398),
    .B(_0488_),
    .X(_0491_));
 sg13g2_nor2_1 _1177_ (.A(net398),
    .B(_0488_),
    .Y(_0492_));
 sg13g2_nor3_1 _1178_ (.A(_0489_),
    .B(_0491_),
    .C(net399),
    .Y(_0114_));
 sg13g2_nand2_1 _1179_ (.Y(_0493_),
    .A(net404),
    .B(_0491_));
 sg13g2_xnor2_1 _1180_ (.Y(_0494_),
    .A(net404),
    .B(_0491_));
 sg13g2_nor2_1 _1181_ (.A(_0489_),
    .B(net405),
    .Y(_0115_));
 sg13g2_xor2_1 _1182_ (.B(_0493_),
    .A(net432),
    .X(_0495_));
 sg13g2_nor2_1 _1183_ (.A(_0489_),
    .B(_0495_),
    .Y(_0116_));
 sg13g2_nand2_1 _1184_ (.Y(_0496_),
    .A(\ltc.sec_u[3] ),
    .B(\ltc.sec_u[1] ));
 sg13g2_nor3_1 _1185_ (.A(net410),
    .B(\ltc.sec_u[0] ),
    .C(_0496_),
    .Y(_0497_));
 sg13g2_and2_1 _1186_ (.A(net346),
    .B(_0497_),
    .X(_0498_));
 sg13g2_nand2_1 _1187_ (.Y(_0499_),
    .A(net178),
    .B(_0487_));
 sg13g2_nor2_1 _1188_ (.A(net346),
    .B(_0497_),
    .Y(_0500_));
 sg13g2_nor3_1 _1189_ (.A(_0498_),
    .B(_0499_),
    .C(net347),
    .Y(_0117_));
 sg13g2_nor2_1 _1190_ (.A(net402),
    .B(_0498_),
    .Y(_0501_));
 sg13g2_and2_1 _1191_ (.A(net402),
    .B(_0498_),
    .X(_0502_));
 sg13g2_nor3_1 _1192_ (.A(_0499_),
    .B(net403),
    .C(_0502_),
    .Y(_0118_));
 sg13g2_xnor2_1 _1193_ (.Y(_0503_),
    .A(net395),
    .B(_0502_));
 sg13g2_nor2_1 _1194_ (.A(_0499_),
    .B(net396),
    .Y(_0119_));
 sg13g2_nor2_1 _1195_ (.A(net428),
    .B(net328),
    .Y(_0504_));
 sg13g2_nor2b_1 _1196_ (.A(\ltc.frm_u[1] ),
    .B_N(\ltc.frm_u[0] ),
    .Y(_0505_));
 sg13g2_a22oi_1 _1197_ (.Y(_0506_),
    .B1(_0505_),
    .B2(_0207_),
    .A2(_0504_),
    .A1(_0333_));
 sg13g2_nand2_1 _1198_ (.Y(_0507_),
    .A(\ltc.frm_u[2] ),
    .B(_0147_));
 sg13g2_nand4_1 _1199_ (.B(\ltc.frm_d[0] ),
    .C(_0334_),
    .A(_0145_),
    .Y(_0508_),
    .D(_0504_));
 sg13g2_o21ai_1 _1200_ (.B1(_0508_),
    .Y(_0509_),
    .A1(_0506_),
    .A2(_0507_));
 sg13g2_nand3_1 _1201_ (.B(net407),
    .C(_0509_),
    .A(_0144_),
    .Y(_0510_));
 sg13g2_nor2_1 _1202_ (.A(_0148_),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_nand2b_2 _1203_ (.Y(_0512_),
    .B(net178),
    .A_N(_0497_));
 sg13g2_a21oi_1 _1204_ (.A1(_0148_),
    .A2(_0510_),
    .Y(_0513_),
    .B1(_0512_));
 sg13g2_nor2b_1 _1205_ (.A(_0511_),
    .B_N(_0513_),
    .Y(_0120_));
 sg13g2_nor2_1 _1206_ (.A(net424),
    .B(_0511_),
    .Y(_0514_));
 sg13g2_and2_1 _1207_ (.A(net424),
    .B(_0511_),
    .X(_0515_));
 sg13g2_nor3_1 _1208_ (.A(_0512_),
    .B(net425),
    .C(_0515_),
    .Y(_0121_));
 sg13g2_nand2_1 _1209_ (.Y(_0516_),
    .A(net410),
    .B(_0515_));
 sg13g2_xnor2_1 _1210_ (.Y(_0517_),
    .A(net410),
    .B(_0515_));
 sg13g2_nor2_1 _1211_ (.A(_0512_),
    .B(net411),
    .Y(_0122_));
 sg13g2_xor2_1 _1212_ (.B(_0516_),
    .A(net435),
    .X(_0518_));
 sg13g2_nor2_1 _1213_ (.A(_0512_),
    .B(_0518_),
    .Y(_0123_));
 sg13g2_nand2_1 _1214_ (.Y(_0519_),
    .A(net179),
    .B(_0510_));
 sg13g2_nand4_1 _1215_ (.B(_0145_),
    .C(net428),
    .A(net445),
    .Y(_0520_),
    .D(_0146_));
 sg13g2_and2_1 _1216_ (.A(_0147_),
    .B(_0520_),
    .X(_0521_));
 sg13g2_nor2_1 _1217_ (.A(_0147_),
    .B(_0520_),
    .Y(_0522_));
 sg13g2_nor3_1 _1218_ (.A(_0519_),
    .B(net470),
    .C(_0522_),
    .Y(_0124_));
 sg13g2_xnor2_1 _1219_ (.Y(_0523_),
    .A(net407),
    .B(_0522_));
 sg13g2_nor2_1 _1220_ (.A(_0519_),
    .B(net408),
    .Y(_0125_));
 sg13g2_nand3_1 _1221_ (.B(_0510_),
    .C(_0520_),
    .A(net128),
    .Y(_0524_));
 sg13g2_o21ai_1 _1222_ (.B1(net180),
    .Y(_0525_),
    .A1(net328),
    .A2(_0451_));
 sg13g2_a21oi_1 _1223_ (.A1(net328),
    .A2(_0524_),
    .Y(_0126_),
    .B1(_0525_));
 sg13g2_nand4_1 _1224_ (.B(net128),
    .C(_0510_),
    .A(net428),
    .Y(_0526_),
    .D(_0520_));
 sg13g2_nand2_1 _1225_ (.Y(_0527_),
    .A(net428),
    .B(net328));
 sg13g2_nand3b_1 _1226_ (.B(_0527_),
    .C(_0451_),
    .Y(_0528_),
    .A_N(_0504_));
 sg13g2_a21oi_1 _1227_ (.A1(_0526_),
    .A2(_0528_),
    .Y(_0127_),
    .B1(net173));
 sg13g2_nand4_1 _1228_ (.B(net128),
    .C(_0510_),
    .A(net413),
    .Y(_0529_),
    .D(_0520_));
 sg13g2_nand2_1 _1229_ (.Y(_0530_),
    .A(_0145_),
    .B(_0527_));
 sg13g2_nand3_1 _1230_ (.B(net428),
    .C(net328),
    .A(net413),
    .Y(_0531_));
 sg13g2_nand2_1 _1231_ (.Y(_0532_),
    .A(_0451_),
    .B(_0531_));
 sg13g2_nand3_1 _1232_ (.B(_0530_),
    .C(_0531_),
    .A(_0451_),
    .Y(_0533_));
 sg13g2_a21oi_1 _1233_ (.A1(_0529_),
    .A2(_0533_),
    .Y(_0128_),
    .B1(net173));
 sg13g2_a21oi_1 _1234_ (.A1(net128),
    .A2(_0520_),
    .Y(_0534_),
    .B1(_0144_));
 sg13g2_or2_1 _1235_ (.X(_0535_),
    .B(_0531_),
    .A(net128));
 sg13g2_a221oi_1 _1236_ (.B2(_0144_),
    .C1(net173),
    .B1(_0535_),
    .A1(_0532_),
    .Y(_0129_),
    .A2(_0534_));
 sg13g2_nor2_1 _1237_ (.A(\ltc.bit_clk ),
    .B(\ltc.output_buffer[79] ),
    .Y(_0536_));
 sg13g2_nor2_1 _1238_ (.A(_0177_),
    .B(_0536_),
    .Y(_0537_));
 sg13g2_o21ai_1 _1239_ (.B1(net181),
    .Y(_0538_),
    .A1(net228),
    .A2(_0537_));
 sg13g2_a21oi_1 _1240_ (.A1(net228),
    .A2(_0537_),
    .Y(_0130_),
    .B1(_0538_));
 sg13g2_and2_1 _1241_ (.A(net361),
    .B(net227),
    .X(_0539_));
 sg13g2_and4_1 _1242_ (.A(net267),
    .B(\ltc.bit_counter[2] ),
    .C(net361),
    .D(net227),
    .X(_0540_));
 sg13g2_nand2_1 _1243_ (.Y(_0541_),
    .A(\ltc.bit_counter[5] ),
    .B(\ltc.bit_counter[4] ));
 sg13g2_and3_2 _1244_ (.X(_0542_),
    .A(net277),
    .B(net437),
    .C(_0540_));
 sg13g2_and3_1 _1245_ (.X(_0543_),
    .A(\ltc.bit_counter[6] ),
    .B(net261),
    .C(_0542_));
 sg13g2_and4_1 _1246_ (.A(\ltc.bit_counter[6] ),
    .B(net261),
    .C(net385),
    .D(_0542_),
    .X(_0544_));
 sg13g2_nand3_1 _1247_ (.B(net462),
    .C(_0544_),
    .A(net440),
    .Y(_0545_));
 sg13g2_xor2_1 _1248_ (.B(_0545_),
    .A(net446),
    .X(_0546_));
 sg13g2_a21o_1 _1249_ (.A2(_0544_),
    .A1(net440),
    .B1(net462),
    .X(_0547_));
 sg13g2_nand2_1 _1250_ (.Y(_0548_),
    .A(_0545_),
    .B(_0547_));
 sg13g2_nand3_1 _1251_ (.B(\ltc.bit_counter[9] ),
    .C(_0207_),
    .A(\ltc.bit_counter[2] ),
    .Y(_0549_));
 sg13g2_nor3_1 _1252_ (.A(\ltc.bit_counter[6] ),
    .B(_0541_),
    .C(_0549_),
    .Y(_0550_));
 sg13g2_nor3_1 _1253_ (.A(\ltc.bit_counter[2] ),
    .B(_0154_),
    .C(\ltc.bit_counter[9] ),
    .Y(_0551_));
 sg13g2_and2_1 _1254_ (.A(_0173_),
    .B(_0334_),
    .X(_0552_));
 sg13g2_a21oi_1 _1255_ (.A1(_0551_),
    .A2(_0552_),
    .Y(_0553_),
    .B1(_0550_));
 sg13g2_nand3_1 _1256_ (.B(\ltc.bit_counter[8] ),
    .C(_0539_),
    .A(\ltc.bit_counter[7] ),
    .Y(_0554_));
 sg13g2_nor3_1 _1257_ (.A(\ltc.bit_counter[3] ),
    .B(_0553_),
    .C(_0554_),
    .Y(_0555_));
 sg13g2_xnor2_1 _1258_ (.Y(_0556_),
    .A(net457),
    .B(_0539_));
 sg13g2_nand3_1 _1259_ (.B(_0175_),
    .C(_0333_),
    .A(_0174_),
    .Y(_0557_));
 sg13g2_nor4_1 _1260_ (.A(\ltc.bit_counter[3] ),
    .B(_0541_),
    .C(_0556_),
    .D(_0557_),
    .Y(_0558_));
 sg13g2_mux2_1 _1261_ (.A0(_0558_),
    .A1(_0555_),
    .S(_0548_),
    .X(_0559_));
 sg13g2_nor2b_1 _1262_ (.A(_0546_),
    .B_N(_0559_),
    .Y(_0560_));
 sg13g2_nand2b_1 _1263_ (.Y(_0561_),
    .B(net178),
    .A_N(_0560_));
 sg13g2_nor2_1 _1264_ (.A(net227),
    .B(net124),
    .Y(_0131_));
 sg13g2_nor3_1 _1265_ (.A(_0171_),
    .B(_0539_),
    .C(net123),
    .Y(_0132_));
 sg13g2_nor2_1 _1266_ (.A(_0556_),
    .B(net123),
    .Y(_0133_));
 sg13g2_a21oi_1 _1267_ (.A1(\ltc.bit_counter[2] ),
    .A2(_0539_),
    .Y(_0562_),
    .B1(net267));
 sg13g2_nor3_1 _1268_ (.A(_0540_),
    .B(net123),
    .C(net268),
    .Y(_0134_));
 sg13g2_xnor2_1 _1269_ (.Y(_0563_),
    .A(net437),
    .B(_0540_));
 sg13g2_nor2_1 _1270_ (.A(net124),
    .B(net438),
    .Y(_0135_));
 sg13g2_a21oi_1 _1271_ (.A1(\ltc.bit_counter[4] ),
    .A2(_0540_),
    .Y(_0564_),
    .B1(net277));
 sg13g2_nor3_1 _1272_ (.A(_0542_),
    .B(net123),
    .C(net278),
    .Y(_0136_));
 sg13g2_xnor2_1 _1273_ (.Y(_0565_),
    .A(net442),
    .B(_0542_));
 sg13g2_nor2_1 _1274_ (.A(net124),
    .B(_0565_),
    .Y(_0137_));
 sg13g2_a21oi_1 _1275_ (.A1(\ltc.bit_counter[6] ),
    .A2(_0542_),
    .Y(_0566_),
    .B1(net261));
 sg13g2_nor3_1 _1276_ (.A(_0543_),
    .B(net124),
    .C(net262),
    .Y(_0138_));
 sg13g2_nor2_1 _1277_ (.A(net385),
    .B(_0543_),
    .Y(_0567_));
 sg13g2_nor3_1 _1278_ (.A(_0544_),
    .B(net123),
    .C(net386),
    .Y(_0139_));
 sg13g2_xnor2_1 _1279_ (.Y(_0568_),
    .A(net440),
    .B(_0544_));
 sg13g2_nor2_1 _1280_ (.A(net123),
    .B(net441),
    .Y(_0140_));
 sg13g2_nor2_1 _1281_ (.A(_0548_),
    .B(net123),
    .Y(_0141_));
 sg13g2_nor2_1 _1282_ (.A(net447),
    .B(net123),
    .Y(_0142_));
 sg13g2_o21ai_1 _1283_ (.B1(net181),
    .Y(_0569_),
    .A1(net231),
    .A2(_0560_));
 sg13g2_a21oi_1 _1284_ (.A1(net231),
    .A2(_0560_),
    .Y(_0143_),
    .B1(_0569_));
 sg13g2_dfrbpq_1 _1285_ (.RESET_B(net105),
    .D(_0000_),
    .Q(\ltc.output_buffer[0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1286_ (.RESET_B(net89),
    .D(_0001_),
    .Q(\ltc.output_buffer[1] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1287_ (.RESET_B(net88),
    .D(_0002_),
    .Q(\ltc.output_buffer[2] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1288_ (.RESET_B(net87),
    .D(_0003_),
    .Q(\ltc.output_buffer[3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1289_ (.RESET_B(net86),
    .D(net248),
    .Q(\ltc.output_buffer[4] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1290_ (.RESET_B(net85),
    .D(_0005_),
    .Q(\ltc.output_buffer[5] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1291_ (.RESET_B(net84),
    .D(net234),
    .Q(\ltc.output_buffer[6] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1292_ (.RESET_B(net83),
    .D(_0007_),
    .Q(\ltc.output_buffer[7] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1293_ (.RESET_B(net82),
    .D(net238),
    .Q(\ltc.output_buffer[8] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1294_ (.RESET_B(net81),
    .D(_0009_),
    .Q(\ltc.output_buffer[9] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1295_ (.RESET_B(net80),
    .D(net246),
    .Q(\ltc.output_buffer[10] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1296_ (.RESET_B(net79),
    .D(net244),
    .Q(\ltc.output_buffer[11] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1297_ (.RESET_B(net78),
    .D(_0012_),
    .Q(\ltc.output_buffer[12] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1298_ (.RESET_B(net77),
    .D(net254),
    .Q(\ltc.output_buffer[13] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1299_ (.RESET_B(net76),
    .D(_0014_),
    .Q(\ltc.output_buffer[14] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1300_ (.RESET_B(net75),
    .D(_0015_),
    .Q(\ltc.output_buffer[15] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1301_ (.RESET_B(net74),
    .D(_0016_),
    .Q(\ltc.output_buffer[16] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1302_ (.RESET_B(net73),
    .D(_0017_),
    .Q(\ltc.output_buffer[17] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1303_ (.RESET_B(net72),
    .D(_0018_),
    .Q(\ltc.output_buffer[18] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1304_ (.RESET_B(net71),
    .D(_0019_),
    .Q(\ltc.output_buffer[19] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1305_ (.RESET_B(net70),
    .D(net283),
    .Q(\ltc.output_buffer[20] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1306_ (.RESET_B(net69),
    .D(_0021_),
    .Q(\ltc.output_buffer[21] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1307_ (.RESET_B(net68),
    .D(_0022_),
    .Q(\ltc.output_buffer[22] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _1308_ (.RESET_B(net67),
    .D(net296),
    .Q(\ltc.output_buffer[23] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1309_ (.RESET_B(net66),
    .D(_0024_),
    .Q(\ltc.output_buffer[24] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1310_ (.RESET_B(net65),
    .D(_0025_),
    .Q(\ltc.output_buffer[25] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1311_ (.RESET_B(net64),
    .D(_0026_),
    .Q(\ltc.output_buffer[26] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1312_ (.RESET_B(net63),
    .D(_0027_),
    .Q(\ltc.output_buffer[27] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1313_ (.RESET_B(net62),
    .D(net290),
    .Q(\ltc.output_buffer[28] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1314_ (.RESET_B(net61),
    .D(net294),
    .Q(\ltc.output_buffer[29] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1315_ (.RESET_B(net60),
    .D(net336),
    .Q(\ltc.output_buffer[30] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1316_ (.RESET_B(net59),
    .D(net332),
    .Q(\ltc.output_buffer[31] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1317_ (.RESET_B(net58),
    .D(_0032_),
    .Q(\ltc.output_buffer[32] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1318_ (.RESET_B(net57),
    .D(_0033_),
    .Q(\ltc.output_buffer[33] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1319_ (.RESET_B(net56),
    .D(_0034_),
    .Q(\ltc.output_buffer[34] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1320_ (.RESET_B(net55),
    .D(_0035_),
    .Q(\ltc.output_buffer[35] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1321_ (.RESET_B(net54),
    .D(_0036_),
    .Q(\ltc.output_buffer[36] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1322_ (.RESET_B(net53),
    .D(net292),
    .Q(\ltc.output_buffer[37] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1323_ (.RESET_B(net52),
    .D(net302),
    .Q(\ltc.output_buffer[38] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1324_ (.RESET_B(net51),
    .D(net308),
    .Q(\ltc.output_buffer[39] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1325_ (.RESET_B(net50),
    .D(_0040_),
    .Q(\ltc.output_buffer[40] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1326_ (.RESET_B(net49),
    .D(_0041_),
    .Q(\ltc.output_buffer[41] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1327_ (.RESET_B(net48),
    .D(_0042_),
    .Q(\ltc.output_buffer[42] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1328_ (.RESET_B(net47),
    .D(_0043_),
    .Q(\ltc.output_buffer[43] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1329_ (.RESET_B(net46),
    .D(net373),
    .Q(\ltc.output_buffer[44] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1330_ (.RESET_B(net45),
    .D(net352),
    .Q(\ltc.output_buffer[45] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1331_ (.RESET_B(net44),
    .D(net300),
    .Q(\ltc.output_buffer[46] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1332_ (.RESET_B(net43),
    .D(net287),
    .Q(\ltc.output_buffer[47] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1333_ (.RESET_B(net42),
    .D(_0048_),
    .Q(\ltc.output_buffer[48] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1334_ (.RESET_B(net41),
    .D(_0049_),
    .Q(\ltc.output_buffer[49] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1335_ (.RESET_B(net40),
    .D(_0050_),
    .Q(\ltc.output_buffer[50] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1336_ (.RESET_B(net39),
    .D(_0051_),
    .Q(\ltc.output_buffer[51] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1337_ (.RESET_B(net38),
    .D(net271),
    .Q(\ltc.output_buffer[52] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1338_ (.RESET_B(net37),
    .D(net304),
    .Q(\ltc.output_buffer[53] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1339_ (.RESET_B(net36),
    .D(net273),
    .Q(\ltc.output_buffer[54] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1340_ (.RESET_B(net35),
    .D(net266),
    .Q(\ltc.output_buffer[55] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1341_ (.RESET_B(net34),
    .D(_0056_),
    .Q(\ltc.output_buffer[56] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1342_ (.RESET_B(net33),
    .D(_0057_),
    .Q(\ltc.output_buffer[57] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1343_ (.RESET_B(net32),
    .D(_0058_),
    .Q(\ltc.output_buffer[58] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1344_ (.RESET_B(net31),
    .D(_0059_),
    .Q(\ltc.output_buffer[59] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1345_ (.RESET_B(net30),
    .D(net367),
    .Q(\ltc.output_buffer[60] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1346_ (.RESET_B(net29),
    .D(net281),
    .Q(\ltc.output_buffer[61] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1347_ (.RESET_B(net28),
    .D(net306),
    .Q(\ltc.output_buffer[62] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _1348_ (.RESET_B(net27),
    .D(net285),
    .Q(\ltc.output_buffer[63] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1349_ (.RESET_B(net26),
    .D(_0064_),
    .Q(\ltc.output_buffer[64] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1350_ (.RESET_B(net25),
    .D(_0065_),
    .Q(\ltc.output_buffer[65] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1351_ (.RESET_B(net24),
    .D(_0066_),
    .Q(\ltc.output_buffer[66] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1352_ (.RESET_B(net23),
    .D(_0067_),
    .Q(\ltc.output_buffer[67] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1353_ (.RESET_B(net225),
    .D(_0068_),
    .Q(\ltc.output_buffer[68] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1354_ (.RESET_B(net224),
    .D(_0069_),
    .Q(\ltc.output_buffer[69] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net223),
    .D(net323),
    .Q(\ltc.output_buffer[70] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1356_ (.RESET_B(net222),
    .D(net363),
    .Q(\ltc.output_buffer[71] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net221),
    .D(_0072_),
    .Q(\ltc.output_buffer[72] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1358_ (.RESET_B(net220),
    .D(_0073_),
    .Q(\ltc.output_buffer[73] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1359_ (.RESET_B(net219),
    .D(_0074_),
    .Q(\ltc.output_buffer[74] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1360_ (.RESET_B(net218),
    .D(_0075_),
    .Q(\ltc.output_buffer[75] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1361_ (.RESET_B(net217),
    .D(net298),
    .Q(\ltc.output_buffer[76] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net216),
    .D(net379),
    .Q(\ltc.output_buffer[77] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net215),
    .D(net314),
    .Q(\ltc.output_buffer[78] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1364_ (.RESET_B(net214),
    .D(net359),
    .Q(\ltc.output_buffer[79] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1365_ (.RESET_B(net213),
    .D(_0080_),
    .Q(\ltc.hrs_u[0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1366_ (.RESET_B(net211),
    .D(_0081_),
    .Q(\ltc.frm_counter[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1367_ (.RESET_B(net210),
    .D(_0082_),
    .Q(\ltc.frm_counter[1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1368_ (.RESET_B(net209),
    .D(net276),
    .Q(\ltc.frm_counter[2] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1369_ (.RESET_B(net208),
    .D(_0084_),
    .Q(\ltc.frm_counter[3] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1370_ (.RESET_B(net207),
    .D(_0085_),
    .Q(\ltc.frm_counter[4] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1371_ (.RESET_B(net206),
    .D(net418),
    .Q(\ltc.frm_counter[5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1372_ (.RESET_B(net205),
    .D(_0087_),
    .Q(\ltc.frm_counter[6] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1373_ (.RESET_B(net204),
    .D(_0088_),
    .Q(\ltc.frm_counter[7] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1374_ (.RESET_B(net203),
    .D(_0089_),
    .Q(\ltc.frm_counter[8] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1375_ (.RESET_B(net202),
    .D(_0090_),
    .Q(\ltc.frm_counter[9] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1376_ (.RESET_B(net201),
    .D(_0091_),
    .Q(\ltc.frm_counter[10] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1377_ (.RESET_B(net200),
    .D(net421),
    .Q(\ltc.frm_counter[11] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1378_ (.RESET_B(net199),
    .D(_0093_),
    .Q(\ltc.frm_counter[12] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1379_ (.RESET_B(net198),
    .D(net461),
    .Q(\ltc.frm_counter[13] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1380_ (.RESET_B(net197),
    .D(_0095_),
    .Q(\ltc.frm_counter[14] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1381_ (.RESET_B(net196),
    .D(_0096_),
    .Q(\ltc.frm_counter[15] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1382_ (.RESET_B(net195),
    .D(_0097_),
    .Q(\ltc.frm_counter[16] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1383_ (.RESET_B(net194),
    .D(_0098_),
    .Q(\ltc.frm_counter[17] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1384_ (.RESET_B(net193),
    .D(_0099_),
    .Q(\ltc.frm_counter[18] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net192),
    .D(net259),
    .Q(\ltc.frm_counter[19] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1386_ (.RESET_B(net191),
    .D(_0101_),
    .Q(\ltc.frm_counter[20] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net190),
    .D(net241),
    .Q(\ltc.frm_counter[21] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1388_ (.RESET_B(net189),
    .D(net357),
    .Q(\ltc.frm_counter[22] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net188),
    .D(_0104_),
    .Q(\ltc.frm_counter[23] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1390_ (.RESET_B(net187),
    .D(net431),
    .Q(\ltc.hrs_d[0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net185),
    .D(_0106_),
    .Q(\ltc.hrs_d[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1392_ (.RESET_B(net183),
    .D(_0107_),
    .Q(\ltc.hrs_u[1] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1393_ (.RESET_B(net122),
    .D(_0108_),
    .Q(\ltc.hrs_u[2] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1394_ (.RESET_B(net120),
    .D(_0109_),
    .Q(\ltc.hrs_u[3] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1395_ (.RESET_B(net118),
    .D(net319),
    .Q(\ltc.min_d[0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1396_ (.RESET_B(net116),
    .D(_0111_),
    .Q(\ltc.min_d[1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1397_ (.RESET_B(net114),
    .D(net382),
    .Q(\ltc.min_d[2] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net112),
    .D(_0113_),
    .Q(\ltc.min_u[0] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1399_ (.RESET_B(net110),
    .D(_0114_),
    .Q(\ltc.min_u[1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1400_ (.RESET_B(net108),
    .D(net406),
    .Q(\ltc.min_u[2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1401_ (.RESET_B(net106),
    .D(net433),
    .Q(\ltc.min_u[3] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net104),
    .D(net348),
    .Q(\ltc.sec_d[0] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1403_ (.RESET_B(net102),
    .D(_0118_),
    .Q(\ltc.sec_d[1] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net100),
    .D(net397),
    .Q(\ltc.sec_d[2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1405_ (.RESET_B(net98),
    .D(_0120_),
    .Q(\ltc.sec_u[0] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net96),
    .D(_0121_),
    .Q(\ltc.sec_u[1] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1407_ (.RESET_B(net94),
    .D(net412),
    .Q(\ltc.sec_u[2] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1408_ (.RESET_B(net92),
    .D(net436),
    .Q(\ltc.sec_u[3] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1409_ (.RESET_B(net90),
    .D(net471),
    .Q(\ltc.frm_d[0] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1410_ (.RESET_B(net186),
    .D(_0125_),
    .Q(\ltc.frm_d[1] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1411_ (.RESET_B(net182),
    .D(_0126_),
    .Q(\ltc.frm_u[0] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _1412_ (.RESET_B(net119),
    .D(_0127_),
    .Q(\ltc.frm_u[1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1413_ (.RESET_B(net115),
    .D(net414),
    .Q(\ltc.frm_u[2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1414_ (.RESET_B(net111),
    .D(_0129_),
    .Q(\ltc.frm_u[3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net107),
    .D(net229),
    .Q(\ltc.timecode ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1416_ (.RESET_B(net103),
    .D(_0131_),
    .Q(\ltc.bit_counter[0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net101),
    .D(_0132_),
    .Q(\ltc.bit_counter[1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1418_ (.RESET_B(net99),
    .D(_0133_),
    .Q(\ltc.bit_counter[2] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1419_ (.RESET_B(net97),
    .D(net269),
    .Q(\ltc.bit_counter[3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1420_ (.RESET_B(net95),
    .D(_0135_),
    .Q(\ltc.bit_counter[4] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1421_ (.RESET_B(net93),
    .D(net279),
    .Q(\ltc.bit_counter[5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1422_ (.RESET_B(net91),
    .D(_0137_),
    .Q(\ltc.bit_counter[6] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1423_ (.RESET_B(net212),
    .D(net263),
    .Q(\ltc.bit_counter[7] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net184),
    .D(net387),
    .Q(\ltc.bit_counter[8] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1425_ (.RESET_B(net121),
    .D(_0140_),
    .Q(\ltc.bit_counter[9] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net117),
    .D(_0141_),
    .Q(\ltc.bit_counter[10] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net113),
    .D(_0142_),
    .Q(\ltc.bit_counter[11] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net109),
    .D(net232),
    .Q(\ltc.bit_clk ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_tiehi _1351__24 (.L_HI(net24));
 sg13g2_tiehi _1350__25 (.L_HI(net25));
 sg13g2_tiehi _1349__26 (.L_HI(net26));
 sg13g2_tiehi _1348__27 (.L_HI(net27));
 sg13g2_tiehi _1347__28 (.L_HI(net28));
 sg13g2_tiehi _1346__29 (.L_HI(net29));
 sg13g2_tiehi _1345__30 (.L_HI(net30));
 sg13g2_tiehi _1344__31 (.L_HI(net31));
 sg13g2_tiehi _1343__32 (.L_HI(net32));
 sg13g2_tiehi _1342__33 (.L_HI(net33));
 sg13g2_tiehi _1341__34 (.L_HI(net34));
 sg13g2_tiehi _1340__35 (.L_HI(net35));
 sg13g2_tiehi _1339__36 (.L_HI(net36));
 sg13g2_tiehi _1338__37 (.L_HI(net37));
 sg13g2_tiehi _1337__38 (.L_HI(net38));
 sg13g2_tiehi _1336__39 (.L_HI(net39));
 sg13g2_tiehi _1335__40 (.L_HI(net40));
 sg13g2_tiehi _1334__41 (.L_HI(net41));
 sg13g2_tiehi _1333__42 (.L_HI(net42));
 sg13g2_tiehi _1332__43 (.L_HI(net43));
 sg13g2_tiehi _1331__44 (.L_HI(net44));
 sg13g2_tiehi _1330__45 (.L_HI(net45));
 sg13g2_tiehi _1329__46 (.L_HI(net46));
 sg13g2_tiehi _1328__47 (.L_HI(net47));
 sg13g2_tiehi _1327__48 (.L_HI(net48));
 sg13g2_tiehi _1326__49 (.L_HI(net49));
 sg13g2_tiehi _1325__50 (.L_HI(net50));
 sg13g2_tiehi _1324__51 (.L_HI(net51));
 sg13g2_tiehi _1323__52 (.L_HI(net52));
 sg13g2_tiehi _1322__53 (.L_HI(net53));
 sg13g2_tiehi _1321__54 (.L_HI(net54));
 sg13g2_tiehi _1320__55 (.L_HI(net55));
 sg13g2_tiehi _1319__56 (.L_HI(net56));
 sg13g2_tiehi _1318__57 (.L_HI(net57));
 sg13g2_tiehi _1317__58 (.L_HI(net58));
 sg13g2_tiehi _1316__59 (.L_HI(net59));
 sg13g2_tiehi _1315__60 (.L_HI(net60));
 sg13g2_tiehi _1314__61 (.L_HI(net61));
 sg13g2_tiehi _1313__62 (.L_HI(net62));
 sg13g2_tiehi _1312__63 (.L_HI(net63));
 sg13g2_tiehi _1311__64 (.L_HI(net64));
 sg13g2_tiehi _1310__65 (.L_HI(net65));
 sg13g2_tiehi _1309__66 (.L_HI(net66));
 sg13g2_tiehi _1308__67 (.L_HI(net67));
 sg13g2_tiehi _1307__68 (.L_HI(net68));
 sg13g2_tiehi _1306__69 (.L_HI(net69));
 sg13g2_tiehi _1305__70 (.L_HI(net70));
 sg13g2_tiehi _1304__71 (.L_HI(net71));
 sg13g2_tiehi _1303__72 (.L_HI(net72));
 sg13g2_tiehi _1302__73 (.L_HI(net73));
 sg13g2_tiehi _1301__74 (.L_HI(net74));
 sg13g2_tiehi _1300__75 (.L_HI(net75));
 sg13g2_tiehi _1299__76 (.L_HI(net76));
 sg13g2_tiehi _1298__77 (.L_HI(net77));
 sg13g2_tiehi _1297__78 (.L_HI(net78));
 sg13g2_tiehi _1296__79 (.L_HI(net79));
 sg13g2_tiehi _1295__80 (.L_HI(net80));
 sg13g2_tiehi _1294__81 (.L_HI(net81));
 sg13g2_tiehi _1293__82 (.L_HI(net82));
 sg13g2_tiehi _1292__83 (.L_HI(net83));
 sg13g2_tiehi _1291__84 (.L_HI(net84));
 sg13g2_tiehi _1290__85 (.L_HI(net85));
 sg13g2_tiehi _1289__86 (.L_HI(net86));
 sg13g2_tiehi _1288__87 (.L_HI(net87));
 sg13g2_tiehi _1287__88 (.L_HI(net88));
 sg13g2_tiehi _1286__89 (.L_HI(net89));
 sg13g2_tiehi _1409__90 (.L_HI(net90));
 sg13g2_tiehi _1422__91 (.L_HI(net91));
 sg13g2_tiehi _1408__92 (.L_HI(net92));
 sg13g2_tiehi _1421__93 (.L_HI(net93));
 sg13g2_tiehi _1407__94 (.L_HI(net94));
 sg13g2_tiehi _1420__95 (.L_HI(net95));
 sg13g2_tiehi _1406__96 (.L_HI(net96));
 sg13g2_tiehi _1419__97 (.L_HI(net97));
 sg13g2_tiehi _1405__98 (.L_HI(net98));
 sg13g2_tiehi _1418__99 (.L_HI(net99));
 sg13g2_tiehi _1404__100 (.L_HI(net100));
 sg13g2_tiehi _1417__101 (.L_HI(net101));
 sg13g2_tiehi _1403__102 (.L_HI(net102));
 sg13g2_tiehi _1416__103 (.L_HI(net103));
 sg13g2_tiehi _1402__104 (.L_HI(net104));
 sg13g2_tiehi _1285__105 (.L_HI(net105));
 sg13g2_tiehi _1401__106 (.L_HI(net106));
 sg13g2_tiehi _1415__107 (.L_HI(net107));
 sg13g2_tiehi _1400__108 (.L_HI(net108));
 sg13g2_tiehi _1428__109 (.L_HI(net109));
 sg13g2_tiehi _1399__110 (.L_HI(net110));
 sg13g2_tiehi _1414__111 (.L_HI(net111));
 sg13g2_tiehi _1398__112 (.L_HI(net112));
 sg13g2_tiehi _1427__113 (.L_HI(net113));
 sg13g2_tiehi _1397__114 (.L_HI(net114));
 sg13g2_tiehi _1413__115 (.L_HI(net115));
 sg13g2_tiehi _1396__116 (.L_HI(net116));
 sg13g2_tiehi _1426__117 (.L_HI(net117));
 sg13g2_tiehi _1395__118 (.L_HI(net118));
 sg13g2_tiehi _1412__119 (.L_HI(net119));
 sg13g2_tiehi _1394__120 (.L_HI(net120));
 sg13g2_tiehi _1425__121 (.L_HI(net121));
 sg13g2_tiehi _1393__122 (.L_HI(net122));
 sg13g2_tiehi _1411__123 (.L_HI(net182));
 sg13g2_tiehi _1392__124 (.L_HI(net183));
 sg13g2_tiehi _1424__125 (.L_HI(net184));
 sg13g2_tiehi _1391__126 (.L_HI(net185));
 sg13g2_tiehi _1410__127 (.L_HI(net186));
 sg13g2_tiehi _1390__128 (.L_HI(net187));
 sg13g2_tiehi _1389__129 (.L_HI(net188));
 sg13g2_tiehi _1388__130 (.L_HI(net189));
 sg13g2_tiehi _1387__131 (.L_HI(net190));
 sg13g2_tiehi _1386__132 (.L_HI(net191));
 sg13g2_tiehi _1385__133 (.L_HI(net192));
 sg13g2_tiehi _1384__134 (.L_HI(net193));
 sg13g2_tiehi _1383__135 (.L_HI(net194));
 sg13g2_tiehi _1382__136 (.L_HI(net195));
 sg13g2_tiehi _1381__137 (.L_HI(net196));
 sg13g2_tiehi _1380__138 (.L_HI(net197));
 sg13g2_tiehi _1379__139 (.L_HI(net198));
 sg13g2_tiehi _1378__140 (.L_HI(net199));
 sg13g2_tiehi _1377__141 (.L_HI(net200));
 sg13g2_tiehi _1376__142 (.L_HI(net201));
 sg13g2_tiehi _1375__143 (.L_HI(net202));
 sg13g2_tiehi _1374__144 (.L_HI(net203));
 sg13g2_tiehi _1373__145 (.L_HI(net204));
 sg13g2_tiehi _1372__146 (.L_HI(net205));
 sg13g2_tiehi _1371__147 (.L_HI(net206));
 sg13g2_tiehi _1370__148 (.L_HI(net207));
 sg13g2_tiehi _1369__149 (.L_HI(net208));
 sg13g2_tiehi _1368__150 (.L_HI(net209));
 sg13g2_tiehi _1367__151 (.L_HI(net210));
 sg13g2_tiehi _1366__152 (.L_HI(net211));
 sg13g2_tiehi _1423__153 (.L_HI(net212));
 sg13g2_tiehi _1365__154 (.L_HI(net213));
 sg13g2_tiehi _1364__155 (.L_HI(net214));
 sg13g2_tiehi _1363__156 (.L_HI(net215));
 sg13g2_tiehi _1362__157 (.L_HI(net216));
 sg13g2_tiehi _1361__158 (.L_HI(net217));
 sg13g2_tiehi _1360__159 (.L_HI(net218));
 sg13g2_tiehi _1359__160 (.L_HI(net219));
 sg13g2_tiehi _1358__161 (.L_HI(net220));
 sg13g2_tiehi _1357__162 (.L_HI(net221));
 sg13g2_tiehi _1356__163 (.L_HI(net222));
 sg13g2_tiehi _1355__164 (.L_HI(net223));
 sg13g2_tiehi _1354__165 (.L_HI(net224));
 sg13g2_tiehi _1353__166 (.L_HI(net225));
 sg13g2_tiehi tt_um_flummer_ltc_167 (.L_HI(net226));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_flummer_ltc_10 (.L_LO(net10));
 sg13g2_tielo tt_um_flummer_ltc_11 (.L_LO(net11));
 sg13g2_tielo tt_um_flummer_ltc_12 (.L_LO(net12));
 sg13g2_tielo tt_um_flummer_ltc_13 (.L_LO(net13));
 sg13g2_tielo tt_um_flummer_ltc_14 (.L_LO(net14));
 sg13g2_tielo tt_um_flummer_ltc_15 (.L_LO(net15));
 sg13g2_tielo tt_um_flummer_ltc_16 (.L_LO(net16));
 sg13g2_tielo tt_um_flummer_ltc_17 (.L_LO(net17));
 sg13g2_tielo tt_um_flummer_ltc_18 (.L_LO(net18));
 sg13g2_tielo tt_um_flummer_ltc_19 (.L_LO(net19));
 sg13g2_tielo tt_um_flummer_ltc_20 (.L_LO(net20));
 sg13g2_tielo tt_um_flummer_ltc_21 (.L_LO(net21));
 sg13g2_tielo tt_um_flummer_ltc_22 (.L_LO(net22));
 sg13g2_tiehi _1352__23 (.L_HI(net23));
 sg13g2_buf_2 _1588_ (.A(\ltc.timecode ),
    .X(uio_out[7]));
 sg13g2_buf_1 _1589_ (.A(uio_in[0]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1590_ (.A(uio_in[1]),
    .X(uo_out[2]));
 sg13g2_buf_1 _1591_ (.A(uio_in[2]),
    .X(uo_out[3]));
 sg13g2_buf_1 _1592_ (.A(uio_in[3]),
    .X(uo_out[4]));
 sg13g2_buf_1 _1593_ (.A(uio_in[4]),
    .X(uo_out[5]));
 sg13g2_buf_1 _1594_ (.A(uio_in[5]),
    .X(uo_out[6]));
 sg13g2_buf_1 _1595_ (.A(uio_in[6]),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout123 (.A(_0561_),
    .X(net123));
 sg13g2_buf_1 fanout124 (.A(_0561_),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(net127),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(net127),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(_0453_),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(_0452_),
    .X(net128));
 sg13g2_buf_8 fanout129 (.A(net130),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(net137),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_8 fanout132 (.A(net137),
    .X(net132));
 sg13g2_buf_1 fanout133 (.A(net137),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(net136),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(net136),
    .X(net135));
 sg13g2_buf_8 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_0196_),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(net139),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(_0194_),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(net141),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(_0194_),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(net143),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(_0193_),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0193_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(net147),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(_0179_),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(net149),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(_0179_),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(net157),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(net157),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(net153),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(net157),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net157),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net164),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(net162),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(net162),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(net162),
    .X(net160));
 sg13g2_buf_1 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(net164),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net164),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(_0178_),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net168),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net167),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(net168),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net174),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net174),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net173),
    .X(net171));
 sg13g2_buf_1 fanout172 (.A(net173),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_0155_),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(rst_n),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net181),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(net181),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(rst_n),
    .X(net181));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_flummer_ltc_9 (.L_LO(net9));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ltc.bit_counter[0] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ltc.timecode ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0130_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ltc.frm_counter[0] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold5 (.A(\ltc.bit_clk ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0143_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold7 (.A(\ltc.output_buffer[6] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0006_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ltc.output_buffer[14] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0198_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold11 (.A(\ltc.output_buffer[8] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0008_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ltc.frm_counter[21] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0464_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0102_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold16 (.A(\ltc.output_buffer[7] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold17 (.A(\ltc.output_buffer[11] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0011_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold19 (.A(\ltc.output_buffer[10] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0010_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold21 (.A(\ltc.output_buffer[4] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0004_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold23 (.A(\ltc.output_buffer[15] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold24 (.A(\ltc.output_buffer[5] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold25 (.A(\ltc.output_buffer[1] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0197_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold27 (.A(\ltc.output_buffer[13] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0013_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ltc.output_buffer[9] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ltc.output_buffer[12] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold31 (.A(\ltc.frm_counter[19] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0461_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0100_),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ltc.output_buffer[2] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold35 (.A(\ltc.bit_counter[7] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0566_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0138_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold38 (.A(\ltc.output_buffer[3] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ltc.output_buffer[54] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0055_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ltc.bit_counter[3] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0562_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0134_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold44 (.A(\ltc.output_buffer[51] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0052_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold46 (.A(\ltc.output_buffer[53] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0054_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ltc.frm_counter[2] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0456_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0083_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold51 (.A(\ltc.bit_counter[5] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0564_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0136_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ltc.output_buffer[60] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0061_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold56 (.A(\ltc.output_buffer[19] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0020_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold58 (.A(\ltc.output_buffer[62] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0063_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold60 (.A(\ltc.output_buffer[46] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0047_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ltc.output_buffer[16] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold63 (.A(\ltc.output_buffer[27] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0028_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ltc.output_buffer[36] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0037_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold67 (.A(\ltc.output_buffer[28] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0029_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ltc.output_buffer[22] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0023_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ltc.output_buffer[75] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0076_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ltc.output_buffer[45] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0046_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ltc.output_buffer[37] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0038_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ltc.output_buffer[52] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0053_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ltc.output_buffer[61] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0062_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold81 (.A(\ltc.output_buffer[38] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0039_),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ltc.output_buffer[26] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0284_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ltc.output_buffer[42] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0314_),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold87 (.A(\ltc.output_buffer[77] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0078_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold89 (.A(\ltc.output_buffer[66] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0366_),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ltc.min_d[0] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0483_),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0110_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold94 (.A(\ltc.output_buffer[64] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0364_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold96 (.A(\ltc.output_buffer[69] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0070_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ltc.output_buffer[34] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0300_),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold100 (.A(\ltc.output_buffer[18] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0202_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold102 (.A(\ltc.frm_u[0] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold103 (.A(\ltc.output_buffer[72] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0376_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ltc.output_buffer[30] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0031_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold107 (.A(\ltc.output_buffer[32] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0298_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ltc.output_buffer[29] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0030_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ltc.output_buffer[56] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0348_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold113 (.A(\ltc.output_buffer[74] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0378_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold115 (.A(\ltc.output_buffer[35] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold116 (.A(\ltc.output_buffer[49] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0329_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold118 (.A(\ltc.output_buffer[57] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold119 (.A(\ltc.output_buffer[58] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ltc.sec_d[0] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0500_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0117_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold123 (.A(\ltc.output_buffer[68] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0368_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold125 (.A(\ltc.output_buffer[44] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0045_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold127 (.A(\ltc.output_buffer[24] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0282_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold129 (.A(\ltc.frm_counter[22] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0465_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0103_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ltc.output_buffer[78] ),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0079_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold134 (.A(\ltc.output_buffer[17] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold135 (.A(\ltc.bit_counter[1] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ltc.output_buffer[70] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0071_),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ltc.output_buffer[40] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0312_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ltc.output_buffer[59] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0060_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold142 (.A(\ltc.output_buffer[21] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0275_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold144 (.A(\ltc.output_buffer[50] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold145 (.A(\ltc.output_buffer[25] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold146 (.A(\ltc.output_buffer[43] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0044_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ltc.frm_counter[23] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0467_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold150 (.A(\ltc.output_buffer[65] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold151 (.A(\ltc.output_buffer[67] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold152 (.A(\ltc.output_buffer[76] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0077_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold154 (.A(\ltc.min_d[2] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0486_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold156 (.A(_0112_),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold157 (.A(\ltc.output_buffer[48] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0328_),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ltc.bit_counter[8] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0567_),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0139_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ltc.output_buffer[41] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold163 (.A(\ltc.output_buffer[73] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ltc.frm_counter[20] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0462_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold166 (.A(\ltc.output_buffer[33] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold167 (.A(\ltc.hrs_u[1] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0475_),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold169 (.A(\ltc.sec_d[2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0503_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0119_),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold172 (.A(\ltc.min_u[1] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0492_),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold174 (.A(\ltc.min_d[1] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0484_),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold176 (.A(\ltc.sec_d[1] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0501_),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold178 (.A(\ltc.min_u[2] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0494_),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0115_),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ltc.frm_d[1] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0523_),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold183 (.A(\ltc.hrs_d[1] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold184 (.A(\ltc.sec_u[2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0517_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0122_),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold187 (.A(\ltc.frm_u[2] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0128_),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold189 (.A(\ltc.output_buffer[0] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ltc.frm_counter[5] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0459_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0086_),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold193 (.A(\ltc.frm_counter[11] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0432_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0092_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold196 (.A(\ltc.frm_counter[4] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0458_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold198 (.A(\ltc.sec_u[1] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0514_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold200 (.A(\ltc.hrs_u[0] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0399_),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ltc.frm_u[1] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold203 (.A(\ltc.hrs_d[0] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0471_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0105_),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold206 (.A(\ltc.min_u[3] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0116_),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold208 (.A(\ltc.hrs_u[2] ),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold209 (.A(\ltc.sec_u[3] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0123_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold211 (.A(\ltc.bit_counter[4] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0563_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold213 (.A(\ltc.hrs_u[3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold214 (.A(\ltc.bit_counter[9] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0568_),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ltc.bit_counter[6] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold217 (.A(\ltc.frm_counter[3] ),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0457_),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold219 (.A(\ltc.frm_u[3] ),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold220 (.A(\ltc.bit_counter[11] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0546_),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold222 (.A(\ltc.frm_counter[18] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold223 (.A(_0416_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold224 (.A(\ltc.frm_counter[1] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold225 (.A(\ltc.frm_counter[6] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold226 (.A(\ltc.min_u[0] ),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold227 (.A(\ltc.frm_counter[10] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold228 (.A(_0433_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold229 (.A(\ltc.frm_counter[15] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0436_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold231 (.A(\ltc.bit_counter[2] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold232 (.A(\ltc.frm_counter[16] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0419_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold234 (.A(\ltc.frm_counter[13] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0094_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold236 (.A(\ltc.bit_counter[10] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold237 (.A(\ltc.frm_counter[8] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold238 (.A(\ltc.sec_u[0] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold239 (.A(\ltc.frm_counter[7] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold240 (.A(\ltc.frm_counter[9] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0437_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold242 (.A(\ltc.frm_counter[12] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold243 (.A(\ltc.frm_d[0] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0521_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0124_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold246 (.A(\ltc.frm_counter[14] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold247 (.A(\ltc.frm_counter[17] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold248 (.A(\ltc.frm_counter[13] ),
    .X(net474));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_4 FILLER_4_259 ();
 sg13g2_fill_1 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_fill_2 FILLER_5_196 ();
 sg13g2_fill_1 FILLER_5_198 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_decap_8 FILLER_5_241 ();
 sg13g2_decap_4 FILLER_5_248 ();
 sg13g2_fill_2 FILLER_5_279 ();
 sg13g2_fill_1 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_fill_2 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_4 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_193 ();
 sg13g2_fill_2 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_232 ();
 sg13g2_fill_2 FILLER_6_261 ();
 sg13g2_fill_1 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_fill_1 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_decap_4 FILLER_7_250 ();
 sg13g2_fill_1 FILLER_7_254 ();
 sg13g2_fill_1 FILLER_7_286 ();
 sg13g2_fill_1 FILLER_7_300 ();
 sg13g2_decap_8 FILLER_7_310 ();
 sg13g2_decap_8 FILLER_7_317 ();
 sg13g2_decap_8 FILLER_7_324 ();
 sg13g2_decap_8 FILLER_7_331 ();
 sg13g2_decap_8 FILLER_7_338 ();
 sg13g2_decap_8 FILLER_7_345 ();
 sg13g2_decap_8 FILLER_7_352 ();
 sg13g2_decap_8 FILLER_7_359 ();
 sg13g2_decap_8 FILLER_7_366 ();
 sg13g2_decap_8 FILLER_7_373 ();
 sg13g2_decap_8 FILLER_7_380 ();
 sg13g2_decap_8 FILLER_7_387 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_189 ();
 sg13g2_fill_1 FILLER_8_191 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_222 ();
 sg13g2_decap_4 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_fill_1 FILLER_8_255 ();
 sg13g2_decap_4 FILLER_8_260 ();
 sg13g2_fill_1 FILLER_8_264 ();
 sg13g2_fill_1 FILLER_8_269 ();
 sg13g2_fill_2 FILLER_8_274 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_decap_8 FILLER_8_307 ();
 sg13g2_decap_8 FILLER_8_314 ();
 sg13g2_decap_8 FILLER_8_321 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_4 FILLER_9_175 ();
 sg13g2_fill_2 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_191 ();
 sg13g2_fill_2 FILLER_9_206 ();
 sg13g2_fill_2 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_257 ();
 sg13g2_fill_2 FILLER_9_285 ();
 sg13g2_fill_1 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_fill_2 FILLER_10_168 ();
 sg13g2_fill_1 FILLER_10_170 ();
 sg13g2_fill_2 FILLER_10_236 ();
 sg13g2_fill_1 FILLER_10_238 ();
 sg13g2_fill_2 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_285 ();
 sg13g2_decap_8 FILLER_10_302 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_fill_2 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_4 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_4 FILLER_11_175 ();
 sg13g2_fill_2 FILLER_11_179 ();
 sg13g2_fill_2 FILLER_11_220 ();
 sg13g2_fill_1 FILLER_11_246 ();
 sg13g2_decap_4 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_fill_2 FILLER_11_319 ();
 sg13g2_fill_2 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_370 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_4 FILLER_12_182 ();
 sg13g2_decap_4 FILLER_12_215 ();
 sg13g2_fill_1 FILLER_12_219 ();
 sg13g2_decap_4 FILLER_12_224 ();
 sg13g2_decap_4 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_263 ();
 sg13g2_fill_2 FILLER_12_276 ();
 sg13g2_fill_2 FILLER_12_286 ();
 sg13g2_fill_2 FILLER_12_296 ();
 sg13g2_fill_1 FILLER_12_298 ();
 sg13g2_decap_4 FILLER_12_309 ();
 sg13g2_fill_2 FILLER_12_313 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_fill_1 FILLER_13_204 ();
 sg13g2_decap_8 FILLER_13_209 ();
 sg13g2_fill_1 FILLER_13_216 ();
 sg13g2_fill_2 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_259 ();
 sg13g2_fill_2 FILLER_13_277 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_4 FILLER_14_168 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_236 ();
 sg13g2_fill_1 FILLER_14_238 ();
 sg13g2_fill_1 FILLER_14_266 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_322 ();
 sg13g2_fill_2 FILLER_14_351 ();
 sg13g2_fill_2 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_1 FILLER_15_177 ();
 sg13g2_fill_1 FILLER_15_265 ();
 sg13g2_fill_1 FILLER_15_295 ();
 sg13g2_fill_1 FILLER_15_345 ();
 sg13g2_decap_8 FILLER_15_395 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_4 FILLER_16_182 ();
 sg13g2_fill_1 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_218 ();
 sg13g2_fill_2 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_4 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_fill_2 FILLER_17_207 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_fill_2 FILLER_17_257 ();
 sg13g2_fill_1 FILLER_17_299 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_decap_4 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_fill_1 FILLER_18_196 ();
 sg13g2_fill_2 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_218 ();
 sg13g2_fill_2 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_253 ();
 sg13g2_fill_2 FILLER_18_259 ();
 sg13g2_fill_2 FILLER_18_274 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_decap_4 FILLER_18_347 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_fill_2 FILLER_19_189 ();
 sg13g2_fill_2 FILLER_19_209 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_fill_1 FILLER_19_275 ();
 sg13g2_decap_4 FILLER_19_329 ();
 sg13g2_fill_1 FILLER_19_333 ();
 sg13g2_fill_1 FILLER_19_355 ();
 sg13g2_decap_8 FILLER_19_383 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_228 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_2 FILLER_20_267 ();
 sg13g2_fill_1 FILLER_20_273 ();
 sg13g2_decap_4 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_fill_1 FILLER_20_326 ();
 sg13g2_decap_4 FILLER_20_331 ();
 sg13g2_fill_1 FILLER_20_341 ();
 sg13g2_fill_2 FILLER_20_351 ();
 sg13g2_fill_1 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_387 ();
 sg13g2_decap_8 FILLER_20_394 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_fill_2 FILLER_21_301 ();
 sg13g2_fill_1 FILLER_21_307 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_223 ();
 sg13g2_decap_4 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_307 ();
 sg13g2_fill_1 FILLER_22_309 ();
 sg13g2_decap_4 FILLER_22_345 ();
 sg13g2_fill_2 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_decap_4 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_2 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_fill_2 FILLER_23_314 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_fill_2 FILLER_23_344 ();
 sg13g2_fill_1 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_4 FILLER_24_189 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_decap_4 FILLER_24_223 ();
 sg13g2_fill_2 FILLER_24_227 ();
 sg13g2_fill_1 FILLER_24_233 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_252 ();
 sg13g2_decap_8 FILLER_24_259 ();
 sg13g2_decap_4 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_296 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_fill_1 FILLER_24_308 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_fill_2 FILLER_24_343 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_4 FILLER_25_196 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_decap_8 FILLER_25_233 ();
 sg13g2_decap_4 FILLER_25_245 ();
 sg13g2_decap_4 FILLER_25_252 ();
 sg13g2_fill_2 FILLER_25_256 ();
 sg13g2_decap_4 FILLER_25_280 ();
 sg13g2_fill_1 FILLER_25_284 ();
 sg13g2_decap_4 FILLER_25_302 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_355 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_decap_8 FILLER_25_369 ();
 sg13g2_decap_8 FILLER_25_376 ();
 sg13g2_decap_8 FILLER_25_383 ();
 sg13g2_decap_8 FILLER_25_390 ();
 sg13g2_decap_8 FILLER_25_397 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_4 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_fill_2 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_242 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_4 FILLER_27_196 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_2 FILLER_27_260 ();
 sg13g2_decap_4 FILLER_27_293 ();
 sg13g2_decap_8 FILLER_27_372 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_decap_8 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_262 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_decap_8 FILLER_29_175 ();
 sg13g2_decap_8 FILLER_29_182 ();
 sg13g2_decap_4 FILLER_29_189 ();
 sg13g2_decap_4 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_244 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_274 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_fill_2 FILLER_29_285 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_370 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_fill_2 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_fill_2 FILLER_31_189 ();
 sg13g2_fill_1 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_244 ();
 sg13g2_decap_8 FILLER_31_267 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_352 ();
 sg13g2_decap_8 FILLER_31_359 ();
 sg13g2_decap_8 FILLER_31_366 ();
 sg13g2_decap_8 FILLER_31_373 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_decap_8 FILLER_32_175 ();
 sg13g2_decap_8 FILLER_32_182 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_255 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_decap_8 FILLER_32_352 ();
 sg13g2_decap_8 FILLER_32_359 ();
 sg13g2_decap_8 FILLER_32_366 ();
 sg13g2_decap_8 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_fill_2 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_fill_1 FILLER_33_312 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_fill_1 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_decap_8 FILLER_34_147 ();
 sg13g2_decap_8 FILLER_34_154 ();
 sg13g2_decap_8 FILLER_34_161 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_decap_8 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_189 ();
 sg13g2_decap_4 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_280 ();
 sg13g2_fill_1 FILLER_34_295 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_decap_4 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_4 FILLER_35_203 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_1 FILLER_35_227 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_fill_2 FILLER_36_203 ();
 sg13g2_fill_2 FILLER_36_232 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_fill_2 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_fill_2 FILLER_37_221 ();
 sg13g2_decap_4 FILLER_37_226 ();
 sg13g2_decap_4 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_238 ();
 sg13g2_fill_2 FILLER_37_287 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_1 FILLER_37_317 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_fill_2 FILLER_37_406 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_fill_2 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_258 ();
 sg13g2_fill_2 FILLER_38_263 ();
 sg13g2_fill_1 FILLER_38_265 ();
 sg13g2_decap_4 FILLER_38_300 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_4 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_4 FILLER_39_203 ();
 sg13g2_fill_2 FILLER_39_207 ();
 sg13g2_decap_8 FILLER_39_257 ();
 sg13g2_decap_4 FILLER_39_264 ();
 sg13g2_fill_1 FILLER_39_268 ();
 sg13g2_fill_2 FILLER_39_283 ();
 sg13g2_fill_1 FILLER_39_308 ();
 sg13g2_fill_1 FILLER_39_318 ();
 sg13g2_fill_2 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_348 ();
 sg13g2_decap_8 FILLER_39_355 ();
 sg13g2_decap_8 FILLER_39_362 ();
 sg13g2_decap_8 FILLER_39_369 ();
 sg13g2_decap_8 FILLER_39_376 ();
 sg13g2_decap_8 FILLER_39_383 ();
 sg13g2_decap_8 FILLER_39_390 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_decap_4 FILLER_39_404 ();
 sg13g2_fill_1 FILLER_39_408 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_fill_2 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_198 ();
 sg13g2_fill_2 FILLER_40_207 ();
 sg13g2_fill_1 FILLER_40_209 ();
 sg13g2_fill_2 FILLER_40_245 ();
 sg13g2_fill_1 FILLER_40_247 ();
 sg13g2_fill_2 FILLER_40_275 ();
 sg13g2_decap_8 FILLER_40_341 ();
 sg13g2_decap_8 FILLER_40_348 ();
 sg13g2_decap_8 FILLER_40_355 ();
 sg13g2_decap_8 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_decap_8 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_383 ();
 sg13g2_decap_8 FILLER_40_390 ();
 sg13g2_decap_8 FILLER_40_397 ();
 sg13g2_decap_4 FILLER_40_404 ();
 sg13g2_fill_1 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_fill_2 FILLER_41_196 ();
 sg13g2_fill_1 FILLER_41_198 ();
 sg13g2_fill_1 FILLER_41_221 ();
 sg13g2_decap_4 FILLER_41_267 ();
 sg13g2_fill_1 FILLER_41_271 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_decap_4 FILLER_41_303 ();
 sg13g2_fill_2 FILLER_41_315 ();
 sg13g2_fill_2 FILLER_41_332 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_fill_2 FILLER_41_406 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_decap_8 FILLER_42_70 ();
 sg13g2_decap_8 FILLER_42_77 ();
 sg13g2_decap_8 FILLER_42_84 ();
 sg13g2_decap_8 FILLER_42_91 ();
 sg13g2_decap_8 FILLER_42_98 ();
 sg13g2_decap_8 FILLER_42_105 ();
 sg13g2_decap_8 FILLER_42_112 ();
 sg13g2_decap_8 FILLER_42_119 ();
 sg13g2_decap_8 FILLER_42_126 ();
 sg13g2_decap_8 FILLER_42_133 ();
 sg13g2_decap_8 FILLER_42_140 ();
 sg13g2_decap_8 FILLER_42_147 ();
 sg13g2_decap_8 FILLER_42_154 ();
 sg13g2_decap_8 FILLER_42_161 ();
 sg13g2_decap_8 FILLER_42_168 ();
 sg13g2_decap_8 FILLER_42_175 ();
 sg13g2_decap_8 FILLER_42_182 ();
 sg13g2_decap_8 FILLER_42_189 ();
 sg13g2_fill_2 FILLER_42_196 ();
 sg13g2_fill_2 FILLER_42_236 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_fill_1 FILLER_42_262 ();
 sg13g2_decap_8 FILLER_42_279 ();
 sg13g2_fill_2 FILLER_42_286 ();
 sg13g2_decap_4 FILLER_42_301 ();
 sg13g2_fill_1 FILLER_42_305 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_364 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_decap_8 FILLER_42_378 ();
 sg13g2_decap_8 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_decap_8 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_406 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_278 ();
 sg13g2_fill_1 FILLER_43_280 ();
 sg13g2_fill_1 FILLER_43_291 ();
 sg13g2_fill_2 FILLER_43_318 ();
 sg13g2_fill_1 FILLER_43_320 ();
 sg13g2_decap_8 FILLER_43_348 ();
 sg13g2_decap_8 FILLER_43_355 ();
 sg13g2_decap_8 FILLER_43_362 ();
 sg13g2_decap_8 FILLER_43_369 ();
 sg13g2_decap_8 FILLER_43_376 ();
 sg13g2_decap_8 FILLER_43_383 ();
 sg13g2_decap_8 FILLER_43_390 ();
 sg13g2_decap_8 FILLER_43_397 ();
 sg13g2_decap_4 FILLER_43_404 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_56 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_8 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_77 ();
 sg13g2_decap_8 FILLER_44_84 ();
 sg13g2_decap_8 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_98 ();
 sg13g2_decap_8 FILLER_44_105 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_8 FILLER_44_119 ();
 sg13g2_decap_8 FILLER_44_126 ();
 sg13g2_decap_8 FILLER_44_133 ();
 sg13g2_decap_8 FILLER_44_140 ();
 sg13g2_decap_8 FILLER_44_147 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_161 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_decap_8 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_196 ();
 sg13g2_decap_4 FILLER_44_203 ();
 sg13g2_fill_1 FILLER_44_261 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_8 FILLER_44_277 ();
 sg13g2_decap_8 FILLER_44_284 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_decap_4 FILLER_44_298 ();
 sg13g2_fill_2 FILLER_44_302 ();
 sg13g2_decap_4 FILLER_44_321 ();
 sg13g2_fill_1 FILLER_44_325 ();
 sg13g2_decap_8 FILLER_44_330 ();
 sg13g2_decap_8 FILLER_44_337 ();
 sg13g2_decap_8 FILLER_44_344 ();
 sg13g2_decap_8 FILLER_44_351 ();
 sg13g2_decap_8 FILLER_44_358 ();
 sg13g2_decap_8 FILLER_44_365 ();
 sg13g2_decap_8 FILLER_44_372 ();
 sg13g2_decap_8 FILLER_44_379 ();
 sg13g2_decap_8 FILLER_44_386 ();
 sg13g2_decap_8 FILLER_44_393 ();
 sg13g2_decap_8 FILLER_44_400 ();
 sg13g2_fill_2 FILLER_44_407 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_fill_2 FILLER_45_210 ();
 sg13g2_decap_4 FILLER_45_216 ();
 sg13g2_fill_2 FILLER_45_220 ();
 sg13g2_fill_1 FILLER_45_239 ();
 sg13g2_fill_1 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_fill_2 FILLER_45_326 ();
 sg13g2_fill_1 FILLER_45_328 ();
 sg13g2_decap_8 FILLER_45_335 ();
 sg13g2_fill_2 FILLER_45_342 ();
 sg13g2_decap_8 FILLER_45_353 ();
 sg13g2_decap_8 FILLER_45_360 ();
 sg13g2_decap_8 FILLER_45_367 ();
 sg13g2_decap_8 FILLER_45_374 ();
 sg13g2_decap_8 FILLER_45_381 ();
 sg13g2_decap_8 FILLER_45_388 ();
 sg13g2_decap_8 FILLER_45_395 ();
 sg13g2_decap_8 FILLER_45_402 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_fill_2 FILLER_46_224 ();
 sg13g2_fill_2 FILLER_46_298 ();
 sg13g2_fill_1 FILLER_46_327 ();
 sg13g2_decap_8 FILLER_46_356 ();
 sg13g2_decap_8 FILLER_46_363 ();
 sg13g2_decap_8 FILLER_46_370 ();
 sg13g2_decap_8 FILLER_46_377 ();
 sg13g2_decap_8 FILLER_46_384 ();
 sg13g2_decap_8 FILLER_46_391 ();
 sg13g2_decap_8 FILLER_46_398 ();
 sg13g2_decap_4 FILLER_46_405 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_247 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_286 ();
 sg13g2_fill_1 FILLER_47_311 ();
 sg13g2_fill_2 FILLER_47_325 ();
 sg13g2_decap_8 FILLER_47_344 ();
 sg13g2_decap_8 FILLER_47_351 ();
 sg13g2_decap_8 FILLER_47_358 ();
 sg13g2_decap_8 FILLER_47_365 ();
 sg13g2_decap_8 FILLER_47_372 ();
 sg13g2_decap_8 FILLER_47_379 ();
 sg13g2_decap_8 FILLER_47_386 ();
 sg13g2_decap_8 FILLER_47_393 ();
 sg13g2_decap_8 FILLER_47_400 ();
 sg13g2_fill_2 FILLER_47_407 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_4 FILLER_48_221 ();
 sg13g2_fill_2 FILLER_48_234 ();
 sg13g2_decap_4 FILLER_48_250 ();
 sg13g2_decap_8 FILLER_48_260 ();
 sg13g2_decap_8 FILLER_48_267 ();
 sg13g2_decap_4 FILLER_48_274 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_317 ();
 sg13g2_fill_1 FILLER_48_319 ();
 sg13g2_fill_2 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_341 ();
 sg13g2_decap_8 FILLER_48_351 ();
 sg13g2_decap_8 FILLER_48_358 ();
 sg13g2_decap_8 FILLER_48_365 ();
 sg13g2_decap_8 FILLER_48_372 ();
 sg13g2_decap_8 FILLER_48_379 ();
 sg13g2_decap_8 FILLER_48_386 ();
 sg13g2_decap_8 FILLER_48_393 ();
 sg13g2_decap_8 FILLER_48_400 ();
 sg13g2_fill_2 FILLER_48_407 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_fill_2 FILLER_49_203 ();
 sg13g2_fill_1 FILLER_49_205 ();
 sg13g2_fill_2 FILLER_49_210 ();
 sg13g2_fill_2 FILLER_49_225 ();
 sg13g2_fill_1 FILLER_49_254 ();
 sg13g2_decap_8 FILLER_49_281 ();
 sg13g2_fill_1 FILLER_49_288 ();
 sg13g2_fill_1 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_358 ();
 sg13g2_decap_8 FILLER_49_365 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_decap_8 FILLER_49_386 ();
 sg13g2_decap_8 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_4 FILLER_50_196 ();
 sg13g2_fill_1 FILLER_50_200 ();
 sg13g2_decap_4 FILLER_50_228 ();
 sg13g2_fill_2 FILLER_50_240 ();
 sg13g2_decap_4 FILLER_50_281 ();
 sg13g2_fill_1 FILLER_50_285 ();
 sg13g2_fill_1 FILLER_50_321 ();
 sg13g2_decap_8 FILLER_50_355 ();
 sg13g2_decap_8 FILLER_50_362 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_decap_8 FILLER_50_390 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_decap_8 FILLER_51_56 ();
 sg13g2_decap_8 FILLER_51_63 ();
 sg13g2_decap_8 FILLER_51_70 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_decap_8 FILLER_51_91 ();
 sg13g2_decap_8 FILLER_51_98 ();
 sg13g2_decap_8 FILLER_51_105 ();
 sg13g2_decap_8 FILLER_51_112 ();
 sg13g2_decap_8 FILLER_51_119 ();
 sg13g2_decap_8 FILLER_51_126 ();
 sg13g2_decap_8 FILLER_51_133 ();
 sg13g2_decap_8 FILLER_51_140 ();
 sg13g2_decap_8 FILLER_51_147 ();
 sg13g2_decap_8 FILLER_51_154 ();
 sg13g2_decap_8 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_168 ();
 sg13g2_decap_8 FILLER_51_175 ();
 sg13g2_decap_8 FILLER_51_182 ();
 sg13g2_decap_8 FILLER_51_189 ();
 sg13g2_decap_4 FILLER_51_196 ();
 sg13g2_fill_1 FILLER_51_200 ();
 sg13g2_decap_8 FILLER_51_214 ();
 sg13g2_fill_2 FILLER_51_230 ();
 sg13g2_fill_1 FILLER_51_250 ();
 sg13g2_fill_2 FILLER_51_260 ();
 sg13g2_decap_8 FILLER_51_307 ();
 sg13g2_fill_1 FILLER_51_314 ();
 sg13g2_fill_1 FILLER_51_337 ();
 sg13g2_decap_8 FILLER_51_351 ();
 sg13g2_decap_8 FILLER_51_358 ();
 sg13g2_decap_8 FILLER_51_365 ();
 sg13g2_decap_8 FILLER_51_372 ();
 sg13g2_decap_8 FILLER_51_379 ();
 sg13g2_decap_8 FILLER_51_386 ();
 sg13g2_decap_8 FILLER_51_393 ();
 sg13g2_decap_8 FILLER_51_400 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_8 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_fill_2 FILLER_52_196 ();
 sg13g2_fill_1 FILLER_52_198 ();
 sg13g2_fill_2 FILLER_52_220 ();
 sg13g2_fill_2 FILLER_52_254 ();
 sg13g2_fill_1 FILLER_52_256 ();
 sg13g2_fill_1 FILLER_52_267 ();
 sg13g2_decap_4 FILLER_52_285 ();
 sg13g2_fill_2 FILLER_52_289 ();
 sg13g2_fill_2 FILLER_52_295 ();
 sg13g2_fill_1 FILLER_52_297 ();
 sg13g2_fill_1 FILLER_52_302 ();
 sg13g2_decap_4 FILLER_52_322 ();
 sg13g2_fill_1 FILLER_52_326 ();
 sg13g2_decap_8 FILLER_52_349 ();
 sg13g2_decap_8 FILLER_52_356 ();
 sg13g2_decap_8 FILLER_52_363 ();
 sg13g2_decap_8 FILLER_52_370 ();
 sg13g2_decap_8 FILLER_52_377 ();
 sg13g2_decap_8 FILLER_52_384 ();
 sg13g2_decap_8 FILLER_52_391 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_4 FILLER_53_182 ();
 sg13g2_fill_1 FILLER_53_186 ();
 sg13g2_decap_4 FILLER_53_215 ();
 sg13g2_fill_1 FILLER_53_236 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_decap_4 FILLER_53_289 ();
 sg13g2_fill_2 FILLER_53_293 ();
 sg13g2_fill_2 FILLER_53_335 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_fill_2 FILLER_53_406 ();
 sg13g2_fill_1 FILLER_53_408 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_8 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_63 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_8 FILLER_54_77 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_decap_8 FILLER_54_91 ();
 sg13g2_decap_8 FILLER_54_98 ();
 sg13g2_decap_8 FILLER_54_105 ();
 sg13g2_decap_8 FILLER_54_112 ();
 sg13g2_decap_8 FILLER_54_119 ();
 sg13g2_decap_8 FILLER_54_126 ();
 sg13g2_decap_8 FILLER_54_133 ();
 sg13g2_decap_8 FILLER_54_140 ();
 sg13g2_decap_8 FILLER_54_147 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_decap_8 FILLER_54_161 ();
 sg13g2_decap_8 FILLER_54_168 ();
 sg13g2_decap_4 FILLER_54_175 ();
 sg13g2_fill_2 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_206 ();
 sg13g2_fill_2 FILLER_54_278 ();
 sg13g2_fill_1 FILLER_54_280 ();
 sg13g2_fill_2 FILLER_54_309 ();
 sg13g2_decap_8 FILLER_54_345 ();
 sg13g2_decap_8 FILLER_54_352 ();
 sg13g2_decap_8 FILLER_54_359 ();
 sg13g2_decap_8 FILLER_54_366 ();
 sg13g2_decap_8 FILLER_54_373 ();
 sg13g2_decap_8 FILLER_54_380 ();
 sg13g2_decap_8 FILLER_54_387 ();
 sg13g2_decap_8 FILLER_54_394 ();
 sg13g2_decap_8 FILLER_54_401 ();
 sg13g2_fill_1 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_fill_2 FILLER_55_253 ();
 sg13g2_fill_1 FILLER_55_268 ();
 sg13g2_decap_8 FILLER_55_317 ();
 sg13g2_fill_1 FILLER_55_324 ();
 sg13g2_decap_8 FILLER_55_330 ();
 sg13g2_decap_8 FILLER_55_337 ();
 sg13g2_decap_8 FILLER_55_344 ();
 sg13g2_decap_8 FILLER_55_351 ();
 sg13g2_decap_8 FILLER_55_358 ();
 sg13g2_decap_8 FILLER_55_365 ();
 sg13g2_decap_8 FILLER_55_372 ();
 sg13g2_decap_8 FILLER_55_379 ();
 sg13g2_decap_8 FILLER_55_386 ();
 sg13g2_decap_8 FILLER_55_393 ();
 sg13g2_decap_8 FILLER_55_400 ();
 sg13g2_fill_2 FILLER_55_407 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_8 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_70 ();
 sg13g2_decap_8 FILLER_56_77 ();
 sg13g2_decap_8 FILLER_56_84 ();
 sg13g2_decap_8 FILLER_56_91 ();
 sg13g2_decap_8 FILLER_56_98 ();
 sg13g2_decap_8 FILLER_56_105 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_8 FILLER_56_126 ();
 sg13g2_decap_8 FILLER_56_133 ();
 sg13g2_decap_8 FILLER_56_140 ();
 sg13g2_decap_8 FILLER_56_147 ();
 sg13g2_decap_8 FILLER_56_154 ();
 sg13g2_decap_8 FILLER_56_161 ();
 sg13g2_decap_8 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_175 ();
 sg13g2_decap_8 FILLER_56_182 ();
 sg13g2_decap_4 FILLER_56_189 ();
 sg13g2_fill_2 FILLER_56_193 ();
 sg13g2_decap_4 FILLER_56_233 ();
 sg13g2_fill_2 FILLER_56_260 ();
 sg13g2_fill_2 FILLER_56_275 ();
 sg13g2_fill_1 FILLER_56_277 ();
 sg13g2_decap_8 FILLER_56_350 ();
 sg13g2_decap_8 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_decap_8 FILLER_56_378 ();
 sg13g2_decap_8 FILLER_56_385 ();
 sg13g2_decap_8 FILLER_56_392 ();
 sg13g2_decap_8 FILLER_56_399 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_fill_1 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_209 ();
 sg13g2_fill_1 FILLER_57_216 ();
 sg13g2_decap_4 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_228 ();
 sg13g2_decap_8 FILLER_57_235 ();
 sg13g2_fill_1 FILLER_57_242 ();
 sg13g2_fill_1 FILLER_57_252 ();
 sg13g2_decap_4 FILLER_57_266 ();
 sg13g2_fill_1 FILLER_57_283 ();
 sg13g2_fill_2 FILLER_57_313 ();
 sg13g2_decap_8 FILLER_57_347 ();
 sg13g2_decap_8 FILLER_57_354 ();
 sg13g2_decap_8 FILLER_57_361 ();
 sg13g2_decap_8 FILLER_57_368 ();
 sg13g2_decap_8 FILLER_57_375 ();
 sg13g2_decap_8 FILLER_57_382 ();
 sg13g2_decap_8 FILLER_57_389 ();
 sg13g2_decap_8 FILLER_57_396 ();
 sg13g2_decap_4 FILLER_57_403 ();
 sg13g2_fill_2 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_decap_8 FILLER_58_140 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_fill_1 FILLER_58_196 ();
 sg13g2_fill_1 FILLER_58_266 ();
 sg13g2_decap_4 FILLER_58_308 ();
 sg13g2_fill_1 FILLER_58_312 ();
 sg13g2_fill_2 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_328 ();
 sg13g2_decap_8 FILLER_58_335 ();
 sg13g2_decap_8 FILLER_58_342 ();
 sg13g2_decap_8 FILLER_58_349 ();
 sg13g2_decap_8 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_363 ();
 sg13g2_decap_8 FILLER_58_370 ();
 sg13g2_decap_8 FILLER_58_377 ();
 sg13g2_decap_8 FILLER_58_384 ();
 sg13g2_decap_8 FILLER_58_391 ();
 sg13g2_decap_8 FILLER_58_398 ();
 sg13g2_decap_4 FILLER_58_405 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_decap_8 FILLER_59_84 ();
 sg13g2_decap_8 FILLER_59_91 ();
 sg13g2_decap_8 FILLER_59_98 ();
 sg13g2_decap_8 FILLER_59_105 ();
 sg13g2_decap_8 FILLER_59_112 ();
 sg13g2_decap_8 FILLER_59_119 ();
 sg13g2_decap_8 FILLER_59_126 ();
 sg13g2_decap_8 FILLER_59_133 ();
 sg13g2_decap_8 FILLER_59_140 ();
 sg13g2_decap_8 FILLER_59_147 ();
 sg13g2_decap_8 FILLER_59_154 ();
 sg13g2_decap_8 FILLER_59_161 ();
 sg13g2_decap_8 FILLER_59_168 ();
 sg13g2_decap_8 FILLER_59_175 ();
 sg13g2_decap_8 FILLER_59_182 ();
 sg13g2_decap_8 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_196 ();
 sg13g2_fill_2 FILLER_59_203 ();
 sg13g2_fill_2 FILLER_59_214 ();
 sg13g2_fill_2 FILLER_59_243 ();
 sg13g2_fill_2 FILLER_59_258 ();
 sg13g2_fill_1 FILLER_59_260 ();
 sg13g2_fill_2 FILLER_59_269 ();
 sg13g2_fill_1 FILLER_59_271 ();
 sg13g2_decap_8 FILLER_59_304 ();
 sg13g2_decap_8 FILLER_59_311 ();
 sg13g2_decap_8 FILLER_59_318 ();
 sg13g2_decap_4 FILLER_59_325 ();
 sg13g2_fill_1 FILLER_59_329 ();
 sg13g2_decap_8 FILLER_59_346 ();
 sg13g2_decap_8 FILLER_59_353 ();
 sg13g2_decap_8 FILLER_59_360 ();
 sg13g2_decap_8 FILLER_59_367 ();
 sg13g2_decap_8 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_decap_8 FILLER_59_388 ();
 sg13g2_decap_8 FILLER_59_395 ();
 sg13g2_decap_8 FILLER_59_402 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_decap_8 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_91 ();
 sg13g2_decap_8 FILLER_60_98 ();
 sg13g2_decap_8 FILLER_60_105 ();
 sg13g2_decap_8 FILLER_60_112 ();
 sg13g2_decap_8 FILLER_60_119 ();
 sg13g2_decap_8 FILLER_60_126 ();
 sg13g2_decap_8 FILLER_60_133 ();
 sg13g2_decap_8 FILLER_60_140 ();
 sg13g2_decap_8 FILLER_60_147 ();
 sg13g2_decap_8 FILLER_60_154 ();
 sg13g2_decap_8 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_182 ();
 sg13g2_decap_8 FILLER_60_189 ();
 sg13g2_decap_4 FILLER_60_196 ();
 sg13g2_fill_2 FILLER_60_200 ();
 sg13g2_decap_4 FILLER_60_206 ();
 sg13g2_fill_1 FILLER_60_210 ();
 sg13g2_fill_2 FILLER_60_216 ();
 sg13g2_fill_1 FILLER_60_218 ();
 sg13g2_fill_1 FILLER_60_232 ();
 sg13g2_fill_1 FILLER_60_275 ();
 sg13g2_fill_2 FILLER_60_285 ();
 sg13g2_decap_8 FILLER_60_306 ();
 sg13g2_fill_2 FILLER_60_313 ();
 sg13g2_fill_1 FILLER_60_315 ();
 sg13g2_decap_8 FILLER_60_344 ();
 sg13g2_decap_8 FILLER_60_351 ();
 sg13g2_decap_8 FILLER_60_358 ();
 sg13g2_decap_8 FILLER_60_365 ();
 sg13g2_decap_8 FILLER_60_372 ();
 sg13g2_decap_8 FILLER_60_379 ();
 sg13g2_decap_8 FILLER_60_386 ();
 sg13g2_decap_8 FILLER_60_393 ();
 sg13g2_decap_8 FILLER_60_400 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_decap_8 FILLER_61_77 ();
 sg13g2_decap_8 FILLER_61_84 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_decap_8 FILLER_61_98 ();
 sg13g2_decap_8 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_112 ();
 sg13g2_decap_8 FILLER_61_119 ();
 sg13g2_decap_8 FILLER_61_126 ();
 sg13g2_decap_8 FILLER_61_133 ();
 sg13g2_decap_8 FILLER_61_140 ();
 sg13g2_decap_8 FILLER_61_147 ();
 sg13g2_decap_8 FILLER_61_154 ();
 sg13g2_decap_8 FILLER_61_161 ();
 sg13g2_decap_8 FILLER_61_168 ();
 sg13g2_decap_8 FILLER_61_175 ();
 sg13g2_decap_8 FILLER_61_182 ();
 sg13g2_decap_8 FILLER_61_189 ();
 sg13g2_decap_8 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_203 ();
 sg13g2_decap_8 FILLER_61_210 ();
 sg13g2_fill_2 FILLER_61_285 ();
 sg13g2_fill_1 FILLER_61_287 ();
 sg13g2_fill_2 FILLER_61_302 ();
 sg13g2_fill_1 FILLER_61_304 ();
 sg13g2_fill_2 FILLER_61_333 ();
 sg13g2_decap_8 FILLER_61_344 ();
 sg13g2_decap_8 FILLER_61_351 ();
 sg13g2_decap_8 FILLER_61_358 ();
 sg13g2_decap_4 FILLER_61_369 ();
 sg13g2_fill_2 FILLER_61_373 ();
 sg13g2_decap_8 FILLER_61_384 ();
 sg13g2_decap_8 FILLER_61_391 ();
 sg13g2_decap_8 FILLER_61_398 ();
 sg13g2_decap_4 FILLER_61_405 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_decap_8 FILLER_62_91 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_4 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_204 ();
 sg13g2_decap_8 FILLER_62_211 ();
 sg13g2_decap_4 FILLER_62_218 ();
 sg13g2_fill_2 FILLER_62_222 ();
 sg13g2_decap_8 FILLER_62_269 ();
 sg13g2_fill_2 FILLER_62_276 ();
 sg13g2_fill_1 FILLER_62_278 ();
 sg13g2_decap_4 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_299 ();
 sg13g2_fill_1 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_383 ();
 sg13g2_decap_8 FILLER_62_390 ();
 sg13g2_decap_8 FILLER_62_397 ();
 sg13g2_decap_4 FILLER_62_404 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_4 FILLER_63_189 ();
 sg13g2_fill_2 FILLER_63_193 ();
 sg13g2_decap_4 FILLER_63_227 ();
 sg13g2_fill_2 FILLER_63_231 ();
 sg13g2_fill_2 FILLER_63_237 ();
 sg13g2_fill_1 FILLER_63_239 ();
 sg13g2_fill_2 FILLER_63_253 ();
 sg13g2_fill_2 FILLER_63_259 ();
 sg13g2_fill_1 FILLER_63_261 ();
 sg13g2_decap_8 FILLER_63_274 ();
 sg13g2_decap_8 FILLER_63_281 ();
 sg13g2_fill_2 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_348 ();
 sg13g2_fill_1 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_388 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_8 FILLER_64_70 ();
 sg13g2_decap_8 FILLER_64_77 ();
 sg13g2_decap_8 FILLER_64_84 ();
 sg13g2_decap_8 FILLER_64_91 ();
 sg13g2_decap_8 FILLER_64_98 ();
 sg13g2_decap_8 FILLER_64_105 ();
 sg13g2_decap_8 FILLER_64_112 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_8 FILLER_64_140 ();
 sg13g2_decap_8 FILLER_64_147 ();
 sg13g2_decap_8 FILLER_64_154 ();
 sg13g2_decap_8 FILLER_64_161 ();
 sg13g2_decap_8 FILLER_64_168 ();
 sg13g2_decap_8 FILLER_64_175 ();
 sg13g2_decap_8 FILLER_64_182 ();
 sg13g2_fill_1 FILLER_64_189 ();
 sg13g2_decap_8 FILLER_64_232 ();
 sg13g2_decap_8 FILLER_64_239 ();
 sg13g2_decap_8 FILLER_64_246 ();
 sg13g2_fill_2 FILLER_64_253 ();
 sg13g2_fill_1 FILLER_64_295 ();
 sg13g2_fill_2 FILLER_64_307 ();
 sg13g2_fill_1 FILLER_64_327 ();
 sg13g2_fill_1 FILLER_64_383 ();
 sg13g2_decap_8 FILLER_64_397 ();
 sg13g2_decap_4 FILLER_64_404 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_4 FILLER_65_182 ();
 sg13g2_decap_4 FILLER_65_214 ();
 sg13g2_decap_8 FILLER_65_227 ();
 sg13g2_fill_2 FILLER_65_234 ();
 sg13g2_decap_4 FILLER_65_240 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_332 ();
 sg13g2_decap_4 FILLER_65_346 ();
 sg13g2_fill_1 FILLER_65_364 ();
 sg13g2_fill_1 FILLER_65_370 ();
 sg13g2_decap_4 FILLER_65_403 ();
 sg13g2_fill_2 FILLER_65_407 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_decap_8 FILLER_66_84 ();
 sg13g2_decap_8 FILLER_66_91 ();
 sg13g2_decap_8 FILLER_66_98 ();
 sg13g2_decap_8 FILLER_66_105 ();
 sg13g2_decap_8 FILLER_66_112 ();
 sg13g2_decap_8 FILLER_66_119 ();
 sg13g2_decap_8 FILLER_66_126 ();
 sg13g2_decap_8 FILLER_66_133 ();
 sg13g2_decap_8 FILLER_66_140 ();
 sg13g2_decap_8 FILLER_66_147 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_161 ();
 sg13g2_decap_8 FILLER_66_168 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_decap_4 FILLER_66_182 ();
 sg13g2_decap_4 FILLER_66_323 ();
 sg13g2_fill_1 FILLER_66_327 ();
 sg13g2_fill_2 FILLER_66_345 ();
 sg13g2_fill_2 FILLER_66_375 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_fill_2 FILLER_67_182 ();
 sg13g2_fill_1 FILLER_67_184 ();
 sg13g2_fill_2 FILLER_67_219 ();
 sg13g2_fill_2 FILLER_67_249 ();
 sg13g2_fill_1 FILLER_67_251 ();
 sg13g2_fill_1 FILLER_67_257 ();
 sg13g2_decap_8 FILLER_67_289 ();
 sg13g2_decap_4 FILLER_67_301 ();
 sg13g2_fill_1 FILLER_67_305 ();
 sg13g2_decap_8 FILLER_67_310 ();
 sg13g2_decap_8 FILLER_67_317 ();
 sg13g2_fill_2 FILLER_67_332 ();
 sg13g2_fill_1 FILLER_67_334 ();
 sg13g2_fill_1 FILLER_67_363 ();
 sg13g2_decap_8 FILLER_67_401 ();
 sg13g2_fill_1 FILLER_67_408 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_8 FILLER_68_77 ();
 sg13g2_decap_8 FILLER_68_84 ();
 sg13g2_decap_8 FILLER_68_91 ();
 sg13g2_decap_8 FILLER_68_98 ();
 sg13g2_decap_8 FILLER_68_105 ();
 sg13g2_decap_8 FILLER_68_112 ();
 sg13g2_decap_8 FILLER_68_119 ();
 sg13g2_decap_8 FILLER_68_126 ();
 sg13g2_decap_8 FILLER_68_133 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_decap_8 FILLER_68_147 ();
 sg13g2_decap_8 FILLER_68_154 ();
 sg13g2_decap_8 FILLER_68_161 ();
 sg13g2_decap_8 FILLER_68_168 ();
 sg13g2_decap_8 FILLER_68_175 ();
 sg13g2_decap_8 FILLER_68_182 ();
 sg13g2_fill_1 FILLER_68_189 ();
 sg13g2_fill_2 FILLER_68_194 ();
 sg13g2_fill_2 FILLER_68_200 ();
 sg13g2_decap_8 FILLER_68_233 ();
 sg13g2_decap_8 FILLER_68_240 ();
 sg13g2_fill_1 FILLER_68_247 ();
 sg13g2_fill_2 FILLER_68_252 ();
 sg13g2_fill_1 FILLER_68_254 ();
 sg13g2_fill_1 FILLER_68_263 ();
 sg13g2_decap_4 FILLER_68_279 ();
 sg13g2_fill_2 FILLER_68_283 ();
 sg13g2_decap_8 FILLER_68_296 ();
 sg13g2_decap_8 FILLER_68_303 ();
 sg13g2_fill_2 FILLER_68_310 ();
 sg13g2_fill_1 FILLER_68_365 ();
 sg13g2_fill_2 FILLER_68_388 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_decap_8 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_98 ();
 sg13g2_decap_8 FILLER_69_105 ();
 sg13g2_decap_8 FILLER_69_112 ();
 sg13g2_decap_8 FILLER_69_119 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_decap_8 FILLER_69_133 ();
 sg13g2_decap_8 FILLER_69_140 ();
 sg13g2_decap_8 FILLER_69_147 ();
 sg13g2_decap_8 FILLER_69_154 ();
 sg13g2_decap_8 FILLER_69_161 ();
 sg13g2_decap_8 FILLER_69_168 ();
 sg13g2_decap_8 FILLER_69_175 ();
 sg13g2_decap_4 FILLER_69_182 ();
 sg13g2_fill_2 FILLER_69_186 ();
 sg13g2_decap_4 FILLER_69_202 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_211 ();
 sg13g2_fill_2 FILLER_69_231 ();
 sg13g2_fill_1 FILLER_69_233 ();
 sg13g2_fill_1 FILLER_69_280 ();
 sg13g2_decap_8 FILLER_69_284 ();
 sg13g2_decap_8 FILLER_69_291 ();
 sg13g2_fill_1 FILLER_69_298 ();
 sg13g2_fill_2 FILLER_69_356 ();
 sg13g2_fill_2 FILLER_69_376 ();
 sg13g2_fill_1 FILLER_69_378 ();
 sg13g2_fill_2 FILLER_69_407 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_fill_2 FILLER_70_175 ();
 sg13g2_decap_4 FILLER_70_240 ();
 sg13g2_fill_1 FILLER_70_266 ();
 sg13g2_decap_4 FILLER_70_296 ();
 sg13g2_fill_2 FILLER_70_328 ();
 sg13g2_decap_8 FILLER_70_402 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_decap_8 FILLER_71_70 ();
 sg13g2_decap_8 FILLER_71_77 ();
 sg13g2_decap_8 FILLER_71_84 ();
 sg13g2_decap_8 FILLER_71_91 ();
 sg13g2_decap_8 FILLER_71_98 ();
 sg13g2_decap_8 FILLER_71_105 ();
 sg13g2_decap_8 FILLER_71_112 ();
 sg13g2_decap_8 FILLER_71_119 ();
 sg13g2_decap_8 FILLER_71_126 ();
 sg13g2_decap_8 FILLER_71_133 ();
 sg13g2_decap_8 FILLER_71_140 ();
 sg13g2_decap_8 FILLER_71_147 ();
 sg13g2_decap_8 FILLER_71_154 ();
 sg13g2_decap_8 FILLER_71_161 ();
 sg13g2_decap_8 FILLER_71_168 ();
 sg13g2_decap_8 FILLER_71_175 ();
 sg13g2_fill_2 FILLER_71_186 ();
 sg13g2_decap_4 FILLER_71_237 ();
 sg13g2_decap_4 FILLER_71_246 ();
 sg13g2_fill_2 FILLER_71_269 ();
 sg13g2_fill_1 FILLER_71_281 ();
 sg13g2_decap_8 FILLER_71_310 ();
 sg13g2_fill_2 FILLER_71_317 ();
 sg13g2_fill_2 FILLER_71_328 ();
 sg13g2_fill_1 FILLER_71_347 ();
 sg13g2_fill_2 FILLER_71_393 ();
 sg13g2_decap_4 FILLER_71_404 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_fill_2 FILLER_72_175 ();
 sg13g2_fill_2 FILLER_72_236 ();
 sg13g2_fill_1 FILLER_72_238 ();
 sg13g2_fill_1 FILLER_72_276 ();
 sg13g2_fill_2 FILLER_72_282 ();
 sg13g2_decap_8 FILLER_72_299 ();
 sg13g2_fill_2 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_308 ();
 sg13g2_fill_1 FILLER_72_346 ();
 sg13g2_fill_1 FILLER_72_355 ();
 sg13g2_fill_2 FILLER_72_379 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_8 FILLER_73_91 ();
 sg13g2_decap_8 FILLER_73_98 ();
 sg13g2_decap_8 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_112 ();
 sg13g2_decap_8 FILLER_73_119 ();
 sg13g2_decap_8 FILLER_73_126 ();
 sg13g2_decap_8 FILLER_73_133 ();
 sg13g2_decap_8 FILLER_73_140 ();
 sg13g2_decap_8 FILLER_73_147 ();
 sg13g2_decap_8 FILLER_73_154 ();
 sg13g2_decap_8 FILLER_73_161 ();
 sg13g2_decap_8 FILLER_73_168 ();
 sg13g2_decap_8 FILLER_73_175 ();
 sg13g2_decap_4 FILLER_73_186 ();
 sg13g2_fill_2 FILLER_73_219 ();
 sg13g2_decap_8 FILLER_73_262 ();
 sg13g2_decap_8 FILLER_73_269 ();
 sg13g2_fill_2 FILLER_73_276 ();
 sg13g2_fill_1 FILLER_73_278 ();
 sg13g2_decap_8 FILLER_73_288 ();
 sg13g2_decap_4 FILLER_73_295 ();
 sg13g2_fill_1 FILLER_73_299 ();
 sg13g2_fill_2 FILLER_73_335 ();
 sg13g2_fill_2 FILLER_73_346 ();
 sg13g2_fill_1 FILLER_73_348 ();
 sg13g2_decap_4 FILLER_73_405 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_84 ();
 sg13g2_decap_8 FILLER_74_91 ();
 sg13g2_decap_8 FILLER_74_98 ();
 sg13g2_decap_8 FILLER_74_105 ();
 sg13g2_decap_8 FILLER_74_112 ();
 sg13g2_decap_8 FILLER_74_119 ();
 sg13g2_decap_8 FILLER_74_126 ();
 sg13g2_decap_8 FILLER_74_133 ();
 sg13g2_decap_8 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_147 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_4 FILLER_74_175 ();
 sg13g2_fill_2 FILLER_74_179 ();
 sg13g2_fill_1 FILLER_74_221 ();
 sg13g2_decap_4 FILLER_74_259 ();
 sg13g2_decap_8 FILLER_74_272 ();
 sg13g2_decap_4 FILLER_74_279 ();
 sg13g2_fill_1 FILLER_74_287 ();
 sg13g2_decap_4 FILLER_74_300 ();
 sg13g2_fill_2 FILLER_74_304 ();
 sg13g2_fill_1 FILLER_74_325 ();
 sg13g2_fill_1 FILLER_74_341 ();
 sg13g2_decap_4 FILLER_74_346 ();
 sg13g2_decap_4 FILLER_74_363 ();
 sg13g2_fill_1 FILLER_74_367 ();
 sg13g2_fill_1 FILLER_74_372 ();
 sg13g2_fill_2 FILLER_74_381 ();
 sg13g2_fill_1 FILLER_74_383 ();
 sg13g2_decap_8 FILLER_74_402 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_4 FILLER_75_182 ();
 sg13g2_decap_4 FILLER_75_190 ();
 sg13g2_fill_2 FILLER_75_194 ();
 sg13g2_fill_1 FILLER_75_208 ();
 sg13g2_fill_1 FILLER_75_315 ();
 sg13g2_fill_2 FILLER_75_326 ();
 sg13g2_decap_8 FILLER_75_352 ();
 sg13g2_fill_2 FILLER_75_359 ();
 sg13g2_fill_1 FILLER_75_361 ();
 sg13g2_decap_8 FILLER_75_387 ();
 sg13g2_decap_8 FILLER_75_394 ();
 sg13g2_decap_8 FILLER_75_401 ();
 sg13g2_fill_1 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_8 FILLER_76_84 ();
 sg13g2_decap_8 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_98 ();
 sg13g2_decap_8 FILLER_76_105 ();
 sg13g2_decap_8 FILLER_76_112 ();
 sg13g2_decap_8 FILLER_76_119 ();
 sg13g2_decap_8 FILLER_76_126 ();
 sg13g2_decap_8 FILLER_76_133 ();
 sg13g2_decap_8 FILLER_76_140 ();
 sg13g2_decap_8 FILLER_76_147 ();
 sg13g2_decap_8 FILLER_76_154 ();
 sg13g2_decap_8 FILLER_76_161 ();
 sg13g2_decap_8 FILLER_76_168 ();
 sg13g2_decap_8 FILLER_76_175 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_4 FILLER_76_189 ();
 sg13g2_fill_2 FILLER_76_243 ();
 sg13g2_fill_1 FILLER_76_245 ();
 sg13g2_fill_1 FILLER_76_274 ();
 sg13g2_fill_2 FILLER_76_284 ();
 sg13g2_fill_1 FILLER_76_286 ();
 sg13g2_fill_1 FILLER_76_309 ();
 sg13g2_fill_1 FILLER_76_337 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_390 ();
 sg13g2_decap_8 FILLER_76_397 ();
 sg13g2_decap_4 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_4 FILLER_77_182 ();
 sg13g2_fill_2 FILLER_77_186 ();
 sg13g2_fill_1 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_263 ();
 sg13g2_fill_1 FILLER_77_306 ();
 sg13g2_fill_2 FILLER_77_323 ();
 sg13g2_fill_2 FILLER_77_338 ();
 sg13g2_decap_8 FILLER_77_386 ();
 sg13g2_decap_8 FILLER_77_393 ();
 sg13g2_decap_8 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_11 ();
 sg13g2_decap_8 FILLER_78_18 ();
 sg13g2_decap_8 FILLER_78_25 ();
 sg13g2_decap_8 FILLER_78_32 ();
 sg13g2_decap_8 FILLER_78_39 ();
 sg13g2_decap_8 FILLER_78_46 ();
 sg13g2_decap_8 FILLER_78_53 ();
 sg13g2_decap_8 FILLER_78_60 ();
 sg13g2_decap_8 FILLER_78_67 ();
 sg13g2_decap_8 FILLER_78_74 ();
 sg13g2_decap_8 FILLER_78_81 ();
 sg13g2_decap_8 FILLER_78_88 ();
 sg13g2_decap_8 FILLER_78_95 ();
 sg13g2_decap_8 FILLER_78_102 ();
 sg13g2_decap_8 FILLER_78_109 ();
 sg13g2_decap_8 FILLER_78_116 ();
 sg13g2_decap_8 FILLER_78_123 ();
 sg13g2_decap_8 FILLER_78_130 ();
 sg13g2_decap_8 FILLER_78_137 ();
 sg13g2_decap_8 FILLER_78_144 ();
 sg13g2_decap_8 FILLER_78_151 ();
 sg13g2_decap_8 FILLER_78_158 ();
 sg13g2_decap_8 FILLER_78_165 ();
 sg13g2_decap_8 FILLER_78_172 ();
 sg13g2_decap_8 FILLER_78_179 ();
 sg13g2_fill_2 FILLER_78_186 ();
 sg13g2_fill_1 FILLER_78_246 ();
 sg13g2_fill_2 FILLER_78_255 ();
 sg13g2_fill_1 FILLER_78_278 ();
 sg13g2_fill_1 FILLER_78_297 ();
 sg13g2_decap_8 FILLER_78_379 ();
 sg13g2_decap_8 FILLER_78_386 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_decap_8 FILLER_78_400 ();
 sg13g2_fill_2 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_12 ();
 sg13g2_decap_8 FILLER_79_19 ();
 sg13g2_decap_8 FILLER_79_26 ();
 sg13g2_decap_8 FILLER_79_33 ();
 sg13g2_decap_8 FILLER_79_40 ();
 sg13g2_decap_8 FILLER_79_47 ();
 sg13g2_decap_8 FILLER_79_54 ();
 sg13g2_decap_8 FILLER_79_61 ();
 sg13g2_decap_8 FILLER_79_68 ();
 sg13g2_decap_8 FILLER_79_75 ();
 sg13g2_decap_8 FILLER_79_82 ();
 sg13g2_decap_8 FILLER_79_89 ();
 sg13g2_decap_8 FILLER_79_96 ();
 sg13g2_decap_8 FILLER_79_103 ();
 sg13g2_decap_8 FILLER_79_110 ();
 sg13g2_decap_8 FILLER_79_117 ();
 sg13g2_decap_8 FILLER_79_124 ();
 sg13g2_decap_8 FILLER_79_131 ();
 sg13g2_decap_8 FILLER_79_138 ();
 sg13g2_decap_8 FILLER_79_145 ();
 sg13g2_decap_8 FILLER_79_152 ();
 sg13g2_decap_8 FILLER_79_159 ();
 sg13g2_decap_8 FILLER_79_166 ();
 sg13g2_decap_8 FILLER_79_173 ();
 sg13g2_decap_8 FILLER_79_180 ();
 sg13g2_decap_8 FILLER_79_187 ();
 sg13g2_fill_1 FILLER_79_194 ();
 sg13g2_decap_8 FILLER_79_203 ();
 sg13g2_fill_1 FILLER_79_210 ();
 sg13g2_fill_1 FILLER_79_220 ();
 sg13g2_fill_1 FILLER_79_249 ();
 sg13g2_fill_1 FILLER_79_351 ();
 sg13g2_fill_2 FILLER_79_361 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_decap_8 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_399 ();
 sg13g2_fill_2 FILLER_79_406 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_8 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_123 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_decap_4 FILLER_80_132 ();
 sg13g2_decap_4 FILLER_80_140 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_fill_1 FILLER_80_215 ();
 sg13g2_decap_4 FILLER_80_232 ();
 sg13g2_decap_4 FILLER_80_245 ();
 sg13g2_decap_4 FILLER_80_253 ();
 sg13g2_fill_2 FILLER_80_257 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_fill_2 FILLER_80_270 ();
 sg13g2_decap_8 FILLER_80_276 ();
 sg13g2_decap_8 FILLER_80_283 ();
 sg13g2_decap_4 FILLER_80_290 ();
 sg13g2_decap_4 FILLER_80_307 ();
 sg13g2_fill_1 FILLER_80_311 ();
 sg13g2_fill_1 FILLER_80_324 ();
 sg13g2_fill_2 FILLER_80_337 ();
 sg13g2_fill_1 FILLER_80_339 ();
 sg13g2_decap_8 FILLER_80_383 ();
 sg13g2_decap_8 FILLER_80_390 ();
 sg13g2_decap_8 FILLER_80_397 ();
 sg13g2_decap_4 FILLER_80_404 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net226;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
endmodule
