module tt_um_vga_example (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire clknet_0_clk;
 wire \color_state[0] ;
 wire \color_state[1] ;
 wire \color_state[2] ;
 wire \dog_pos_x[0] ;
 wire \dog_pos_x[1] ;
 wire \dog_pos_x[2] ;
 wire \dog_pos_x[3] ;
 wire \dog_pos_x[4] ;
 wire \dog_pos_x[5] ;
 wire \dog_pos_x[6] ;
 wire \dog_pos_x[7] ;
 wire \dog_pos_x[8] ;
 wire \dog_pos_x[9] ;
 wire \dog_pos_y[0] ;
 wire \dog_pos_y[1] ;
 wire \dog_pos_y[2] ;
 wire \dog_pos_y[3] ;
 wire \dog_pos_y[4] ;
 wire \dog_pos_y[5] ;
 wire \dog_pos_y[6] ;
 wire \dog_pos_y[7] ;
 wire \dog_pos_y[8] ;
 wire \dog_pos_y[9] ;
 wire horz_dir;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \square_x_pos[0] ;
 wire \square_x_pos[1] ;
 wire \square_x_pos[2] ;
 wire \square_x_pos[3] ;
 wire \square_x_pos[4] ;
 wire \square_x_pos[5] ;
 wire \square_x_pos[6] ;
 wire \square_x_pos[7] ;
 wire \square_x_pos[8] ;
 wire \square_x_pos[9] ;
 wire \square_y_pos[0] ;
 wire \square_y_pos[1] ;
 wire \square_y_pos[2] ;
 wire \square_y_pos[3] ;
 wire \square_y_pos[4] ;
 wire \square_y_pos[5] ;
 wire \square_y_pos[6] ;
 wire \square_y_pos[7] ;
 wire \square_y_pos[8] ;
 wire \square_y_pos[9] ;
 wire \tick_count[0] ;
 wire \tick_count[1] ;
 wire \tick_count[2] ;
 wire \tick_count[3] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire vert_dir;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;

 sg13g2_inv_2 _1148_ (.Y(_0317_),
    .A(net452));
 sg13g2_inv_4 _1149_ (.A(net359),
    .Y(_0318_));
 sg13g2_inv_2 _1150_ (.Y(_0319_),
    .A(net449));
 sg13g2_inv_1 _1151_ (.Y(_0320_),
    .A(net354));
 sg13g2_inv_2 _1152_ (.Y(_0321_),
    .A(net352));
 sg13g2_inv_2 _1153_ (.Y(_0322_),
    .A(net356));
 sg13g2_inv_2 _1154_ (.Y(_0323_),
    .A(net440));
 sg13g2_inv_1 _1155_ (.Y(_0324_),
    .A(net441));
 sg13g2_inv_4 _1156_ (.A(net444),
    .Y(_0325_));
 sg13g2_inv_2 _1157_ (.Y(_0326_),
    .A(net446));
 sg13g2_inv_4 _1158_ (.A(net348),
    .Y(_0327_));
 sg13g2_inv_4 _1159_ (.A(net351),
    .Y(_0328_));
 sg13g2_inv_4 _1160_ (.A(net50),
    .Y(_0329_));
 sg13g2_inv_1 _1161_ (.Y(_0330_),
    .A(net378));
 sg13g2_inv_2 _1162_ (.Y(_0331_),
    .A(net380));
 sg13g2_inv_1 _1163_ (.Y(_0332_),
    .A(net382));
 sg13g2_inv_2 _1164_ (.Y(_0333_),
    .A(net372));
 sg13g2_inv_4 _1165_ (.A(net407),
    .Y(_0334_));
 sg13g2_inv_2 _1166_ (.Y(_0335_),
    .A(\dog_pos_x[6] ));
 sg13g2_inv_4 _1167_ (.A(net410),
    .Y(_0336_));
 sg13g2_inv_2 _1168_ (.Y(_0337_),
    .A(net413));
 sg13g2_inv_1 _1169_ (.Y(_0338_),
    .A(net415));
 sg13g2_inv_2 _1170_ (.Y(_0339_),
    .A(net418));
 sg13g2_inv_2 _1171_ (.Y(_0340_),
    .A(net421));
 sg13g2_inv_4 _1172_ (.A(\dog_pos_x[9] ),
    .Y(_0341_));
 sg13g2_inv_2 _1173_ (.Y(_0342_),
    .A(\dog_pos_x[7] ));
 sg13g2_inv_2 _1174_ (.Y(_0343_),
    .A(\color_state[0] ));
 sg13g2_inv_2 _1175_ (.Y(_0344_),
    .A(\color_state[1] ));
 sg13g2_inv_1 _1176_ (.Y(_0000_),
    .A(\tick_count[0] ));
 sg13g2_inv_1 _1177_ (.Y(_0345_),
    .A(net344));
 sg13g2_inv_1 _1178_ (.Y(_0346_),
    .A(net345));
 sg13g2_inv_1 _1179_ (.Y(_0347_),
    .A(net2));
 sg13g2_inv_1 _1180_ (.Y(_0348_),
    .A(\square_y_pos[9] ));
 sg13g2_inv_1 _1181_ (.Y(_0349_),
    .A(\square_x_pos[4] ));
 sg13g2_inv_2 _1182_ (.Y(_0350_),
    .A(\square_x_pos[5] ));
 sg13g2_inv_1 _1183_ (.Y(_0351_),
    .A(\square_x_pos[7] ));
 sg13g2_inv_2 _1184_ (.Y(_0352_),
    .A(\square_x_pos[8] ));
 sg13g2_inv_2 _1185_ (.Y(_0353_),
    .A(net1));
 sg13g2_inv_1 _1186_ (.Y(_0354_),
    .A(net4));
 sg13g2_inv_2 _1187_ (.Y(_0355_),
    .A(\dog_pos_y[9] ));
 sg13g2_inv_4 _1188_ (.A(net422),
    .Y(_0356_));
 sg13g2_inv_2 _1189_ (.Y(_0357_),
    .A(net450));
 sg13g2_inv_1 _1190_ (.Y(_0358_),
    .A(net7));
 sg13g2_inv_1 _1191_ (.Y(_0359_),
    .A(\square_x_pos[3] ));
 sg13g2_inv_1 _1192_ (.Y(_0360_),
    .A(\square_y_pos[0] ));
 sg13g2_and3_2 _1193_ (.X(_0361_),
    .A(net386),
    .B(net391),
    .C(net396));
 sg13g2_nand3_1 _1194_ (.B(net391),
    .C(net395),
    .A(net386),
    .Y(_0362_));
 sg13g2_a21oi_2 _1195_ (.B1(net387),
    .Y(_0363_),
    .A2(net395),
    .A1(net391));
 sg13g2_a21o_2 _1196_ (.A2(net396),
    .A1(net391),
    .B1(net386),
    .X(_0364_));
 sg13g2_a21oi_1 _1197_ (.A1(_0362_),
    .A2(_0364_),
    .Y(_0365_),
    .B1(net423));
 sg13g2_nor2b_1 _1198_ (.A(net395),
    .B_N(\hvsync_gen.hpos[0] ),
    .Y(_0366_));
 sg13g2_nor2b_1 _1199_ (.A(net424),
    .B_N(net390),
    .Y(_0367_));
 sg13g2_nand2b_1 _1200_ (.Y(_0368_),
    .B(net390),
    .A_N(net424));
 sg13g2_nor2b_1 _1201_ (.A(net390),
    .B_N(net425),
    .Y(_0369_));
 sg13g2_nand2b_1 _1202_ (.Y(_0370_),
    .B(net425),
    .A_N(net391));
 sg13g2_a221oi_1 _1203_ (.B2(_0368_),
    .C1(_0369_),
    .B1(_0366_),
    .A1(net390),
    .Y(_0371_),
    .A2(net395));
 sg13g2_nand3_1 _1204_ (.B(_0362_),
    .C(_0364_),
    .A(net423),
    .Y(_0372_));
 sg13g2_o21ai_1 _1205_ (.B1(_0372_),
    .Y(_0373_),
    .A1(_0365_),
    .A2(_0371_));
 sg13g2_xnor2_1 _1206_ (.Y(_0374_),
    .A(net334),
    .B(_0363_));
 sg13g2_a21o_1 _1207_ (.A2(_0374_),
    .A1(net420),
    .B1(_0373_),
    .X(_0375_));
 sg13g2_o21ai_1 _1208_ (.B1(net336),
    .Y(_0376_),
    .A1(net334),
    .A2(_0363_));
 sg13g2_nand3_1 _1209_ (.B(net382),
    .C(_0364_),
    .A(net379),
    .Y(_0377_));
 sg13g2_a21oi_1 _1210_ (.A1(_0376_),
    .A2(_0377_),
    .Y(_0378_),
    .B1(net418));
 sg13g2_nor2_1 _1211_ (.A(net420),
    .B(_0374_),
    .Y(_0379_));
 sg13g2_nor2_1 _1212_ (.A(_0378_),
    .B(_0379_),
    .Y(_0380_));
 sg13g2_nand3_1 _1213_ (.B(_0376_),
    .C(_0377_),
    .A(net418),
    .Y(_0381_));
 sg13g2_xnor2_1 _1214_ (.Y(_0382_),
    .A(net337),
    .B(_0376_));
 sg13g2_a22oi_1 _1215_ (.Y(_0383_),
    .B1(_0382_),
    .B2(net415),
    .A2(_0380_),
    .A1(_0375_));
 sg13g2_o21ai_1 _1216_ (.B1(net375),
    .Y(_0384_),
    .A1(net376),
    .A2(_0376_));
 sg13g2_nand3b_1 _1217_ (.B(net330),
    .C(net338),
    .Y(_0385_),
    .A_N(_0376_));
 sg13g2_and2_1 _1218_ (.A(_0384_),
    .B(_0385_),
    .X(_0386_));
 sg13g2_nor2_1 _1219_ (.A(net415),
    .B(_0382_),
    .Y(_0387_));
 sg13g2_a221oi_1 _1220_ (.B2(net401),
    .C1(_0387_),
    .B1(_0386_),
    .A1(_0381_),
    .Y(_0388_),
    .A2(_0383_));
 sg13g2_and2_1 _1221_ (.A(net375),
    .B(net373),
    .X(_0389_));
 sg13g2_nand2_2 _1222_ (.Y(_0390_),
    .A(net374),
    .B(\dog_pos_x[7] ));
 sg13g2_o21ai_1 _1223_ (.B1(_0389_),
    .Y(_0391_),
    .A1(net376),
    .A2(_0376_));
 sg13g2_xnor2_1 _1224_ (.Y(_0392_),
    .A(net329),
    .B(_0384_));
 sg13g2_nand2_1 _1225_ (.Y(_0393_),
    .A(net412),
    .B(_0392_));
 sg13g2_o21ai_1 _1226_ (.B1(_0393_),
    .Y(_0394_),
    .A1(net401),
    .A2(_0386_));
 sg13g2_or2_1 _1227_ (.X(_0395_),
    .B(_0391_),
    .A(net332));
 sg13g2_xnor2_1 _1228_ (.Y(_0396_),
    .A(net332),
    .B(_0391_));
 sg13g2_nor2_1 _1229_ (.A(net408),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_nor2_1 _1230_ (.A(net410),
    .B(_0392_),
    .Y(_0398_));
 sg13g2_nor2_1 _1231_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_o21ai_1 _1232_ (.B1(_0399_),
    .Y(_0400_),
    .A1(_0388_),
    .A2(_0394_));
 sg13g2_xnor2_1 _1233_ (.Y(_0401_),
    .A(_0341_),
    .B(_0395_));
 sg13g2_a22oi_1 _1234_ (.Y(_0402_),
    .B1(_0401_),
    .B2(net405),
    .A2(_0396_),
    .A1(net408));
 sg13g2_nor2b_2 _1235_ (.A(\dog_pos_x[9] ),
    .B_N(net405),
    .Y(_0403_));
 sg13g2_nand2_2 _1236_ (.Y(_0404_),
    .A(net405),
    .B(_0341_));
 sg13g2_nand2b_2 _1237_ (.Y(_0405_),
    .B(\dog_pos_x[9] ),
    .A_N(net405));
 sg13g2_nand2_1 _1238_ (.Y(_0406_),
    .A(_0395_),
    .B(_0405_));
 sg13g2_a22oi_1 _1239_ (.Y(_0407_),
    .B1(_0404_),
    .B2(_0406_),
    .A2(_0402_),
    .A1(_0400_));
 sg13g2_nand2_2 _1240_ (.Y(_0408_),
    .A(net353),
    .B(net352));
 sg13g2_a21oi_2 _1241_ (.B1(net355),
    .Y(_0409_),
    .A2(net357),
    .A1(net362));
 sg13g2_nor2_2 _1242_ (.A(_0408_),
    .B(_0409_),
    .Y(_0410_));
 sg13g2_xnor2_1 _1243_ (.Y(_0411_),
    .A(net349),
    .B(_0410_));
 sg13g2_and2_1 _1244_ (.A(net439),
    .B(_0411_),
    .X(_0412_));
 sg13g2_o21ai_1 _1245_ (.B1(net341),
    .Y(_0413_),
    .A1(net342),
    .A2(_0409_));
 sg13g2_nand2b_1 _1246_ (.Y(_0414_),
    .B(_0413_),
    .A_N(_0410_));
 sg13g2_nor2_1 _1247_ (.A(net442),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_nand3_1 _1248_ (.B(net358),
    .C(net355),
    .A(net362),
    .Y(_0416_));
 sg13g2_nor2b_1 _1249_ (.A(_0409_),
    .B_N(_0416_),
    .Y(_0417_));
 sg13g2_xnor2_1 _1250_ (.Y(_0418_),
    .A(net447),
    .B(_0417_));
 sg13g2_xnor2_1 _1251_ (.Y(_0419_),
    .A(net353),
    .B(_0409_));
 sg13g2_inv_1 _1252_ (.Y(_0420_),
    .A(_0419_));
 sg13g2_nand2_1 _1253_ (.Y(_0421_),
    .A(_0325_),
    .B(_0419_));
 sg13g2_xnor2_1 _1254_ (.Y(_0422_),
    .A(net444),
    .B(_0419_));
 sg13g2_nor2b_1 _1255_ (.A(_0418_),
    .B_N(_0422_),
    .Y(_0423_));
 sg13g2_nand2b_1 _1256_ (.Y(_0424_),
    .B(_0422_),
    .A_N(_0418_));
 sg13g2_xnor2_1 _1257_ (.Y(_0425_),
    .A(net361),
    .B(net358));
 sg13g2_nor2_1 _1258_ (.A(net448),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_and2_1 _1259_ (.A(\hvsync_gen.vpos[3] ),
    .B(_0425_),
    .X(_0427_));
 sg13g2_nor2_1 _1260_ (.A(net361),
    .B(net451),
    .Y(_0428_));
 sg13g2_and2_1 _1261_ (.A(\hvsync_gen.vpos[1] ),
    .B(\hvsync_gen.vpos[0] ),
    .X(_0429_));
 sg13g2_nand2b_1 _1262_ (.Y(_0430_),
    .B(net368),
    .A_N(\hvsync_gen.vpos[0] ));
 sg13g2_nor2_1 _1263_ (.A(net452),
    .B(net48),
    .Y(_0431_));
 sg13g2_a21oi_1 _1264_ (.A1(net368),
    .A2(_0431_),
    .Y(_0432_),
    .B1(net364));
 sg13g2_a21o_1 _1265_ (.A2(_0430_),
    .A1(net452),
    .B1(_0432_),
    .X(_0433_));
 sg13g2_a221oi_1 _1266_ (.B2(net452),
    .C1(_0432_),
    .B1(_0430_),
    .A1(net361),
    .Y(_0434_),
    .A2(net451));
 sg13g2_nor3_1 _1267_ (.A(_0426_),
    .B(_0428_),
    .C(_0434_),
    .Y(_0435_));
 sg13g2_o21ai_1 _1268_ (.B1(_0423_),
    .Y(_0436_),
    .A1(_0427_),
    .A2(_0435_));
 sg13g2_and3_1 _1269_ (.X(_0437_),
    .A(net447),
    .B(_0417_),
    .C(_0421_));
 sg13g2_a221oi_1 _1270_ (.B2(net444),
    .C1(_0437_),
    .B1(_0420_),
    .A1(\hvsync_gen.vpos[6] ),
    .Y(_0438_),
    .A2(_0414_));
 sg13g2_a21oi_1 _1271_ (.A1(_0436_),
    .A2(_0438_),
    .Y(_0439_),
    .B1(_0415_));
 sg13g2_nor2_1 _1272_ (.A(net439),
    .B(_0411_),
    .Y(_0440_));
 sg13g2_nand3_1 _1273_ (.B(net350),
    .C(_0410_),
    .A(net347),
    .Y(_0441_));
 sg13g2_a21o_1 _1274_ (.A2(_0410_),
    .A1(net349),
    .B1(net347),
    .X(_0442_));
 sg13g2_nand2_1 _1275_ (.Y(_0443_),
    .A(_0441_),
    .B(_0442_));
 sg13g2_nor2_1 _1276_ (.A(net435),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_nor2_1 _1277_ (.A(_0440_),
    .B(_0444_),
    .Y(_0445_));
 sg13g2_o21ai_1 _1278_ (.B1(_0445_),
    .Y(_0446_),
    .A1(_0412_),
    .A2(_0439_));
 sg13g2_nor2_2 _1279_ (.A(_0329_),
    .B(\dog_pos_y[9] ),
    .Y(_0447_));
 sg13g2_nand2_2 _1280_ (.Y(_0448_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0355_));
 sg13g2_a22oi_1 _1281_ (.Y(_0449_),
    .B1(_0447_),
    .B2(_0441_),
    .A2(_0443_),
    .A1(net435));
 sg13g2_nand2_1 _1282_ (.Y(_0450_),
    .A(_0446_),
    .B(_0449_));
 sg13g2_nor2_2 _1283_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0355_),
    .Y(_0451_));
 sg13g2_nand2_2 _1284_ (.Y(_0452_),
    .A(_0329_),
    .B(\dog_pos_y[9] ));
 sg13g2_nand2_1 _1285_ (.Y(_0453_),
    .A(_0441_),
    .B(_0452_));
 sg13g2_nand2_1 _1286_ (.Y(_0454_),
    .A(_0448_),
    .B(_0453_));
 sg13g2_a22oi_1 _1287_ (.Y(_0455_),
    .B1(_0453_),
    .B2(_0448_),
    .A2(_0449_),
    .A1(_0446_));
 sg13g2_and3_2 _1288_ (.X(_0456_),
    .A(net388),
    .B(net384),
    .C(net393));
 sg13g2_nand3_1 _1289_ (.B(net384),
    .C(net393),
    .A(net388),
    .Y(_0457_));
 sg13g2_a21oi_2 _1290_ (.B1(net384),
    .Y(_0458_),
    .A2(net393),
    .A1(net388));
 sg13g2_a21o_2 _1291_ (.A2(net393),
    .A1(net388),
    .B1(net384),
    .X(_0459_));
 sg13g2_nand2_1 _1292_ (.Y(_0460_),
    .A(_0457_),
    .B(_0459_));
 sg13g2_nand3_1 _1293_ (.B(_0457_),
    .C(_0459_),
    .A(net421),
    .Y(_0461_));
 sg13g2_xor2_1 _1294_ (.B(net392),
    .A(net387),
    .X(_0462_));
 sg13g2_nand2_1 _1295_ (.Y(_0463_),
    .A(_0356_),
    .B(_0462_));
 sg13g2_nor2_1 _1296_ (.A(_0356_),
    .B(_0462_),
    .Y(_0464_));
 sg13g2_nor2_1 _1297_ (.A(net425),
    .B(net392),
    .Y(_0465_));
 sg13g2_or2_1 _1298_ (.X(_0466_),
    .B(net390),
    .A(net424));
 sg13g2_nand2_1 _1299_ (.Y(_0467_),
    .A(net425),
    .B(net392));
 sg13g2_nor2b_1 _1300_ (.A(\hvsync_gen.hpos[0] ),
    .B_N(net395),
    .Y(_0468_));
 sg13g2_o21ai_1 _1301_ (.B1(_0467_),
    .Y(_0469_),
    .A1(_0465_),
    .A2(_0468_));
 sg13g2_a21oi_1 _1302_ (.A1(_0463_),
    .A2(_0469_),
    .Y(_0470_),
    .B1(_0464_));
 sg13g2_o21ai_1 _1303_ (.B1(net398),
    .Y(_0471_),
    .A1(_0456_),
    .A2(_0458_));
 sg13g2_xnor2_1 _1304_ (.Y(_0472_),
    .A(net380),
    .B(_0458_));
 sg13g2_nor2_1 _1305_ (.A(net419),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_a21oi_1 _1306_ (.A1(_0461_),
    .A2(_0470_),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_nor3_2 _1307_ (.A(net378),
    .B(net380),
    .C(_0459_),
    .Y(_0475_));
 sg13g2_a21oi_1 _1308_ (.A1(net335),
    .A2(_0458_),
    .Y(_0476_),
    .B1(net338));
 sg13g2_nor2_1 _1309_ (.A(_0475_),
    .B(_0476_),
    .Y(_0477_));
 sg13g2_and2_1 _1310_ (.A(net419),
    .B(_0472_),
    .X(_0478_));
 sg13g2_a221oi_1 _1311_ (.B2(net416),
    .C1(_0478_),
    .B1(_0477_),
    .A1(_0471_),
    .Y(_0479_),
    .A2(_0474_));
 sg13g2_o21ai_1 _1312_ (.B1(net400),
    .Y(_0480_),
    .A1(_0475_),
    .A2(_0476_));
 sg13g2_xnor2_1 _1313_ (.Y(_0481_),
    .A(net331),
    .B(_0475_));
 sg13g2_o21ai_1 _1314_ (.B1(_0480_),
    .Y(_0482_),
    .A1(net413),
    .A2(_0481_));
 sg13g2_nor2_1 _1315_ (.A(_0390_),
    .B(_0475_),
    .Y(_0483_));
 sg13g2_o21ai_1 _1316_ (.B1(_0342_),
    .Y(_0484_),
    .A1(net331),
    .A2(_0475_));
 sg13g2_nand2b_1 _1317_ (.Y(_0485_),
    .B(_0484_),
    .A_N(_0483_));
 sg13g2_a22oi_1 _1318_ (.Y(_0486_),
    .B1(_0485_),
    .B2(net411),
    .A2(_0481_),
    .A1(net413));
 sg13g2_o21ai_1 _1319_ (.B1(_0486_),
    .Y(_0487_),
    .A1(_0479_),
    .A2(_0482_));
 sg13g2_nand2_1 _1320_ (.Y(_0488_),
    .A(net371),
    .B(_0483_));
 sg13g2_xnor2_1 _1321_ (.Y(_0489_),
    .A(net372),
    .B(_0483_));
 sg13g2_nand2b_1 _1322_ (.Y(_0490_),
    .B(_0334_),
    .A_N(_0489_));
 sg13g2_o21ai_1 _1323_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net412),
    .A2(_0485_));
 sg13g2_nand2b_1 _1324_ (.Y(_0492_),
    .B(_0487_),
    .A_N(_0491_));
 sg13g2_a22oi_1 _1325_ (.Y(_0493_),
    .B1(_0489_),
    .B2(net408),
    .A2(_0488_),
    .A1(_0403_));
 sg13g2_nand2_1 _1326_ (.Y(_0494_),
    .A(_0405_),
    .B(_0488_));
 sg13g2_a22oi_1 _1327_ (.Y(_0495_),
    .B1(_0494_),
    .B2(_0404_),
    .A2(_0493_),
    .A1(_0492_));
 sg13g2_o21ai_1 _1328_ (.B1(_0407_),
    .Y(_0496_),
    .A1(_0455_),
    .A2(_0495_));
 sg13g2_a221oi_1 _1329_ (.B2(_0469_),
    .C1(_0464_),
    .B1(_0463_),
    .A1(net421),
    .Y(_0497_),
    .A2(_0460_));
 sg13g2_nand3_1 _1330_ (.B(_0457_),
    .C(_0459_),
    .A(net398),
    .Y(_0498_));
 sg13g2_xnor2_1 _1331_ (.Y(_0499_),
    .A(net335),
    .B(_0456_));
 sg13g2_o21ai_1 _1332_ (.B1(_0498_),
    .Y(_0500_),
    .A1(net419),
    .A2(_0499_));
 sg13g2_or2_1 _1333_ (.X(_0501_),
    .B(_0500_),
    .A(_0497_));
 sg13g2_a21oi_2 _1334_ (.B1(net338),
    .Y(_0502_),
    .A2(_0457_),
    .A1(_0331_));
 sg13g2_o21ai_1 _1335_ (.B1(net378),
    .Y(_0503_),
    .A1(net380),
    .A2(_0456_));
 sg13g2_nor3_1 _1336_ (.A(net378),
    .B(net380),
    .C(_0456_),
    .Y(_0504_));
 sg13g2_or2_1 _1337_ (.X(_0505_),
    .B(_0504_),
    .A(_0502_));
 sg13g2_a22oi_1 _1338_ (.Y(_0506_),
    .B1(_0505_),
    .B2(net416),
    .A2(_0499_),
    .A1(net419));
 sg13g2_nor2_1 _1339_ (.A(net416),
    .B(_0505_),
    .Y(_0507_));
 sg13g2_xnor2_1 _1340_ (.Y(_0508_),
    .A(net331),
    .B(_0502_));
 sg13g2_xnor2_1 _1341_ (.Y(_0509_),
    .A(net374),
    .B(_0502_));
 sg13g2_a221oi_1 _1342_ (.B2(_0337_),
    .C1(_0507_),
    .B1(_0508_),
    .A1(_0501_),
    .Y(_0510_),
    .A2(_0506_));
 sg13g2_nand2_1 _1343_ (.Y(_0511_),
    .A(net413),
    .B(_0509_));
 sg13g2_nor2_1 _1344_ (.A(_0390_),
    .B(_0503_),
    .Y(_0512_));
 sg13g2_a21oi_1 _1345_ (.A1(net374),
    .A2(_0502_),
    .Y(_0513_),
    .B1(net373));
 sg13g2_nor2_1 _1346_ (.A(_0512_),
    .B(_0513_),
    .Y(_0514_));
 sg13g2_o21ai_1 _1347_ (.B1(_0511_),
    .Y(_0515_),
    .A1(_0336_),
    .A2(_0514_));
 sg13g2_xnor2_1 _1348_ (.Y(_0516_),
    .A(net333),
    .B(_0512_));
 sg13g2_a22oi_1 _1349_ (.Y(_0517_),
    .B1(_0516_),
    .B2(_0334_),
    .A2(_0514_),
    .A1(_0336_));
 sg13g2_o21ai_1 _1350_ (.B1(_0517_),
    .Y(_0518_),
    .A1(_0510_),
    .A2(_0515_));
 sg13g2_nor2_1 _1351_ (.A(_0334_),
    .B(_0516_),
    .Y(_0519_));
 sg13g2_nor4_1 _1352_ (.A(net333),
    .B(_0341_),
    .C(_0390_),
    .D(_0503_),
    .Y(_0520_));
 sg13g2_a21oi_1 _1353_ (.A1(net372),
    .A2(_0512_),
    .Y(_0521_),
    .B1(\dog_pos_x[9] ));
 sg13g2_or2_1 _1354_ (.X(_0522_),
    .B(_0521_),
    .A(_0520_));
 sg13g2_a21oi_1 _1355_ (.A1(net405),
    .A2(_0522_),
    .Y(_0523_),
    .B1(_0519_));
 sg13g2_nor2_1 _1356_ (.A(net405),
    .B(_0521_),
    .Y(_0524_));
 sg13g2_or2_1 _1357_ (.X(_0525_),
    .B(_0524_),
    .A(_0520_));
 sg13g2_a21oi_1 _1358_ (.A1(_0518_),
    .A2(_0523_),
    .Y(_0526_),
    .B1(_0525_));
 sg13g2_and3_2 _1359_ (.X(_0527_),
    .A(net365),
    .B(net360),
    .C(net357));
 sg13g2_nand3_1 _1360_ (.B(net360),
    .C(net357),
    .A(net364),
    .Y(_0528_));
 sg13g2_a21oi_2 _1361_ (.B1(net357),
    .Y(_0529_),
    .A2(net360),
    .A1(net364));
 sg13g2_a21o_1 _1362_ (.A2(net360),
    .A1(net364),
    .B1(net357),
    .X(_0530_));
 sg13g2_o21ai_1 _1363_ (.B1(net449),
    .Y(_0531_),
    .A1(_0527_),
    .A2(_0529_));
 sg13g2_nand3_1 _1364_ (.B(_0528_),
    .C(_0530_),
    .A(_0319_),
    .Y(_0532_));
 sg13g2_xor2_1 _1365_ (.B(net360),
    .A(net364),
    .X(_0533_));
 sg13g2_and2_1 _1366_ (.A(_0357_),
    .B(_0533_),
    .X(_0534_));
 sg13g2_nand2b_1 _1367_ (.Y(_0535_),
    .B(net450),
    .A_N(_0533_));
 sg13g2_xnor2_1 _1368_ (.Y(_0536_),
    .A(_0357_),
    .B(_0533_));
 sg13g2_a21oi_1 _1369_ (.A1(_0531_),
    .A2(_0532_),
    .Y(_0537_),
    .B1(_0536_));
 sg13g2_a21oi_1 _1370_ (.A1(net452),
    .A2(_0430_),
    .Y(_0538_),
    .B1(net364));
 sg13g2_a21o_1 _1371_ (.A2(_0431_),
    .A1(net368),
    .B1(_0538_),
    .X(_0539_));
 sg13g2_nor3_1 _1372_ (.A(net364),
    .B(net360),
    .C(net357),
    .Y(_0540_));
 sg13g2_o21ai_1 _1373_ (.B1(net357),
    .Y(_0541_),
    .A1(net364),
    .A2(net360));
 sg13g2_nand2b_1 _1374_ (.Y(_0542_),
    .B(_0541_),
    .A_N(_0540_));
 sg13g2_a221oi_1 _1375_ (.B2(_0319_),
    .C1(_0537_),
    .B1(_0542_),
    .A1(_0536_),
    .Y(_0543_),
    .A2(_0539_));
 sg13g2_nor2_1 _1376_ (.A(_0319_),
    .B(_0542_),
    .Y(_0544_));
 sg13g2_and2_1 _1377_ (.A(net340),
    .B(_0540_),
    .X(_0545_));
 sg13g2_xnor2_1 _1378_ (.Y(_0546_),
    .A(net355),
    .B(_0540_));
 sg13g2_or2_1 _1379_ (.X(_0547_),
    .B(_0546_),
    .A(net446));
 sg13g2_o21ai_1 _1380_ (.B1(_0547_),
    .Y(_0548_),
    .A1(_0543_),
    .A2(_0544_));
 sg13g2_xnor2_1 _1381_ (.Y(_0549_),
    .A(net342),
    .B(_0545_));
 sg13g2_a22oi_1 _1382_ (.Y(_0550_),
    .B1(_0549_),
    .B2(net445),
    .A2(_0546_),
    .A1(net446));
 sg13g2_nor2_2 _1383_ (.A(_0408_),
    .B(_0545_),
    .Y(_0551_));
 sg13g2_o21ai_1 _1384_ (.B1(net341),
    .Y(_0552_),
    .A1(net342),
    .A2(_0545_));
 sg13g2_nand2b_1 _1385_ (.Y(_0553_),
    .B(_0552_),
    .A_N(_0551_));
 sg13g2_nand2b_1 _1386_ (.Y(_0554_),
    .B(_0325_),
    .A_N(_0549_));
 sg13g2_o21ai_1 _1387_ (.B1(_0554_),
    .Y(_0555_),
    .A1(net441),
    .A2(_0553_));
 sg13g2_a21o_1 _1388_ (.A2(_0550_),
    .A1(_0548_),
    .B1(_0555_),
    .X(_0556_));
 sg13g2_xnor2_1 _1389_ (.Y(_0557_),
    .A(net349),
    .B(_0551_));
 sg13g2_a22oi_1 _1390_ (.Y(_0558_),
    .B1(_0557_),
    .B2(net440),
    .A2(_0553_),
    .A1(net441));
 sg13g2_nand2b_1 _1391_ (.Y(_0559_),
    .B(_0323_),
    .A_N(_0557_));
 sg13g2_nand3_1 _1392_ (.B(net349),
    .C(_0551_),
    .A(net347),
    .Y(_0560_));
 sg13g2_a21o_1 _1393_ (.A2(_0551_),
    .A1(net349),
    .B1(net347),
    .X(_0561_));
 sg13g2_nand2_1 _1394_ (.Y(_0562_),
    .A(_0560_),
    .B(_0561_));
 sg13g2_o21ai_1 _1395_ (.B1(_0559_),
    .Y(_0563_),
    .A1(net434),
    .A2(_0562_));
 sg13g2_a21o_1 _1396_ (.A2(_0558_),
    .A1(_0556_),
    .B1(_0563_),
    .X(_0564_));
 sg13g2_xnor2_1 _1397_ (.Y(_0565_),
    .A(_0355_),
    .B(_0560_));
 sg13g2_a22oi_1 _1398_ (.Y(_0566_),
    .B1(_0565_),
    .B2(\hvsync_gen.vpos[9] ),
    .A2(_0562_),
    .A1(net435));
 sg13g2_a21oi_1 _1399_ (.A1(_0452_),
    .A2(_0560_),
    .Y(_0567_),
    .B1(_0447_));
 sg13g2_a21o_1 _1400_ (.A2(_0566_),
    .A1(_0564_),
    .B1(_0567_),
    .X(_0568_));
 sg13g2_a21o_1 _1401_ (.A2(_0568_),
    .A1(_0526_),
    .B1(_0407_),
    .X(_0569_));
 sg13g2_a21o_2 _1402_ (.A2(net436),
    .A1(_0327_),
    .B1(_0447_),
    .X(_0570_));
 sg13g2_nand2_1 _1403_ (.Y(_0571_),
    .A(_0452_),
    .B(_0570_));
 sg13g2_nor2_1 _1404_ (.A(_0327_),
    .B(net435),
    .Y(_0572_));
 sg13g2_nor2_1 _1405_ (.A(_0451_),
    .B(_0572_),
    .Y(_0573_));
 sg13g2_nand2_1 _1406_ (.Y(_0574_),
    .A(net340),
    .B(_0528_));
 sg13g2_a21oi_1 _1407_ (.A1(net340),
    .A2(_0528_),
    .Y(_0575_),
    .B1(_0408_));
 sg13g2_nand2_1 _1408_ (.Y(_0576_),
    .A(net350),
    .B(_0575_));
 sg13g2_nand2_1 _1409_ (.Y(_0577_),
    .A(_0573_),
    .B(_0576_));
 sg13g2_nor2_1 _1410_ (.A(_0448_),
    .B(_0572_),
    .Y(_0578_));
 sg13g2_o21ai_1 _1411_ (.B1(_0570_),
    .Y(_0579_),
    .A1(_0576_),
    .A2(_0578_));
 sg13g2_xnor2_1 _1412_ (.Y(_0580_),
    .A(net350),
    .B(_0575_));
 sg13g2_a21o_1 _1413_ (.A2(_0539_),
    .A1(_0535_),
    .B1(_0534_),
    .X(_0581_));
 sg13g2_xnor2_1 _1414_ (.Y(_0582_),
    .A(net340),
    .B(_0527_));
 sg13g2_o21ai_1 _1415_ (.B1(_0532_),
    .Y(_0583_),
    .A1(net446),
    .A2(_0582_));
 sg13g2_a21oi_1 _1416_ (.A1(_0531_),
    .A2(_0581_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_xnor2_1 _1417_ (.Y(_0585_),
    .A(net353),
    .B(_0574_));
 sg13g2_a221oi_1 _1418_ (.B2(net443),
    .C1(_0584_),
    .B1(_0585_),
    .A1(net446),
    .Y(_0586_),
    .A2(_0582_));
 sg13g2_a21oi_1 _1419_ (.A1(net353),
    .A2(_0574_),
    .Y(_0587_),
    .B1(net352));
 sg13g2_or2_1 _1420_ (.X(_0588_),
    .B(_0587_),
    .A(_0575_));
 sg13g2_nand2b_1 _1421_ (.Y(_0589_),
    .B(net403),
    .A_N(_0588_));
 sg13g2_o21ai_1 _1422_ (.B1(_0589_),
    .Y(_0590_),
    .A1(net445),
    .A2(_0585_));
 sg13g2_a22oi_1 _1423_ (.Y(_0591_),
    .B1(_0588_),
    .B2(net442),
    .A2(_0580_),
    .A1(net438));
 sg13g2_o21ai_1 _1424_ (.B1(_0591_),
    .Y(_0592_),
    .A1(_0586_),
    .A2(_0590_));
 sg13g2_o21ai_1 _1425_ (.B1(_0592_),
    .Y(_0593_),
    .A1(net439),
    .A2(_0580_));
 sg13g2_a22oi_1 _1426_ (.Y(_0594_),
    .B1(_0579_),
    .B2(_0593_),
    .A2(_0577_),
    .A1(_0571_));
 sg13g2_nand3_1 _1427_ (.B(_0569_),
    .C(_0594_),
    .A(_0496_),
    .Y(_0595_));
 sg13g2_or3_1 _1428_ (.A(net388),
    .B(net384),
    .C(net393),
    .X(_0596_));
 sg13g2_nor4_2 _1429_ (.A(net386),
    .B(net382),
    .C(net391),
    .Y(_0597_),
    .D(net396));
 sg13g2_or4_1 _1430_ (.A(net387),
    .B(net383),
    .C(net392),
    .D(net397),
    .X(_0598_));
 sg13g2_nor3_2 _1431_ (.A(net337),
    .B(net336),
    .C(_0597_),
    .Y(_0599_));
 sg13g2_nand4_1 _1432_ (.B(net379),
    .C(net375),
    .A(net377),
    .Y(_0600_),
    .D(_0598_));
 sg13g2_xnor2_1 _1433_ (.Y(_0601_),
    .A(net329),
    .B(_0600_));
 sg13g2_xnor2_1 _1434_ (.Y(_0602_),
    .A(net330),
    .B(_0599_));
 sg13g2_nor2_1 _1435_ (.A(net401),
    .B(_0602_),
    .Y(_0603_));
 sg13g2_a21oi_1 _1436_ (.A1(net411),
    .A2(_0601_),
    .Y(_0604_),
    .B1(_0603_));
 sg13g2_xnor2_1 _1437_ (.Y(_0605_),
    .A(net379),
    .B(_0597_));
 sg13g2_a21oi_1 _1438_ (.A1(net379),
    .A2(_0598_),
    .Y(_0606_),
    .B1(net377));
 sg13g2_nor2_1 _1439_ (.A(_0599_),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_o21ai_1 _1440_ (.B1(net416),
    .Y(_0608_),
    .A1(_0599_),
    .A2(_0606_));
 sg13g2_o21ai_1 _1441_ (.B1(_0608_),
    .Y(_0609_),
    .A1(net399),
    .A2(_0605_));
 sg13g2_or3_1 _1442_ (.A(net386),
    .B(net390),
    .C(net395),
    .X(_0610_));
 sg13g2_a21oi_1 _1443_ (.A1(net382),
    .A2(_0610_),
    .Y(_0611_),
    .B1(_0597_));
 sg13g2_nand2_1 _1444_ (.Y(_0612_),
    .A(net421),
    .B(_0611_));
 sg13g2_o21ai_1 _1445_ (.B1(net386),
    .Y(_0613_),
    .A1(net390),
    .A2(net395));
 sg13g2_a21o_1 _1446_ (.A2(_0613_),
    .A1(_0610_),
    .B1(net422),
    .X(_0614_));
 sg13g2_and3_1 _1447_ (.X(_0615_),
    .A(net422),
    .B(_0610_),
    .C(_0613_));
 sg13g2_mux2_1 _1448_ (.A0(net395),
    .A1(net424),
    .S(net390),
    .X(_0616_));
 sg13g2_and2_1 _1449_ (.A(net47),
    .B(net424),
    .X(_0617_));
 sg13g2_a21o_1 _1450_ (.A2(_0466_),
    .A1(_0366_),
    .B1(_0616_),
    .X(_0618_));
 sg13g2_a21oi_1 _1451_ (.A1(_0614_),
    .A2(_0618_),
    .Y(_0619_),
    .B1(_0615_));
 sg13g2_nor2_1 _1452_ (.A(net421),
    .B(_0611_),
    .Y(_0620_));
 sg13g2_and2_1 _1453_ (.A(net398),
    .B(_0611_),
    .X(_0621_));
 sg13g2_nand2b_1 _1454_ (.Y(_0622_),
    .B(net421),
    .A_N(_0611_));
 sg13g2_a221oi_1 _1455_ (.B2(_0619_),
    .C1(_0620_),
    .B1(_0612_),
    .A1(net399),
    .Y(_0623_),
    .A2(_0605_));
 sg13g2_a22oi_1 _1456_ (.Y(_0624_),
    .B1(_0607_),
    .B2(net400),
    .A2(_0602_),
    .A1(net401));
 sg13g2_o21ai_1 _1457_ (.B1(_0624_),
    .Y(_0625_),
    .A1(_0609_),
    .A2(_0623_));
 sg13g2_nand2b_1 _1458_ (.Y(_0626_),
    .B(_0336_),
    .A_N(_0601_));
 sg13g2_nand3_1 _1459_ (.B(_0389_),
    .C(_0599_),
    .A(net371),
    .Y(_0627_));
 sg13g2_o21ai_1 _1460_ (.B1(net332),
    .Y(_0628_),
    .A1(net329),
    .A2(_0600_));
 sg13g2_nand2_1 _1461_ (.Y(_0629_),
    .A(_0627_),
    .B(_0628_));
 sg13g2_o21ai_1 _1462_ (.B1(_0626_),
    .Y(_0630_),
    .A1(net408),
    .A2(_0629_));
 sg13g2_a21o_1 _1463_ (.A2(_0625_),
    .A1(_0604_),
    .B1(_0630_),
    .X(_0631_));
 sg13g2_a22oi_1 _1464_ (.Y(_0632_),
    .B1(_0629_),
    .B2(net408),
    .A2(_0627_),
    .A1(_0403_));
 sg13g2_o21ai_1 _1465_ (.B1(_0405_),
    .Y(_0633_),
    .A1(_0403_),
    .A2(_0627_));
 sg13g2_a21o_1 _1466_ (.A2(_0632_),
    .A1(_0631_),
    .B1(_0633_),
    .X(_0634_));
 sg13g2_nand4_1 _1467_ (.B(net383),
    .C(net392),
    .A(net387),
    .Y(_0635_),
    .D(net397));
 sg13g2_and2_1 _1468_ (.A(net335),
    .B(_0635_),
    .X(_0636_));
 sg13g2_xnor2_1 _1469_ (.Y(_0637_),
    .A(net335),
    .B(_0635_));
 sg13g2_xnor2_1 _1470_ (.Y(_0638_),
    .A(net334),
    .B(_0361_));
 sg13g2_xnor2_1 _1471_ (.Y(_0639_),
    .A(net383),
    .B(_0361_));
 sg13g2_nor2_1 _1472_ (.A(_0340_),
    .B(_0638_),
    .Y(_0640_));
 sg13g2_o21ai_1 _1473_ (.B1(net423),
    .Y(_0641_),
    .A1(_0361_),
    .A2(_0363_));
 sg13g2_nor3_1 _1474_ (.A(net423),
    .B(_0361_),
    .C(_0363_),
    .Y(_0642_));
 sg13g2_a21oi_1 _1475_ (.A1(_0371_),
    .A2(_0641_),
    .Y(_0643_),
    .B1(_0642_));
 sg13g2_a22oi_1 _1476_ (.Y(_0644_),
    .B1(_0638_),
    .B2(_0340_),
    .A2(_0637_),
    .A1(net399));
 sg13g2_o21ai_1 _1477_ (.B1(_0644_),
    .Y(_0645_),
    .A1(_0640_),
    .A2(_0643_));
 sg13g2_a21o_2 _1478_ (.A2(_0635_),
    .A1(net335),
    .B1(net339),
    .X(_0646_));
 sg13g2_xnor2_1 _1479_ (.Y(_0647_),
    .A(net339),
    .B(_0636_));
 sg13g2_nor2_1 _1480_ (.A(_0339_),
    .B(_0637_),
    .Y(_0648_));
 sg13g2_a21oi_1 _1481_ (.A1(net416),
    .A2(_0647_),
    .Y(_0649_),
    .B1(_0648_));
 sg13g2_nor2_1 _1482_ (.A(net417),
    .B(_0647_),
    .Y(_0650_));
 sg13g2_xnor2_1 _1483_ (.Y(_0651_),
    .A(net375),
    .B(_0646_));
 sg13g2_xnor2_1 _1484_ (.Y(_0652_),
    .A(net331),
    .B(_0646_));
 sg13g2_a221oi_1 _1485_ (.B2(net401),
    .C1(_0650_),
    .B1(_0651_),
    .A1(_0645_),
    .Y(_0653_),
    .A2(_0649_));
 sg13g2_nand2_1 _1486_ (.Y(_0654_),
    .A(net413),
    .B(_0652_));
 sg13g2_nor2_1 _1487_ (.A(_0390_),
    .B(_0646_),
    .Y(_0655_));
 sg13g2_o21ai_1 _1488_ (.B1(_0342_),
    .Y(_0656_),
    .A1(net331),
    .A2(_0646_));
 sg13g2_nor2b_1 _1489_ (.A(_0655_),
    .B_N(_0656_),
    .Y(_0657_));
 sg13g2_o21ai_1 _1490_ (.B1(_0654_),
    .Y(_0658_),
    .A1(_0336_),
    .A2(_0657_));
 sg13g2_nand2_1 _1491_ (.Y(_0659_),
    .A(net372),
    .B(_0655_));
 sg13g2_xnor2_1 _1492_ (.Y(_0660_),
    .A(net333),
    .B(_0655_));
 sg13g2_a22oi_1 _1493_ (.Y(_0661_),
    .B1(_0660_),
    .B2(_0334_),
    .A2(_0657_),
    .A1(_0336_));
 sg13g2_o21ai_1 _1494_ (.B1(_0661_),
    .Y(_0662_),
    .A1(_0653_),
    .A2(_0658_));
 sg13g2_nor2_1 _1495_ (.A(_0334_),
    .B(_0660_),
    .Y(_0663_));
 sg13g2_xnor2_1 _1496_ (.Y(_0664_),
    .A(_0341_),
    .B(_0659_));
 sg13g2_a21oi_1 _1497_ (.A1(net406),
    .A2(_0664_),
    .Y(_0665_),
    .B1(_0663_));
 sg13g2_nand2_1 _1498_ (.Y(_0666_),
    .A(_0405_),
    .B(_0659_));
 sg13g2_a22oi_1 _1499_ (.Y(_0667_),
    .B1(_0666_),
    .B2(_0404_),
    .A2(_0665_),
    .A1(_0662_));
 sg13g2_nand3_1 _1500_ (.B(net408),
    .C(_0405_),
    .A(net332),
    .Y(_0668_));
 sg13g2_nand2_2 _1501_ (.Y(_0669_),
    .A(_0404_),
    .B(_0668_));
 sg13g2_nand2_1 _1502_ (.Y(_0670_),
    .A(net375),
    .B(net401));
 sg13g2_a221oi_1 _1503_ (.B2(_0468_),
    .C1(_0367_),
    .B1(_0370_),
    .A1(net386),
    .Y(_0671_),
    .A2(_0356_));
 sg13g2_nand2b_1 _1504_ (.Y(_0672_),
    .B(net423),
    .A_N(net386));
 sg13g2_o21ai_1 _1505_ (.B1(_0672_),
    .Y(_0673_),
    .A1(net383),
    .A2(net398));
 sg13g2_a22oi_1 _1506_ (.Y(_0674_),
    .B1(net398),
    .B2(net383),
    .A2(_0339_),
    .A1(net379));
 sg13g2_o21ai_1 _1507_ (.B1(_0674_),
    .Y(_0675_),
    .A1(_0671_),
    .A2(_0673_));
 sg13g2_a22oi_1 _1508_ (.Y(_0676_),
    .B1(\hvsync_gen.hpos[4] ),
    .B2(net335),
    .A2(net416),
    .A1(net339));
 sg13g2_o21ai_1 _1509_ (.B1(_0670_),
    .Y(_0677_),
    .A1(net339),
    .A2(net416));
 sg13g2_a21o_1 _1510_ (.A2(_0676_),
    .A1(_0675_),
    .B1(_0677_),
    .X(_0678_));
 sg13g2_a22oi_1 _1511_ (.Y(_0679_),
    .B1(net329),
    .B2(net412),
    .A2(net413),
    .A1(net330));
 sg13g2_nand2_1 _1512_ (.Y(_0680_),
    .A(net371),
    .B(_0334_));
 sg13g2_and2_1 _1513_ (.A(_0405_),
    .B(_0680_),
    .X(_0681_));
 sg13g2_o21ai_1 _1514_ (.B1(_0681_),
    .Y(_0682_),
    .A1(net411),
    .A2(net329));
 sg13g2_a221oi_1 _1515_ (.B2(_0679_),
    .C1(_0682_),
    .B1(_0678_),
    .A1(net332),
    .Y(_0683_),
    .A2(net408));
 sg13g2_xnor2_1 _1516_ (.Y(_0684_),
    .A(_0356_),
    .B(_0462_));
 sg13g2_a21o_1 _1517_ (.A2(_0471_),
    .A1(_0461_),
    .B1(_0684_),
    .X(_0685_));
 sg13g2_o21ai_1 _1518_ (.B1(net384),
    .Y(_0686_),
    .A1(net388),
    .A2(net393));
 sg13g2_and3_1 _1519_ (.X(_0687_),
    .A(net421),
    .B(_0596_),
    .C(_0686_));
 sg13g2_a21oi_1 _1520_ (.A1(_0469_),
    .A2(_0684_),
    .Y(_0688_),
    .B1(_0687_));
 sg13g2_a21o_1 _1521_ (.A2(_0686_),
    .A1(_0596_),
    .B1(\hvsync_gen.hpos[3] ),
    .X(_0689_));
 sg13g2_or4_1 _1522_ (.A(net381),
    .B(net388),
    .C(net385),
    .D(net393),
    .X(_0690_));
 sg13g2_xnor2_1 _1523_ (.Y(_0691_),
    .A(net335),
    .B(_0596_));
 sg13g2_o21ai_1 _1524_ (.B1(_0689_),
    .Y(_0692_),
    .A1(net419),
    .A2(_0691_));
 sg13g2_a21o_1 _1525_ (.A2(_0688_),
    .A1(_0685_),
    .B1(_0692_),
    .X(_0693_));
 sg13g2_xnor2_1 _1526_ (.Y(_0694_),
    .A(net338),
    .B(_0690_));
 sg13g2_a22oi_1 _1527_ (.Y(_0695_),
    .B1(_0694_),
    .B2(net417),
    .A2(_0691_),
    .A1(net419));
 sg13g2_or2_1 _1528_ (.X(_0696_),
    .B(_0694_),
    .A(net416));
 sg13g2_nor3_1 _1529_ (.A(net378),
    .B(net374),
    .C(_0690_),
    .Y(_0697_));
 sg13g2_o21ai_1 _1530_ (.B1(net374),
    .Y(_0698_),
    .A1(net378),
    .A2(_0690_));
 sg13g2_nor2b_1 _1531_ (.A(_0697_),
    .B_N(_0698_),
    .Y(_0699_));
 sg13g2_o21ai_1 _1532_ (.B1(_0696_),
    .Y(_0700_),
    .A1(\hvsync_gen.hpos[6] ),
    .A2(_0699_));
 sg13g2_a21o_1 _1533_ (.A2(_0695_),
    .A1(_0693_),
    .B1(_0700_),
    .X(_0701_));
 sg13g2_nor4_2 _1534_ (.A(\dog_pos_x[5] ),
    .B(net374),
    .C(net373),
    .Y(_0702_),
    .D(_0690_));
 sg13g2_xnor2_1 _1535_ (.Y(_0703_),
    .A(net373),
    .B(_0697_));
 sg13g2_a22oi_1 _1536_ (.Y(_0704_),
    .B1(_0703_),
    .B2(net411),
    .A2(_0699_),
    .A1(net413));
 sg13g2_nand2_1 _1537_ (.Y(_0705_),
    .A(net333),
    .B(_0702_));
 sg13g2_nand3_1 _1538_ (.B(_0341_),
    .C(_0702_),
    .A(net333),
    .Y(_0706_));
 sg13g2_o21ai_1 _1539_ (.B1(_0706_),
    .Y(_0707_),
    .A1(net412),
    .A2(_0703_));
 sg13g2_xnor2_1 _1540_ (.Y(_0708_),
    .A(net372),
    .B(_0702_));
 sg13g2_nor2_1 _1541_ (.A(net409),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_or2_1 _1542_ (.X(_0710_),
    .B(_0709_),
    .A(_0707_));
 sg13g2_a21oi_1 _1543_ (.A1(_0701_),
    .A2(_0704_),
    .Y(_0711_),
    .B1(_0710_));
 sg13g2_xnor2_1 _1544_ (.Y(_0712_),
    .A(_0341_),
    .B(_0705_));
 sg13g2_a22oi_1 _1545_ (.Y(_0713_),
    .B1(_0712_),
    .B2(net405),
    .A2(_0708_),
    .A1(net408));
 sg13g2_inv_1 _1546_ (.Y(_0714_),
    .A(_0713_));
 sg13g2_nor2_1 _1547_ (.A(net405),
    .B(_0712_),
    .Y(_0715_));
 sg13g2_nor3_1 _1548_ (.A(_0669_),
    .B(_0683_),
    .C(_0715_),
    .Y(_0716_));
 sg13g2_o21ai_1 _1549_ (.B1(_0716_),
    .Y(_0717_),
    .A1(_0711_),
    .A2(_0714_));
 sg13g2_o21ai_1 _1550_ (.B1(_0717_),
    .Y(_0718_),
    .A1(_0634_),
    .A2(_0667_));
 sg13g2_nand4_1 _1551_ (.B(net359),
    .C(net354),
    .A(net363),
    .Y(_0719_),
    .D(net356));
 sg13g2_nor2_2 _1552_ (.A(net341),
    .B(_0719_),
    .Y(_0720_));
 sg13g2_nand2_2 _1553_ (.Y(_0721_),
    .A(net350),
    .B(_0720_));
 sg13g2_nand2_1 _1554_ (.Y(_0722_),
    .A(_0573_),
    .B(_0721_));
 sg13g2_nand2_1 _1555_ (.Y(_0723_),
    .A(_0571_),
    .B(_0722_));
 sg13g2_o21ai_1 _1556_ (.B1(_0418_),
    .Y(_0724_),
    .A1(_0427_),
    .A2(_0435_));
 sg13g2_xnor2_1 _1557_ (.Y(_0725_),
    .A(net342),
    .B(_0416_));
 sg13g2_nor2_1 _1558_ (.A(net444),
    .B(_0725_),
    .Y(_0726_));
 sg13g2_a21o_1 _1559_ (.A2(_0724_),
    .A1(_0424_),
    .B1(_0726_),
    .X(_0727_));
 sg13g2_xnor2_1 _1560_ (.Y(_0728_),
    .A(_0321_),
    .B(_0719_));
 sg13g2_a22oi_1 _1561_ (.Y(_0729_),
    .B1(_0728_),
    .B2(\hvsync_gen.vpos[6] ),
    .A2(_0725_),
    .A1(net445));
 sg13g2_xnor2_1 _1562_ (.Y(_0730_),
    .A(net351),
    .B(_0720_));
 sg13g2_nand2b_1 _1563_ (.Y(_0731_),
    .B(net403),
    .A_N(_0728_));
 sg13g2_o21ai_1 _1564_ (.B1(_0731_),
    .Y(_0732_),
    .A1(net439),
    .A2(_0730_));
 sg13g2_a21oi_1 _1565_ (.A1(_0727_),
    .A2(_0729_),
    .Y(_0733_),
    .B1(_0732_));
 sg13g2_xnor2_1 _1566_ (.Y(_0734_),
    .A(_0327_),
    .B(_0721_));
 sg13g2_a22oi_1 _1567_ (.Y(_0735_),
    .B1(_0734_),
    .B2(net435),
    .A2(_0730_),
    .A1(net438));
 sg13g2_inv_1 _1568_ (.Y(_0736_),
    .A(_0735_));
 sg13g2_o21ai_1 _1569_ (.B1(_0723_),
    .Y(_0737_),
    .A1(_0733_),
    .A2(_0736_));
 sg13g2_and2_1 _1570_ (.A(net365),
    .B(net368),
    .X(_0738_));
 sg13g2_nand2_2 _1571_ (.Y(_0739_),
    .A(net367),
    .B(net369));
 sg13g2_nand3_1 _1572_ (.B(net360),
    .C(net368),
    .A(net365),
    .Y(_0740_));
 sg13g2_o21ai_1 _1573_ (.B1(net340),
    .Y(_0741_),
    .A1(_0318_),
    .A2(_0740_));
 sg13g2_o21ai_1 _1574_ (.B1(_0741_),
    .Y(_0742_),
    .A1(_0416_),
    .A2(_0739_));
 sg13g2_nand2b_1 _1575_ (.Y(_0743_),
    .B(net402),
    .A_N(_0742_));
 sg13g2_xnor2_1 _1576_ (.Y(_0744_),
    .A(_0318_),
    .B(_0740_));
 sg13g2_xnor2_1 _1577_ (.Y(_0745_),
    .A(net361),
    .B(_0738_));
 sg13g2_or2_1 _1578_ (.X(_0746_),
    .B(net368),
    .A(net365));
 sg13g2_nor2_1 _1579_ (.A(net368),
    .B(\hvsync_gen.vpos[0] ),
    .Y(_0747_));
 sg13g2_nand2b_1 _1580_ (.Y(_0748_),
    .B(net452),
    .A_N(net365));
 sg13g2_xor2_1 _1581_ (.B(net368),
    .A(net365),
    .X(_0749_));
 sg13g2_a22oi_1 _1582_ (.Y(_0750_),
    .B1(_0749_),
    .B2(_0317_),
    .A2(_0748_),
    .A1(_0747_));
 sg13g2_o21ai_1 _1583_ (.B1(_0750_),
    .Y(_0751_),
    .A1(net451),
    .A2(_0745_));
 sg13g2_nor2_1 _1584_ (.A(net448),
    .B(_0744_),
    .Y(_0752_));
 sg13g2_a22oi_1 _1585_ (.Y(_0753_),
    .B1(_0745_),
    .B2(net451),
    .A2(_0744_),
    .A1(net448));
 sg13g2_a21oi_1 _1586_ (.A1(_0751_),
    .A2(_0753_),
    .Y(_0754_),
    .B1(_0752_));
 sg13g2_and2_1 _1587_ (.A(net447),
    .B(_0742_),
    .X(_0755_));
 sg13g2_nor2_1 _1588_ (.A(_0719_),
    .B(_0739_),
    .Y(_0756_));
 sg13g2_o21ai_1 _1589_ (.B1(net342),
    .Y(_0757_),
    .A1(_0416_),
    .A2(_0739_));
 sg13g2_nand2b_1 _1590_ (.Y(_0758_),
    .B(_0757_),
    .A_N(_0756_));
 sg13g2_a221oi_1 _1591_ (.B2(net444),
    .C1(_0755_),
    .B1(_0758_),
    .A1(_0743_),
    .Y(_0759_),
    .A2(_0754_));
 sg13g2_nand2_1 _1592_ (.Y(_0760_),
    .A(_0720_),
    .B(_0738_));
 sg13g2_o21ai_1 _1593_ (.B1(_0760_),
    .Y(_0761_),
    .A1(net352),
    .A2(_0756_));
 sg13g2_nand2b_1 _1594_ (.Y(_0762_),
    .B(_0325_),
    .A_N(_0758_));
 sg13g2_o21ai_1 _1595_ (.B1(_0762_),
    .Y(_0763_),
    .A1(net442),
    .A2(_0761_));
 sg13g2_xnor2_1 _1596_ (.Y(_0764_),
    .A(_0328_),
    .B(_0760_));
 sg13g2_a22oi_1 _1597_ (.Y(_0765_),
    .B1(_0764_),
    .B2(net438),
    .A2(_0761_),
    .A1(net442));
 sg13g2_o21ai_1 _1598_ (.B1(_0765_),
    .Y(_0766_),
    .A1(_0759_),
    .A2(_0763_));
 sg13g2_nor2_1 _1599_ (.A(_0451_),
    .B(_0570_),
    .Y(_0767_));
 sg13g2_nand2b_1 _1600_ (.Y(_0768_),
    .B(_0323_),
    .A_N(_0764_));
 sg13g2_nor4_1 _1601_ (.A(_0447_),
    .B(_0451_),
    .C(_0721_),
    .D(_0739_),
    .Y(_0769_));
 sg13g2_nor2_1 _1602_ (.A(_0572_),
    .B(_0769_),
    .Y(_0770_));
 sg13g2_nor3_1 _1603_ (.A(_0721_),
    .B(_0739_),
    .C(_0767_),
    .Y(_0771_));
 sg13g2_mux2_1 _1604_ (.A0(_0771_),
    .A1(_0767_),
    .S(_0770_),
    .X(_0772_));
 sg13g2_nand3_1 _1605_ (.B(_0768_),
    .C(_0772_),
    .A(_0766_),
    .Y(_0773_));
 sg13g2_nand2_1 _1606_ (.Y(_0774_),
    .A(\dog_pos_y[9] ),
    .B(_0738_));
 sg13g2_nand4_1 _1607_ (.B(net350),
    .C(_0720_),
    .A(net347),
    .Y(_0775_),
    .D(_0774_));
 sg13g2_o21ai_1 _1608_ (.B1(_0448_),
    .Y(_0776_),
    .A1(_0327_),
    .A2(_0721_));
 sg13g2_a22oi_1 _1609_ (.Y(_0777_),
    .B1(_0775_),
    .B2(_0776_),
    .A2(_0773_),
    .A1(_0571_));
 sg13g2_and3_1 _1610_ (.X(_0778_),
    .A(_0718_),
    .B(_0737_),
    .C(_0777_));
 sg13g2_o21ai_1 _1611_ (.B1(net362),
    .Y(_0779_),
    .A1(net366),
    .A2(net369));
 sg13g2_or3_1 _1612_ (.A(net366),
    .B(net362),
    .C(net369),
    .X(_0780_));
 sg13g2_and2_1 _1613_ (.A(_0779_),
    .B(_0780_),
    .X(_0781_));
 sg13g2_nor4_2 _1614_ (.A(net366),
    .B(net362),
    .C(net358),
    .Y(_0782_),
    .D(net369));
 sg13g2_a21oi_1 _1615_ (.A1(net358),
    .A2(_0780_),
    .Y(_0783_),
    .B1(_0782_));
 sg13g2_a22oi_1 _1616_ (.Y(_0784_),
    .B1(_0783_),
    .B2(net448),
    .A2(_0781_),
    .A1(net451));
 sg13g2_o21ai_1 _1617_ (.B1(_0317_),
    .Y(_0785_),
    .A1(_0738_),
    .A2(_0747_));
 sg13g2_a21oi_1 _1618_ (.A1(_0746_),
    .A2(_0785_),
    .Y(_0786_),
    .B1(_0429_));
 sg13g2_xnor2_1 _1619_ (.Y(_0787_),
    .A(net451),
    .B(_0781_));
 sg13g2_o21ai_1 _1620_ (.B1(_0784_),
    .Y(_0788_),
    .A1(_0786_),
    .A2(_0787_));
 sg13g2_nor2_1 _1621_ (.A(net448),
    .B(_0783_),
    .Y(_0789_));
 sg13g2_xnor2_1 _1622_ (.Y(_0790_),
    .A(net355),
    .B(_0782_));
 sg13g2_a21oi_1 _1623_ (.A1(net402),
    .A2(_0790_),
    .Y(_0791_),
    .B1(_0789_));
 sg13g2_nand3b_1 _1624_ (.B(net356),
    .C(net353),
    .Y(_0792_),
    .A_N(_0782_));
 sg13g2_o21ai_1 _1625_ (.B1(_0320_),
    .Y(_0793_),
    .A1(_0322_),
    .A2(_0782_));
 sg13g2_nand2_1 _1626_ (.Y(_0794_),
    .A(_0792_),
    .B(_0793_));
 sg13g2_nor2_1 _1627_ (.A(net402),
    .B(_0790_),
    .Y(_0795_));
 sg13g2_a221oi_1 _1628_ (.B2(net444),
    .C1(_0795_),
    .B1(_0794_),
    .A1(_0788_),
    .Y(_0796_),
    .A2(_0791_));
 sg13g2_nor3_1 _1629_ (.A(_0322_),
    .B(_0408_),
    .C(_0782_),
    .Y(_0797_));
 sg13g2_xnor2_1 _1630_ (.Y(_0798_),
    .A(_0321_),
    .B(_0792_));
 sg13g2_nor2_1 _1631_ (.A(net442),
    .B(_0798_),
    .Y(_0799_));
 sg13g2_nor2_1 _1632_ (.A(net444),
    .B(_0794_),
    .Y(_0800_));
 sg13g2_or2_1 _1633_ (.X(_0801_),
    .B(_0800_),
    .A(_0799_));
 sg13g2_and2_1 _1634_ (.A(net351),
    .B(_0797_),
    .X(_0802_));
 sg13g2_xnor2_1 _1635_ (.Y(_0803_),
    .A(net351),
    .B(_0797_));
 sg13g2_a22oi_1 _1636_ (.Y(_0804_),
    .B1(_0803_),
    .B2(net438),
    .A2(_0798_),
    .A1(net442));
 sg13g2_o21ai_1 _1637_ (.B1(_0804_),
    .Y(_0805_),
    .A1(_0796_),
    .A2(_0801_));
 sg13g2_nor2_1 _1638_ (.A(net438),
    .B(_0803_),
    .Y(_0806_));
 sg13g2_and2_1 _1639_ (.A(net348),
    .B(_0802_),
    .X(_0807_));
 sg13g2_xnor2_1 _1640_ (.Y(_0808_),
    .A(net348),
    .B(_0802_));
 sg13g2_nor2_1 _1641_ (.A(net435),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_nor2_1 _1642_ (.A(_0806_),
    .B(_0809_),
    .Y(_0810_));
 sg13g2_nor2_1 _1643_ (.A(_0448_),
    .B(_0807_),
    .Y(_0811_));
 sg13g2_a221oi_1 _1644_ (.B2(_0805_),
    .C1(_0811_),
    .B1(_0810_),
    .A1(net436),
    .Y(_0812_),
    .A2(_0808_));
 sg13g2_o21ai_1 _1645_ (.B1(_0448_),
    .Y(_0813_),
    .A1(_0451_),
    .A2(_0807_));
 sg13g2_nor2b_1 _1646_ (.A(_0812_),
    .B_N(_0813_),
    .Y(_0814_));
 sg13g2_xnor2_1 _1647_ (.Y(_0815_),
    .A(net361),
    .B(net451));
 sg13g2_nor3_1 _1648_ (.A(_0426_),
    .B(_0427_),
    .C(_0815_),
    .Y(_0816_));
 sg13g2_a221oi_1 _1649_ (.B2(_0815_),
    .C1(_0816_),
    .B1(_0433_),
    .A1(_0318_),
    .Y(_0817_),
    .A2(\hvsync_gen.vpos[3] ));
 sg13g2_a221oi_1 _1650_ (.B2(_0326_),
    .C1(_0817_),
    .B1(net355),
    .A1(net357),
    .Y(_0818_),
    .A2(_0319_));
 sg13g2_nand2_1 _1651_ (.Y(_0819_),
    .A(net342),
    .B(net444));
 sg13g2_o21ai_1 _1652_ (.B1(_0819_),
    .Y(_0820_),
    .A1(net355),
    .A2(_0326_));
 sg13g2_a22oi_1 _1653_ (.Y(_0821_),
    .B1(_0325_),
    .B2(net353),
    .A2(net403),
    .A1(net352));
 sg13g2_o21ai_1 _1654_ (.B1(_0821_),
    .Y(_0822_),
    .A1(_0818_),
    .A2(_0820_));
 sg13g2_a22oi_1 _1655_ (.Y(_0823_),
    .B1(_0328_),
    .B2(net438),
    .A2(net442),
    .A1(net341));
 sg13g2_a22oi_1 _1656_ (.Y(_0824_),
    .B1(_0822_),
    .B2(_0823_),
    .A2(net350),
    .A1(_0323_));
 sg13g2_a22oi_1 _1657_ (.Y(_0825_),
    .B1(_0573_),
    .B2(_0824_),
    .A2(_0570_),
    .A1(_0452_));
 sg13g2_o21ai_1 _1658_ (.B1(_0634_),
    .Y(_0826_),
    .A1(_0669_),
    .A2(_0683_));
 sg13g2_nor3_1 _1659_ (.A(_0814_),
    .B(_0825_),
    .C(_0826_),
    .Y(_0827_));
 sg13g2_nand3_1 _1660_ (.B(net355),
    .C(_0530_),
    .A(net353),
    .Y(_0828_));
 sg13g2_nor2_1 _1661_ (.A(net341),
    .B(_0828_),
    .Y(_0829_));
 sg13g2_xnor2_1 _1662_ (.Y(_0830_),
    .A(net349),
    .B(_0829_));
 sg13g2_nand2_1 _1663_ (.Y(_0831_),
    .A(net439),
    .B(_0830_));
 sg13g2_xnor2_1 _1664_ (.Y(_0832_),
    .A(net341),
    .B(_0828_));
 sg13g2_and2_1 _1665_ (.A(net441),
    .B(_0832_),
    .X(_0833_));
 sg13g2_o21ai_1 _1666_ (.B1(net342),
    .Y(_0834_),
    .A1(net340),
    .A2(_0529_));
 sg13g2_nand2_1 _1667_ (.Y(_0835_),
    .A(_0828_),
    .B(_0834_));
 sg13g2_nor2_1 _1668_ (.A(net443),
    .B(_0835_),
    .Y(_0836_));
 sg13g2_xnor2_1 _1669_ (.Y(_0837_),
    .A(net355),
    .B(_0529_));
 sg13g2_nor2_1 _1670_ (.A(net402),
    .B(_0837_),
    .Y(_0838_));
 sg13g2_a21oi_1 _1671_ (.A1(net443),
    .A2(_0835_),
    .Y(_0839_),
    .B1(_0838_));
 sg13g2_nor3_1 _1672_ (.A(_0319_),
    .B(_0527_),
    .C(_0529_),
    .Y(_0840_));
 sg13g2_a221oi_1 _1673_ (.B2(_0539_),
    .C1(_0534_),
    .B1(_0535_),
    .A1(_0531_),
    .Y(_0841_),
    .A2(_0532_));
 sg13g2_nand2_1 _1674_ (.Y(_0842_),
    .A(net402),
    .B(_0837_));
 sg13g2_o21ai_1 _1675_ (.B1(_0842_),
    .Y(_0843_),
    .A1(_0840_),
    .A2(_0841_));
 sg13g2_a21oi_1 _1676_ (.A1(_0839_),
    .A2(_0843_),
    .Y(_0844_),
    .B1(_0836_));
 sg13g2_nor2_1 _1677_ (.A(net439),
    .B(_0830_),
    .Y(_0845_));
 sg13g2_nor2_1 _1678_ (.A(net441),
    .B(_0832_),
    .Y(_0846_));
 sg13g2_nor2_1 _1679_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_o21ai_1 _1680_ (.B1(_0847_),
    .Y(_0848_),
    .A1(_0833_),
    .A2(_0844_));
 sg13g2_nand3_1 _1681_ (.B(net349),
    .C(_0829_),
    .A(net347),
    .Y(_0849_));
 sg13g2_nor2_1 _1682_ (.A(_0355_),
    .B(_0849_),
    .Y(_0850_));
 sg13g2_xor2_1 _1683_ (.B(_0849_),
    .A(\dog_pos_y[9] ),
    .X(_0851_));
 sg13g2_nand2b_1 _1684_ (.Y(_0852_),
    .B(_0329_),
    .A_N(_0851_));
 sg13g2_a21o_1 _1685_ (.A2(_0829_),
    .A1(net349),
    .B1(net347),
    .X(_0853_));
 sg13g2_nand2_1 _1686_ (.Y(_0854_),
    .A(_0849_),
    .B(_0853_));
 sg13g2_o21ai_1 _1687_ (.B1(_0852_),
    .Y(_0855_),
    .A1(net435),
    .A2(_0854_));
 sg13g2_a21o_1 _1688_ (.A2(_0848_),
    .A1(_0831_),
    .B1(_0855_),
    .X(_0856_));
 sg13g2_and3_1 _1689_ (.X(_0857_),
    .A(net435),
    .B(_0852_),
    .C(_0854_));
 sg13g2_a21oi_1 _1690_ (.A1(\hvsync_gen.vpos[9] ),
    .A2(_0851_),
    .Y(_0858_),
    .B1(_0857_));
 sg13g2_or3_1 _1691_ (.A(_0526_),
    .B(_0634_),
    .C(_0850_),
    .X(_0859_));
 sg13g2_a221oi_1 _1692_ (.B2(_0858_),
    .C1(_0859_),
    .B1(_0856_),
    .A1(_0450_),
    .Y(_0860_),
    .A2(_0454_));
 sg13g2_a21oi_2 _1693_ (.B1(net379),
    .Y(_0861_),
    .A2(_0610_),
    .A1(net382));
 sg13g2_nand3_1 _1694_ (.B(net382),
    .C(_0610_),
    .A(net379),
    .Y(_0862_));
 sg13g2_nand2b_1 _1695_ (.Y(_0863_),
    .B(_0862_),
    .A_N(_0861_));
 sg13g2_nand2_1 _1696_ (.Y(_0864_),
    .A(net399),
    .B(_0863_));
 sg13g2_o21ai_1 _1697_ (.B1(_0622_),
    .Y(_0865_),
    .A1(_0619_),
    .A2(_0621_));
 sg13g2_xnor2_1 _1698_ (.Y(_0866_),
    .A(net337),
    .B(_0861_));
 sg13g2_nor2_1 _1699_ (.A(net399),
    .B(_0863_),
    .Y(_0867_));
 sg13g2_a221oi_1 _1700_ (.B2(net415),
    .C1(_0867_),
    .B1(_0866_),
    .A1(_0864_),
    .Y(_0868_),
    .A2(_0865_));
 sg13g2_nor3_1 _1701_ (.A(net337),
    .B(net330),
    .C(_0861_),
    .Y(_0869_));
 sg13g2_o21ai_1 _1702_ (.B1(net330),
    .Y(_0870_),
    .A1(net337),
    .A2(_0861_));
 sg13g2_nand2b_1 _1703_ (.Y(_0871_),
    .B(_0870_),
    .A_N(_0869_));
 sg13g2_nand2b_1 _1704_ (.Y(_0872_),
    .B(net400),
    .A_N(_0866_));
 sg13g2_o21ai_1 _1705_ (.B1(_0872_),
    .Y(_0873_),
    .A1(net414),
    .A2(_0871_));
 sg13g2_nand2_1 _1706_ (.Y(_0874_),
    .A(net376),
    .B(_0389_));
 sg13g2_xnor2_1 _1707_ (.Y(_0875_),
    .A(net373),
    .B(_0869_));
 sg13g2_a22oi_1 _1708_ (.Y(_0876_),
    .B1(_0875_),
    .B2(net410),
    .A2(_0871_),
    .A1(net414));
 sg13g2_o21ai_1 _1709_ (.B1(_0876_),
    .Y(_0877_),
    .A1(_0868_),
    .A2(_0873_));
 sg13g2_nor3_1 _1710_ (.A(net332),
    .B(_0861_),
    .C(_0874_),
    .Y(_0878_));
 sg13g2_xnor2_1 _1711_ (.Y(_0879_),
    .A(\dog_pos_x[9] ),
    .B(_0878_));
 sg13g2_nor2_1 _1712_ (.A(net404),
    .B(_0879_),
    .Y(_0880_));
 sg13g2_nor2_1 _1713_ (.A(net410),
    .B(_0875_),
    .Y(_0881_));
 sg13g2_o21ai_1 _1714_ (.B1(net332),
    .Y(_0882_),
    .A1(_0861_),
    .A2(_0874_));
 sg13g2_nand2b_1 _1715_ (.Y(_0883_),
    .B(_0882_),
    .A_N(_0878_));
 sg13g2_nor2_1 _1716_ (.A(net407),
    .B(_0883_),
    .Y(_0884_));
 sg13g2_nor3_1 _1717_ (.A(_0880_),
    .B(_0881_),
    .C(_0884_),
    .Y(_0885_));
 sg13g2_nand2_1 _1718_ (.Y(_0886_),
    .A(net404),
    .B(_0879_));
 sg13g2_nand2_1 _1719_ (.Y(_0887_),
    .A(net407),
    .B(_0883_));
 sg13g2_o21ai_1 _1720_ (.B1(_0886_),
    .Y(_0888_),
    .A1(_0880_),
    .A2(_0887_));
 sg13g2_a21o_1 _1721_ (.A2(_0885_),
    .A1(_0877_),
    .B1(_0888_),
    .X(_0889_));
 sg13g2_nand3_1 _1722_ (.B(net334),
    .C(_0362_),
    .A(net336),
    .Y(_0890_));
 sg13g2_nand3_1 _1723_ (.B(net375),
    .C(_0890_),
    .A(net376),
    .Y(_0891_));
 sg13g2_and3_1 _1724_ (.X(_0892_),
    .A(net376),
    .B(_0389_),
    .C(_0890_));
 sg13g2_nand3_1 _1725_ (.B(_0389_),
    .C(_0890_),
    .A(net376),
    .Y(_0893_));
 sg13g2_a21o_1 _1726_ (.A2(_0893_),
    .A1(_0681_),
    .B1(_0669_),
    .X(_0894_));
 sg13g2_a221oi_1 _1727_ (.B2(_0371_),
    .C1(_0642_),
    .B1(_0641_),
    .A1(net398),
    .Y(_0895_),
    .A2(_0639_));
 sg13g2_o21ai_1 _1728_ (.B1(net379),
    .Y(_0896_),
    .A1(net383),
    .A2(_0361_));
 sg13g2_nand2_1 _1729_ (.Y(_0897_),
    .A(_0890_),
    .B(_0896_));
 sg13g2_nand3_1 _1730_ (.B(_0890_),
    .C(_0896_),
    .A(\hvsync_gen.hpos[4] ),
    .Y(_0898_));
 sg13g2_nand2_1 _1731_ (.Y(_0899_),
    .A(\hvsync_gen.hpos[3] ),
    .B(_0638_));
 sg13g2_nand3b_1 _1732_ (.B(_0898_),
    .C(_0899_),
    .Y(_0900_),
    .A_N(_0895_));
 sg13g2_xnor2_1 _1733_ (.Y(_0901_),
    .A(net337),
    .B(_0890_));
 sg13g2_a22oi_1 _1734_ (.Y(_0902_),
    .B1(_0901_),
    .B2(net400),
    .A2(_0897_),
    .A1(_0339_));
 sg13g2_nor2_1 _1735_ (.A(_0338_),
    .B(_0901_),
    .Y(_0903_));
 sg13g2_a21o_1 _1736_ (.A2(_0890_),
    .A1(net376),
    .B1(net375),
    .X(_0904_));
 sg13g2_nand2_1 _1737_ (.Y(_0905_),
    .A(_0891_),
    .B(_0904_));
 sg13g2_a221oi_1 _1738_ (.B2(net413),
    .C1(_0903_),
    .B1(_0905_),
    .A1(_0900_),
    .Y(_0906_),
    .A2(_0902_));
 sg13g2_xnor2_1 _1739_ (.Y(_0907_),
    .A(net329),
    .B(_0891_));
 sg13g2_nand3_1 _1740_ (.B(_0891_),
    .C(_0904_),
    .A(_0337_),
    .Y(_0908_));
 sg13g2_o21ai_1 _1741_ (.B1(_0908_),
    .Y(_0909_),
    .A1(net411),
    .A2(_0907_));
 sg13g2_xnor2_1 _1742_ (.Y(_0910_),
    .A(net371),
    .B(_0892_));
 sg13g2_a22oi_1 _1743_ (.Y(_0911_),
    .B1(_0910_),
    .B2(net409),
    .A2(_0907_),
    .A1(net411));
 sg13g2_o21ai_1 _1744_ (.B1(_0911_),
    .Y(_0912_),
    .A1(_0906_),
    .A2(_0909_));
 sg13g2_a21oi_1 _1745_ (.A1(net371),
    .A2(_0892_),
    .Y(_0913_),
    .B1(_0404_));
 sg13g2_a221oi_1 _1746_ (.B2(_0912_),
    .C1(_0913_),
    .B1(_0894_),
    .A1(\dog_pos_x[9] ),
    .Y(_0914_),
    .A2(_0878_));
 sg13g2_a21oi_2 _1747_ (.B1(net336),
    .Y(_0915_),
    .A2(_0613_),
    .A1(net334));
 sg13g2_a21o_1 _1748_ (.A2(_0613_),
    .A1(net334),
    .B1(net336),
    .X(_0916_));
 sg13g2_nor2_1 _1749_ (.A(net377),
    .B(_0915_),
    .Y(_0917_));
 sg13g2_a21oi_1 _1750_ (.A1(net337),
    .A2(_0916_),
    .Y(_0918_),
    .B1(net330));
 sg13g2_a21oi_1 _1751_ (.A1(net337),
    .A2(_0916_),
    .Y(_0919_),
    .B1(_0390_));
 sg13g2_xnor2_1 _1752_ (.Y(_0920_),
    .A(net373),
    .B(_0918_));
 sg13g2_nand2_1 _1753_ (.Y(_0921_),
    .A(net412),
    .B(_0920_));
 sg13g2_a21oi_1 _1754_ (.A1(_0610_),
    .A2(_0613_),
    .Y(_0922_),
    .B1(_0356_));
 sg13g2_xnor2_1 _1755_ (.Y(_0923_),
    .A(net382),
    .B(_0613_));
 sg13g2_nor2_1 _1756_ (.A(net420),
    .B(_0923_),
    .Y(_0924_));
 sg13g2_nand3_1 _1757_ (.B(_0610_),
    .C(_0613_),
    .A(_0356_),
    .Y(_0925_));
 sg13g2_and3_1 _1758_ (.X(_0926_),
    .A(net336),
    .B(net334),
    .C(_0613_));
 sg13g2_o21ai_1 _1759_ (.B1(net418),
    .Y(_0927_),
    .A1(_0915_),
    .A2(_0926_));
 sg13g2_a221oi_1 _1760_ (.B2(_0618_),
    .C1(_0922_),
    .B1(_0925_),
    .A1(net420),
    .Y(_0928_),
    .A2(_0923_));
 sg13g2_o21ai_1 _1761_ (.B1(_0927_),
    .Y(_0929_),
    .A1(_0924_),
    .A2(_0928_));
 sg13g2_xnor2_1 _1762_ (.Y(_0930_),
    .A(net377),
    .B(_0915_));
 sg13g2_nor3_1 _1763_ (.A(net418),
    .B(_0915_),
    .C(_0926_),
    .Y(_0931_));
 sg13g2_a21oi_1 _1764_ (.A1(net400),
    .A2(_0930_),
    .Y(_0932_),
    .B1(_0931_));
 sg13g2_nor2_1 _1765_ (.A(net400),
    .B(_0930_),
    .Y(_0933_));
 sg13g2_xnor2_1 _1766_ (.Y(_0934_),
    .A(net330),
    .B(_0917_));
 sg13g2_a221oi_1 _1767_ (.B2(net414),
    .C1(_0933_),
    .B1(_0934_),
    .A1(_0929_),
    .Y(_0935_),
    .A2(_0932_));
 sg13g2_nor2_1 _1768_ (.A(net414),
    .B(_0934_),
    .Y(_0936_));
 sg13g2_o21ai_1 _1769_ (.B1(_0921_),
    .Y(_0937_),
    .A1(_0935_),
    .A2(_0936_));
 sg13g2_nor4_1 _1770_ (.A(net332),
    .B(_0341_),
    .C(_0390_),
    .D(_0917_),
    .Y(_0938_));
 sg13g2_a21oi_1 _1771_ (.A1(net371),
    .A2(_0919_),
    .Y(_0939_),
    .B1(\dog_pos_x[9] ));
 sg13g2_nor3_1 _1772_ (.A(net404),
    .B(_0938_),
    .C(_0939_),
    .Y(_0940_));
 sg13g2_nor2_1 _1773_ (.A(net412),
    .B(_0920_),
    .Y(_0941_));
 sg13g2_xnor2_1 _1774_ (.Y(_0942_),
    .A(net371),
    .B(_0919_));
 sg13g2_nor2_1 _1775_ (.A(net407),
    .B(_0942_),
    .Y(_0943_));
 sg13g2_nor3_1 _1776_ (.A(_0940_),
    .B(_0941_),
    .C(_0943_),
    .Y(_0944_));
 sg13g2_o21ai_1 _1777_ (.B1(net404),
    .Y(_0945_),
    .A1(_0938_),
    .A2(_0939_));
 sg13g2_nand2_1 _1778_ (.Y(_0946_),
    .A(net409),
    .B(_0942_));
 sg13g2_o21ai_1 _1779_ (.B1(_0945_),
    .Y(_0947_),
    .A1(_0940_),
    .A2(_0946_));
 sg13g2_a21o_1 _1780_ (.A2(_0944_),
    .A1(_0937_),
    .B1(_0947_),
    .X(_0948_));
 sg13g2_a21oi_2 _1781_ (.B1(net336),
    .Y(_0949_),
    .A2(_0363_),
    .A1(net334));
 sg13g2_o21ai_1 _1782_ (.B1(net381),
    .Y(_0950_),
    .A1(net382),
    .A2(_0364_));
 sg13g2_xnor2_1 _1783_ (.Y(_0951_),
    .A(net338),
    .B(_0949_));
 sg13g2_nand2_1 _1784_ (.Y(_0952_),
    .A(net417),
    .B(_0951_));
 sg13g2_nand3_1 _1785_ (.B(_0332_),
    .C(_0363_),
    .A(net336),
    .Y(_0953_));
 sg13g2_nand2_1 _1786_ (.Y(_0954_),
    .A(_0950_),
    .B(_0953_));
 sg13g2_nor2_1 _1787_ (.A(net418),
    .B(_0954_),
    .Y(_0955_));
 sg13g2_nand2_1 _1788_ (.Y(_0956_),
    .A(net398),
    .B(_0374_));
 sg13g2_nor2_1 _1789_ (.A(net398),
    .B(_0374_),
    .Y(_0957_));
 sg13g2_a221oi_1 _1790_ (.B2(_0373_),
    .C1(_0957_),
    .B1(_0956_),
    .A1(net419),
    .Y(_0958_),
    .A2(_0954_));
 sg13g2_o21ai_1 _1791_ (.B1(_0952_),
    .Y(_0959_),
    .A1(_0955_),
    .A2(_0958_));
 sg13g2_nor2_1 _1792_ (.A(net417),
    .B(_0951_),
    .Y(_0960_));
 sg13g2_o21ai_1 _1793_ (.B1(net375),
    .Y(_0961_),
    .A1(net376),
    .A2(_0949_));
 sg13g2_nand3_1 _1794_ (.B(net330),
    .C(_0950_),
    .A(net338),
    .Y(_0962_));
 sg13g2_nand3_1 _1795_ (.B(_0961_),
    .C(_0962_),
    .A(net401),
    .Y(_0963_));
 sg13g2_nor2b_1 _1796_ (.A(_0960_),
    .B_N(_0963_),
    .Y(_0964_));
 sg13g2_o21ai_1 _1797_ (.B1(_0389_),
    .Y(_0965_),
    .A1(net377),
    .A2(_0949_));
 sg13g2_xnor2_1 _1798_ (.Y(_0966_),
    .A(net329),
    .B(_0961_));
 sg13g2_a21oi_1 _1799_ (.A1(_0961_),
    .A2(_0962_),
    .Y(_0967_),
    .B1(net401));
 sg13g2_a21o_1 _1800_ (.A2(_0966_),
    .A1(net411),
    .B1(_0967_),
    .X(_0968_));
 sg13g2_a21o_1 _1801_ (.A2(_0964_),
    .A1(_0959_),
    .B1(_0968_),
    .X(_0969_));
 sg13g2_nor2_1 _1802_ (.A(net411),
    .B(_0966_),
    .Y(_0970_));
 sg13g2_a21oi_1 _1803_ (.A1(_0681_),
    .A2(_0965_),
    .Y(_0971_),
    .B1(_0669_));
 sg13g2_nor2_1 _1804_ (.A(_0970_),
    .B(_0971_),
    .Y(_0972_));
 sg13g2_a21o_1 _1805_ (.A2(_0965_),
    .A1(_0669_),
    .B1(_0938_),
    .X(_0973_));
 sg13g2_a221oi_1 _1806_ (.B2(_0972_),
    .C1(_0973_),
    .B1(_0969_),
    .A1(_0403_),
    .Y(_0974_),
    .A2(_0680_));
 sg13g2_a22oi_1 _1807_ (.Y(_0975_),
    .B1(_0948_),
    .B2(_0974_),
    .A2(_0914_),
    .A1(_0889_));
 sg13g2_xnor2_1 _1808_ (.Y(_0976_),
    .A(net358),
    .B(_0779_));
 sg13g2_nor2_1 _1809_ (.A(net448),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_nand2_1 _1810_ (.Y(_0978_),
    .A(net448),
    .B(_0976_));
 sg13g2_xnor2_1 _1811_ (.Y(_0979_),
    .A(net448),
    .B(_0783_));
 sg13g2_mux2_1 _1812_ (.A0(_0979_),
    .A1(_0786_),
    .S(_0787_),
    .X(_0980_));
 sg13g2_a21o_1 _1813_ (.A2(_0980_),
    .A1(_0978_),
    .B1(_0977_),
    .X(_0981_));
 sg13g2_a21oi_2 _1814_ (.B1(_0322_),
    .Y(_0982_),
    .A2(_0779_),
    .A1(_0318_));
 sg13g2_nand3_1 _1815_ (.B(net340),
    .C(_0779_),
    .A(_0318_),
    .Y(_0983_));
 sg13g2_nand2b_1 _1816_ (.Y(_0984_),
    .B(_0983_),
    .A_N(_0982_));
 sg13g2_nand2_1 _1817_ (.Y(_0985_),
    .A(net447),
    .B(_0984_));
 sg13g2_xnor2_1 _1818_ (.Y(_0986_),
    .A(net354),
    .B(_0982_));
 sg13g2_nor2_1 _1819_ (.A(net447),
    .B(_0984_),
    .Y(_0987_));
 sg13g2_a221oi_1 _1820_ (.B2(_0325_),
    .C1(_0987_),
    .B1(_0986_),
    .A1(_0981_),
    .Y(_0988_),
    .A2(_0985_));
 sg13g2_o21ai_1 _1821_ (.B1(net352),
    .Y(_0989_),
    .A1(net353),
    .A2(_0982_));
 sg13g2_or3_1 _1822_ (.A(net354),
    .B(\dog_pos_y[6] ),
    .C(_0982_),
    .X(_0990_));
 sg13g2_and2_1 _1823_ (.A(_0989_),
    .B(_0990_),
    .X(_0991_));
 sg13g2_or2_1 _1824_ (.X(_0992_),
    .B(_0986_),
    .A(_0325_));
 sg13g2_o21ai_1 _1825_ (.B1(_0992_),
    .Y(_0993_),
    .A1(net403),
    .A2(_0991_));
 sg13g2_nor2_1 _1826_ (.A(_0328_),
    .B(_0989_),
    .Y(_0994_));
 sg13g2_xnor2_1 _1827_ (.Y(_0995_),
    .A(_0328_),
    .B(_0989_));
 sg13g2_nor2_1 _1828_ (.A(net438),
    .B(_0995_),
    .Y(_0996_));
 sg13g2_a21oi_1 _1829_ (.A1(_0324_),
    .A2(_0991_),
    .Y(_0997_),
    .B1(_0996_));
 sg13g2_o21ai_1 _1830_ (.B1(_0997_),
    .Y(_0998_),
    .A1(_0988_),
    .A2(_0993_));
 sg13g2_nor3_1 _1831_ (.A(_0327_),
    .B(_0328_),
    .C(_0989_),
    .Y(_0999_));
 sg13g2_xnor2_1 _1832_ (.Y(_1000_),
    .A(net348),
    .B(_0994_));
 sg13g2_a22oi_1 _1833_ (.Y(_1001_),
    .B1(_1000_),
    .B2(net436),
    .A2(_0995_),
    .A1(net438));
 sg13g2_a21oi_1 _1834_ (.A1(_0448_),
    .A2(_0999_),
    .Y(_1002_),
    .B1(_0451_));
 sg13g2_o21ai_1 _1835_ (.B1(_1002_),
    .Y(_1003_),
    .A1(net436),
    .A2(_1000_));
 sg13g2_a21oi_1 _1836_ (.A1(_0998_),
    .A2(_1001_),
    .Y(_1004_),
    .B1(_1003_));
 sg13g2_nor2_1 _1837_ (.A(_0448_),
    .B(_0999_),
    .Y(_1005_));
 sg13g2_nor4_1 _1838_ (.A(_0568_),
    .B(_0975_),
    .C(_1004_),
    .D(_1005_),
    .Y(_1006_));
 sg13g2_nor4_1 _1839_ (.A(_0778_),
    .B(_0827_),
    .C(_0860_),
    .D(_1006_),
    .Y(_1007_));
 sg13g2_nor2_1 _1840_ (.A(net407),
    .B(net410),
    .Y(_1008_));
 sg13g2_o21ai_1 _1841_ (.B1(net406),
    .Y(_1009_),
    .A1(net407),
    .A2(net410));
 sg13g2_nand4_1 _1842_ (.B(net441),
    .C(net443),
    .A(net440),
    .Y(_1010_),
    .D(net434));
 sg13g2_nand3_1 _1843_ (.B(_1009_),
    .C(_1010_),
    .A(_0329_),
    .Y(_1011_));
 sg13g2_nand3_1 _1844_ (.B(net415),
    .C(net418),
    .A(net414),
    .Y(_1012_));
 sg13g2_inv_1 _1845_ (.Y(_1013_),
    .A(_1012_));
 sg13g2_nand3_1 _1846_ (.B(net424),
    .C(net422),
    .A(net420),
    .Y(_1014_));
 sg13g2_o21ai_1 _1847_ (.B1(_1008_),
    .Y(_1015_),
    .A1(_1012_),
    .A2(_1014_));
 sg13g2_nand4_1 _1848_ (.B(_0325_),
    .C(net446),
    .A(net452),
    .Y(_1016_),
    .D(net434));
 sg13g2_nand3_1 _1849_ (.B(net440),
    .C(net441),
    .A(net449),
    .Y(_1017_));
 sg13g2_nor3_1 _1850_ (.A(_0357_),
    .B(_1016_),
    .C(_1017_),
    .Y(_1018_));
 sg13g2_nor4_1 _1851_ (.A(net440),
    .B(net441),
    .C(net443),
    .D(net446),
    .Y(_1019_));
 sg13g2_nand2_1 _1852_ (.Y(_1020_),
    .A(_0317_),
    .B(_0357_));
 sg13g2_nor3_1 _1853_ (.A(net449),
    .B(net434),
    .C(_1020_),
    .Y(_1021_));
 sg13g2_a21oi_1 _1854_ (.A1(_1019_),
    .A2(_1021_),
    .Y(_1022_),
    .B1(_1018_));
 sg13g2_nor3_1 _1855_ (.A(net414),
    .B(net415),
    .C(net418),
    .Y(_1023_));
 sg13g2_nor4_1 _1856_ (.A(net404),
    .B(net420),
    .C(net424),
    .D(net423),
    .Y(_1024_));
 sg13g2_and3_1 _1857_ (.X(_1025_),
    .A(_1008_),
    .B(_1023_),
    .C(_1024_));
 sg13g2_a21oi_2 _1858_ (.B1(_1025_),
    .Y(_1026_),
    .A2(_1015_),
    .A1(net404));
 sg13g2_nand3b_1 _1859_ (.B(_1022_),
    .C(_1026_),
    .Y(_1027_),
    .A_N(_1011_));
 sg13g2_a21oi_2 _1860_ (.B1(_1027_),
    .Y(_1028_),
    .A2(_1007_),
    .A1(_0595_));
 sg13g2_a21oi_2 _1861_ (.B1(_1011_),
    .Y(_1029_),
    .A2(_1026_),
    .A1(_1022_));
 sg13g2_nand3_1 _1862_ (.B(\color_state[2] ),
    .C(_0344_),
    .A(_0343_),
    .Y(_1030_));
 sg13g2_nand2b_1 _1863_ (.Y(_1031_),
    .B(\color_state[1] ),
    .A_N(\color_state[2] ));
 sg13g2_nand3_1 _1864_ (.B(_1030_),
    .C(_1031_),
    .A(_1029_),
    .Y(_1032_));
 sg13g2_nand2b_1 _1865_ (.Y(uo_out[0]),
    .B(_1032_),
    .A_N(_1028_));
 sg13g2_nor2_1 _1866_ (.A(_0343_),
    .B(\color_state[2] ),
    .Y(_1033_));
 sg13g2_o21ai_1 _1867_ (.B1(_1029_),
    .Y(_1034_),
    .A1(\color_state[1] ),
    .A2(_1033_));
 sg13g2_nand2b_1 _1868_ (.Y(uo_out[5]),
    .B(_1034_),
    .A_N(_1028_));
 sg13g2_a21oi_1 _1869_ (.A1(\color_state[0] ),
    .A2(\color_state[2] ),
    .Y(uo_out[1]),
    .B1(_1034_));
 sg13g2_nor2_1 _1870_ (.A(_0343_),
    .B(_0344_),
    .Y(_1035_));
 sg13g2_nor2_1 _1871_ (.A(\color_state[2] ),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_nor2b_1 _1872_ (.A(_1036_),
    .B_N(_1029_),
    .Y(uo_out[6]));
 sg13g2_nand2_1 _1873_ (.Y(_1037_),
    .A(\color_state[2] ),
    .B(_1035_));
 sg13g2_and2_1 _1874_ (.A(uo_out[6]),
    .B(_1037_),
    .X(uo_out[2]));
 sg13g2_xor2_1 _1875_ (.B(\tick_count[0] ),
    .A(\tick_count[1] ),
    .X(_0001_));
 sg13g2_nand3_1 _1876_ (.B(\tick_count[1] ),
    .C(\tick_count[0] ),
    .A(\tick_count[2] ),
    .Y(_1038_));
 sg13g2_a21o_1 _1877_ (.A2(\tick_count[0] ),
    .A1(\tick_count[1] ),
    .B1(\tick_count[2] ),
    .X(_1039_));
 sg13g2_and2_1 _1878_ (.A(_1038_),
    .B(_1039_),
    .X(_0002_));
 sg13g2_nand4_1 _1879_ (.B(\tick_count[3] ),
    .C(\tick_count[1] ),
    .A(\tick_count[2] ),
    .Y(_1040_),
    .D(\tick_count[0] ));
 sg13g2_xnor2_1 _1880_ (.Y(_0003_),
    .A(\tick_count[3] ),
    .B(_1038_));
 sg13g2_nand3_1 _1881_ (.B(net450),
    .C(_0429_),
    .A(net449),
    .Y(_1041_));
 sg13g2_nand2_1 _1882_ (.Y(_1042_),
    .A(net402),
    .B(_1041_));
 sg13g2_nor2_1 _1883_ (.A(net450),
    .B(_0429_),
    .Y(_1043_));
 sg13g2_a21oi_1 _1884_ (.A1(net434),
    .A2(_0429_),
    .Y(_1044_),
    .B1(_1043_));
 sg13g2_nand3_1 _1885_ (.B(_0329_),
    .C(_1020_),
    .A(net449),
    .Y(_1045_));
 sg13g2_nor4_1 _1886_ (.A(_1010_),
    .B(_1042_),
    .C(_1044_),
    .D(net57),
    .Y(_0005_));
 sg13g2_nand2_1 _1887_ (.Y(_1046_),
    .A(net404),
    .B(_0334_));
 sg13g2_nor4_1 _1888_ (.A(_0336_),
    .B(_1013_),
    .C(_1023_),
    .D(_1046_),
    .Y(_0004_));
 sg13g2_nor2_1 _1889_ (.A(_1032_),
    .B(_1035_),
    .Y(uo_out[4]));
 sg13g2_nor2_1 _1890_ (.A(_0343_),
    .B(_1040_),
    .Y(_1047_));
 sg13g2_xnor2_1 _1891_ (.Y(_0006_),
    .A(\color_state[0] ),
    .B(_1040_));
 sg13g2_nor3_1 _1892_ (.A(_0343_),
    .B(_0344_),
    .C(_1040_),
    .Y(_1048_));
 sg13g2_xnor2_1 _1893_ (.Y(_0007_),
    .A(_0344_),
    .B(_1047_));
 sg13g2_xor2_1 _1894_ (.B(_1048_),
    .A(\color_state[2] ),
    .X(_0008_));
 sg13g2_nand3_1 _1895_ (.B(net422),
    .C(_0617_),
    .A(net420),
    .Y(_1049_));
 sg13g2_nor2_1 _1896_ (.A(net399),
    .B(_1049_),
    .Y(_1050_));
 sg13g2_or2_1 _1897_ (.X(_1051_),
    .B(_1049_),
    .A(net399));
 sg13g2_nand3_1 _1898_ (.B(net407),
    .C(_0336_),
    .A(net404),
    .Y(_1052_));
 sg13g2_nor4_2 _1899_ (.A(net414),
    .B(net415),
    .C(_1051_),
    .Y(_1053_),
    .D(_1052_));
 sg13g2_nor4_1 _1900_ (.A(net452),
    .B(_0329_),
    .C(net437),
    .D(\hvsync_gen.vpos[0] ),
    .Y(_1054_));
 sg13g2_nand4_1 _1901_ (.B(net450),
    .C(_1019_),
    .A(net449),
    .Y(_1055_),
    .D(_1054_));
 sg13g2_nand3_1 _1902_ (.B(_1053_),
    .C(_1055_),
    .A(net462),
    .Y(_1056_));
 sg13g2_nor2b_1 _1903_ (.A(net48),
    .B_N(_1056_),
    .Y(_1057_));
 sg13g2_nor2b_2 _1904_ (.A(_1053_),
    .B_N(net457),
    .Y(_1058_));
 sg13g2_nand2b_2 _1905_ (.Y(_1059_),
    .B(net457),
    .A_N(_1053_));
 sg13g2_a21oi_1 _1906_ (.A1(net48),
    .A2(net325),
    .Y(_0009_),
    .B1(_1057_));
 sg13g2_or3_1 _1907_ (.A(_0429_),
    .B(_0431_),
    .C(net326),
    .X(_1060_));
 sg13g2_o21ai_1 _1908_ (.B1(_1060_),
    .Y(_0010_),
    .A1(_0317_),
    .A2(net325));
 sg13g2_nand2_1 _1909_ (.Y(_1061_),
    .A(net450),
    .B(_1058_));
 sg13g2_xnor2_1 _1910_ (.Y(_1062_),
    .A(net450),
    .B(_0429_));
 sg13g2_o21ai_1 _1911_ (.B1(_1061_),
    .Y(_0011_),
    .A1(net326),
    .A2(_1062_));
 sg13g2_a21o_1 _1912_ (.A2(_0429_),
    .A1(net450),
    .B1(net449),
    .X(_1063_));
 sg13g2_nand3b_1 _1913_ (.B(_1063_),
    .C(_1041_),
    .Y(_1064_),
    .A_N(_1056_));
 sg13g2_o21ai_1 _1914_ (.B1(_1064_),
    .Y(_0012_),
    .A1(_0319_),
    .A2(_1059_));
 sg13g2_nand2_1 _1915_ (.Y(_1065_),
    .A(net446),
    .B(_1058_));
 sg13g2_nor2_1 _1916_ (.A(net402),
    .B(_1041_),
    .Y(_1066_));
 sg13g2_xnor2_1 _1917_ (.Y(_1067_),
    .A(net402),
    .B(_1041_));
 sg13g2_o21ai_1 _1918_ (.B1(_1065_),
    .Y(_0013_),
    .A1(net326),
    .A2(_1067_));
 sg13g2_nand2_1 _1919_ (.Y(_1068_),
    .A(net443),
    .B(_1058_));
 sg13g2_nand2_1 _1920_ (.Y(_1069_),
    .A(net443),
    .B(_1066_));
 sg13g2_xnor2_1 _1921_ (.Y(_1070_),
    .A(net443),
    .B(_1066_));
 sg13g2_o21ai_1 _1922_ (.B1(_1068_),
    .Y(_0014_),
    .A1(net326),
    .A2(_1070_));
 sg13g2_nor2_1 _1923_ (.A(net403),
    .B(_1069_),
    .Y(_1071_));
 sg13g2_a21oi_1 _1924_ (.A1(net403),
    .A2(_1069_),
    .Y(_1072_),
    .B1(net326));
 sg13g2_nand2b_1 _1925_ (.Y(_1073_),
    .B(_1072_),
    .A_N(_1071_));
 sg13g2_o21ai_1 _1926_ (.B1(_1073_),
    .Y(_0015_),
    .A1(net403),
    .A2(_1059_));
 sg13g2_nor3_1 _1927_ (.A(_0323_),
    .B(net403),
    .C(_1069_),
    .Y(_1074_));
 sg13g2_nand2_1 _1928_ (.Y(_1075_),
    .A(net440),
    .B(_1058_));
 sg13g2_xnor2_1 _1929_ (.Y(_1076_),
    .A(net440),
    .B(_1071_));
 sg13g2_o21ai_1 _1930_ (.B1(_1075_),
    .Y(_0016_),
    .A1(net326),
    .A2(_1076_));
 sg13g2_a21oi_1 _1931_ (.A1(net434),
    .A2(_1074_),
    .Y(_1077_),
    .B1(net326));
 sg13g2_nor2_1 _1932_ (.A(_1058_),
    .B(_1077_),
    .Y(_1078_));
 sg13g2_nor2b_1 _1933_ (.A(net326),
    .B_N(_1074_),
    .Y(_1079_));
 sg13g2_nor2_1 _1934_ (.A(net434),
    .B(_1079_),
    .Y(_1080_));
 sg13g2_nor2_1 _1935_ (.A(_1078_),
    .B(_1080_),
    .Y(_0017_));
 sg13g2_nand3_1 _1936_ (.B(net434),
    .C(_1079_),
    .A(_0329_),
    .Y(_1081_));
 sg13g2_o21ai_1 _1937_ (.B1(_1081_),
    .Y(_0018_),
    .A1(_0329_),
    .A2(_1078_));
 sg13g2_nor2_1 _1938_ (.A(net47),
    .B(net325),
    .Y(_0019_));
 sg13g2_nor2_1 _1939_ (.A(net47),
    .B(net424),
    .Y(_1082_));
 sg13g2_nor3_1 _1940_ (.A(_0617_),
    .B(net325),
    .C(_1082_),
    .Y(_0020_));
 sg13g2_o21ai_1 _1941_ (.B1(net457),
    .Y(_1083_),
    .A1(net422),
    .A2(_0617_));
 sg13g2_a21oi_1 _1942_ (.A1(net422),
    .A2(_0617_),
    .Y(_0021_),
    .B1(_1083_));
 sg13g2_a21oi_1 _1943_ (.A1(net422),
    .A2(_0617_),
    .Y(_1084_),
    .B1(net420));
 sg13g2_nand2_1 _1944_ (.Y(_1085_),
    .A(net457),
    .B(_1049_));
 sg13g2_nor2_1 _1945_ (.A(_1084_),
    .B(_1085_),
    .Y(_0022_));
 sg13g2_nand2_1 _1946_ (.Y(_1086_),
    .A(net457),
    .B(_1051_));
 sg13g2_a21oi_1 _1947_ (.A1(net399),
    .A2(_1049_),
    .Y(_0023_),
    .B1(_1086_));
 sg13g2_o21ai_1 _1948_ (.B1(_1058_),
    .Y(_1087_),
    .A1(net400),
    .A2(_1051_));
 sg13g2_a21oi_1 _1949_ (.A1(net400),
    .A2(_1051_),
    .Y(_0024_),
    .B1(_1087_));
 sg13g2_a21oi_1 _1950_ (.A1(net415),
    .A2(_1050_),
    .Y(_1088_),
    .B1(net414));
 sg13g2_nor2_2 _1951_ (.A(_1012_),
    .B(_1049_),
    .Y(_1089_));
 sg13g2_nor3_1 _1952_ (.A(net325),
    .B(net61),
    .C(_1089_),
    .Y(_0025_));
 sg13g2_xnor2_1 _1953_ (.Y(_1090_),
    .A(net410),
    .B(_1089_));
 sg13g2_nor2_1 _1954_ (.A(net325),
    .B(_1090_),
    .Y(_0026_));
 sg13g2_a21oi_1 _1955_ (.A1(net410),
    .A2(_1089_),
    .Y(_1091_),
    .B1(net407));
 sg13g2_nor4_1 _1956_ (.A(_0334_),
    .B(_0336_),
    .C(_1012_),
    .D(_1049_),
    .Y(_1092_));
 sg13g2_nor3_1 _1957_ (.A(net325),
    .B(_1091_),
    .C(_1092_),
    .Y(_0027_));
 sg13g2_a21oi_1 _1958_ (.A1(net406),
    .A2(_1092_),
    .Y(_1093_),
    .B1(net325));
 sg13g2_o21ai_1 _1959_ (.B1(_1093_),
    .Y(_1094_),
    .A1(net406),
    .A2(_1092_));
 sg13g2_inv_1 _1960_ (.Y(_0028_),
    .A(_1094_));
 sg13g2_nor2_1 _1961_ (.A(\square_x_pos[5] ),
    .B(\square_x_pos[6] ),
    .Y(_1095_));
 sg13g2_or2_1 _1962_ (.X(_1096_),
    .B(\square_x_pos[6] ),
    .A(\square_x_pos[5] ));
 sg13g2_nand2_1 _1963_ (.Y(_1097_),
    .A(net8),
    .B(\square_x_pos[3] ));
 sg13g2_xnor2_1 _1964_ (.Y(_1098_),
    .A(net8),
    .B(\square_x_pos[3] ));
 sg13g2_nor2_1 _1965_ (.A(\square_x_pos[1] ),
    .B(net6),
    .Y(_1099_));
 sg13g2_nand2_1 _1966_ (.Y(_1100_),
    .A(net453),
    .B(\square_x_pos[0] ));
 sg13g2_a22oi_1 _1967_ (.Y(_1101_),
    .B1(net453),
    .B2(\square_x_pos[0] ),
    .A2(net6),
    .A1(\square_x_pos[1] ));
 sg13g2_nand2_1 _1968_ (.Y(_1102_),
    .A(net7),
    .B(\square_x_pos[2] ));
 sg13g2_xor2_1 _1969_ (.B(\square_x_pos[2] ),
    .A(net7),
    .X(_1103_));
 sg13g2_xnor2_1 _1970_ (.Y(_1104_),
    .A(net7),
    .B(\square_x_pos[2] ));
 sg13g2_or3_1 _1971_ (.A(_1099_),
    .B(_1101_),
    .C(_1104_),
    .X(_1105_));
 sg13g2_nor3_1 _1972_ (.A(_1098_),
    .B(_1099_),
    .C(_1104_),
    .Y(_1106_));
 sg13g2_nor3_1 _1973_ (.A(_1098_),
    .B(_1099_),
    .C(_1105_),
    .Y(_1107_));
 sg13g2_nor2_1 _1974_ (.A(_1098_),
    .B(_1102_),
    .Y(_1108_));
 sg13g2_o21ai_1 _1975_ (.B1(_1097_),
    .Y(_1109_),
    .A1(_1098_),
    .A2(_1102_));
 sg13g2_o21ai_1 _1976_ (.B1(\square_x_pos[4] ),
    .Y(_1110_),
    .A1(_1107_),
    .A2(_1109_));
 sg13g2_xnor2_1 _1977_ (.Y(_1111_),
    .A(_0350_),
    .B(_1110_));
 sg13g2_xnor2_1 _1978_ (.Y(_1112_),
    .A(_0349_),
    .B(_1097_));
 sg13g2_o21ai_1 _1979_ (.B1(_1104_),
    .Y(_1113_),
    .A1(_1099_),
    .A2(_1101_));
 sg13g2_xor2_1 _1980_ (.B(net6),
    .A(\square_x_pos[1] ),
    .X(_1114_));
 sg13g2_nor2_1 _1981_ (.A(net453),
    .B(\square_x_pos[0] ),
    .Y(_1115_));
 sg13g2_nand2_1 _1982_ (.Y(_1116_),
    .A(_1114_),
    .B(_1115_));
 sg13g2_o21ai_1 _1983_ (.B1(_1116_),
    .Y(_1117_),
    .A1(_1100_),
    .A2(_1114_));
 sg13g2_xor2_1 _1984_ (.B(_1102_),
    .A(_1098_),
    .X(_1118_));
 sg13g2_nand4_1 _1985_ (.B(_1113_),
    .C(_1117_),
    .A(_1105_),
    .Y(_1119_),
    .D(_1118_));
 sg13g2_nor2_1 _1986_ (.A(_1106_),
    .B(_1108_),
    .Y(_1120_));
 sg13g2_a21o_1 _1987_ (.A2(_1120_),
    .A1(_1119_),
    .B1(_1112_),
    .X(_1121_));
 sg13g2_nand3_1 _1988_ (.B(_1119_),
    .C(_1120_),
    .A(_1112_),
    .Y(_1122_));
 sg13g2_nand3_1 _1989_ (.B(_1121_),
    .C(_1122_),
    .A(_1111_),
    .Y(_1123_));
 sg13g2_nand2_1 _1990_ (.Y(_1124_),
    .A(\square_x_pos[5] ),
    .B(\square_x_pos[6] ));
 sg13g2_a21oi_1 _1991_ (.A1(_0349_),
    .A2(_1097_),
    .Y(_1125_),
    .B1(\square_x_pos[5] ));
 sg13g2_a21oi_1 _1992_ (.A1(\square_x_pos[5] ),
    .A2(\square_x_pos[6] ),
    .Y(_0071_),
    .B1(_1125_));
 sg13g2_a21o_1 _1993_ (.A2(_0071_),
    .A1(_1123_),
    .B1(_1095_),
    .X(_0072_));
 sg13g2_nand3_1 _1994_ (.B(_0352_),
    .C(_0072_),
    .A(_0351_),
    .Y(_0073_));
 sg13g2_nand3_1 _1995_ (.B(_1096_),
    .C(_1124_),
    .A(_0352_),
    .Y(_0074_));
 sg13g2_nor3_1 _1996_ (.A(_1119_),
    .B(_1123_),
    .C(_0074_),
    .Y(_0075_));
 sg13g2_o21ai_1 _1997_ (.B1(_0075_),
    .Y(_0076_),
    .A1(_0351_),
    .A2(_0072_));
 sg13g2_and4_1 _1998_ (.A(net328),
    .B(\square_x_pos[9] ),
    .C(_0073_),
    .D(_0076_),
    .X(_0077_));
 sg13g2_nor2_1 _1999_ (.A(net6),
    .B(net453),
    .Y(_0078_));
 sg13g2_nor4_2 _2000_ (.A(net6),
    .B(net453),
    .C(net7),
    .Y(_0079_),
    .D(net8));
 sg13g2_nor2b_1 _2001_ (.A(net7),
    .B_N(\square_x_pos[2] ),
    .Y(_0080_));
 sg13g2_nand2b_1 _2002_ (.Y(_0081_),
    .B(\square_x_pos[1] ),
    .A_N(net6));
 sg13g2_nand2b_2 _2003_ (.Y(_0082_),
    .B(net453),
    .A_N(\square_x_pos[0] ));
 sg13g2_nand2b_1 _2004_ (.Y(_0083_),
    .B(_0082_),
    .A_N(_1114_));
 sg13g2_a21oi_1 _2005_ (.A1(_0081_),
    .A2(_0083_),
    .Y(_0084_),
    .B1(_1103_));
 sg13g2_or2_1 _2006_ (.X(_0085_),
    .B(_0084_),
    .A(_0080_));
 sg13g2_o21ai_1 _2007_ (.B1(_1098_),
    .Y(_0086_),
    .A1(_0080_),
    .A2(_0084_));
 sg13g2_o21ai_1 _2008_ (.B1(_0086_),
    .Y(_0087_),
    .A1(net8),
    .A2(_0359_));
 sg13g2_nor2_1 _2009_ (.A(\square_x_pos[4] ),
    .B(_0087_),
    .Y(_0088_));
 sg13g2_nor4_1 _2010_ (.A(\square_x_pos[4] ),
    .B(\square_x_pos[7] ),
    .C(_1096_),
    .D(_0087_),
    .Y(_0089_));
 sg13g2_nand2_1 _2011_ (.Y(_0090_),
    .A(_0352_),
    .B(_0089_));
 sg13g2_nor2_1 _2012_ (.A(\square_x_pos[9] ),
    .B(_0090_),
    .Y(_0091_));
 sg13g2_a21oi_1 _2013_ (.A1(net346),
    .A2(_0091_),
    .Y(_0092_),
    .B1(_0079_));
 sg13g2_nor2b_2 _2014_ (.A(_0077_),
    .B_N(_0092_),
    .Y(_0093_));
 sg13g2_nand2_1 _2015_ (.Y(_0094_),
    .A(net453),
    .B(net320));
 sg13g2_nor2b_2 _2016_ (.A(net397),
    .B_N(net453),
    .Y(_0095_));
 sg13g2_and2_1 _2017_ (.A(net321),
    .B(_0095_),
    .X(_0096_));
 sg13g2_a21o_1 _2018_ (.A2(_0094_),
    .A1(net397),
    .B1(_0096_),
    .X(_0029_));
 sg13g2_nor2_1 _2019_ (.A(net393),
    .B(net320),
    .Y(_0097_));
 sg13g2_nor2b_2 _2020_ (.A(net345),
    .B_N(net5),
    .Y(_0098_));
 sg13g2_xnor2_1 _2021_ (.Y(_0099_),
    .A(net6),
    .B(_0098_));
 sg13g2_nand2_1 _2022_ (.Y(_0100_),
    .A(net394),
    .B(_0099_));
 sg13g2_nor2_1 _2023_ (.A(net394),
    .B(_0099_),
    .Y(_0101_));
 sg13g2_xnor2_1 _2024_ (.Y(_0102_),
    .A(net394),
    .B(_0099_));
 sg13g2_xnor2_1 _2025_ (.Y(_0103_),
    .A(_0095_),
    .B(_0102_));
 sg13g2_a21oi_1 _2026_ (.A1(net321),
    .A2(_0103_),
    .Y(_0030_),
    .B1(_0097_));
 sg13g2_nor2_1 _2027_ (.A(net345),
    .B(_0078_),
    .Y(_0104_));
 sg13g2_xnor2_1 _2028_ (.Y(_0105_),
    .A(net7),
    .B(_0104_));
 sg13g2_and2_1 _2029_ (.A(net388),
    .B(_0105_),
    .X(_0106_));
 sg13g2_xor2_1 _2030_ (.B(_0105_),
    .A(net389),
    .X(_0107_));
 sg13g2_o21ai_1 _2031_ (.B1(_0100_),
    .Y(_0108_),
    .A1(_0095_),
    .A2(_0101_));
 sg13g2_xnor2_1 _2032_ (.Y(_0109_),
    .A(_0107_),
    .B(_0108_));
 sg13g2_nor2_1 _2033_ (.A(net389),
    .B(net321),
    .Y(_0110_));
 sg13g2_a21oi_1 _2034_ (.A1(net321),
    .A2(_0109_),
    .Y(_0031_),
    .B1(_0110_));
 sg13g2_a21oi_1 _2035_ (.A1(_0358_),
    .A2(_0078_),
    .Y(_0111_),
    .B1(net345));
 sg13g2_xnor2_1 _2036_ (.Y(_0112_),
    .A(net8),
    .B(_0111_));
 sg13g2_nand2_1 _2037_ (.Y(_0113_),
    .A(net384),
    .B(_0112_));
 sg13g2_xnor2_1 _2038_ (.Y(_0114_),
    .A(net384),
    .B(_0112_));
 sg13g2_a21oi_1 _2039_ (.A1(_0107_),
    .A2(_0108_),
    .Y(_0115_),
    .B1(_0106_));
 sg13g2_xnor2_1 _2040_ (.Y(_0116_),
    .A(_0114_),
    .B(_0115_));
 sg13g2_nor2_1 _2041_ (.A(net385),
    .B(net320),
    .Y(_0117_));
 sg13g2_a21oi_1 _2042_ (.A1(net320),
    .A2(_0116_),
    .Y(_0032_),
    .B1(_0117_));
 sg13g2_nor2_1 _2043_ (.A(net380),
    .B(net320),
    .Y(_0118_));
 sg13g2_nor2_2 _2044_ (.A(net345),
    .B(_0079_),
    .Y(_0119_));
 sg13g2_or2_1 _2045_ (.X(_0120_),
    .B(_0079_),
    .A(net345));
 sg13g2_nor2_1 _2046_ (.A(net335),
    .B(net327),
    .Y(_0121_));
 sg13g2_xnor2_1 _2047_ (.Y(_0122_),
    .A(net380),
    .B(net327));
 sg13g2_o21ai_1 _2048_ (.B1(_0113_),
    .Y(_0123_),
    .A1(_0114_),
    .A2(_0115_));
 sg13g2_xnor2_1 _2049_ (.Y(_0124_),
    .A(_0122_),
    .B(_0123_));
 sg13g2_a21oi_1 _2050_ (.A1(net320),
    .A2(_0124_),
    .Y(_0033_),
    .B1(_0118_));
 sg13g2_xnor2_1 _2051_ (.Y(_0125_),
    .A(net378),
    .B(net327));
 sg13g2_a21oi_1 _2052_ (.A1(_0122_),
    .A2(_0123_),
    .Y(_0126_),
    .B1(_0121_));
 sg13g2_xnor2_1 _2053_ (.Y(_0127_),
    .A(_0125_),
    .B(_0126_));
 sg13g2_nand2_1 _2054_ (.Y(_0128_),
    .A(net320),
    .B(_0127_));
 sg13g2_o21ai_1 _2055_ (.B1(_0128_),
    .Y(_0034_),
    .A1(net338),
    .A2(net320));
 sg13g2_nor2_1 _2056_ (.A(net331),
    .B(net327),
    .Y(_0129_));
 sg13g2_xnor2_1 _2057_ (.Y(_0130_),
    .A(net374),
    .B(net327));
 sg13g2_o21ai_1 _2058_ (.B1(_0120_),
    .Y(_0131_),
    .A1(net378),
    .A2(net380));
 sg13g2_nand3_1 _2059_ (.B(_0123_),
    .C(_0125_),
    .A(_0122_),
    .Y(_0132_));
 sg13g2_nand2_1 _2060_ (.Y(_0133_),
    .A(_0131_),
    .B(_0132_));
 sg13g2_xor2_1 _2061_ (.B(_0133_),
    .A(_0130_),
    .X(_0134_));
 sg13g2_nand2_1 _2062_ (.Y(_0135_),
    .A(net322),
    .B(_0134_));
 sg13g2_o21ai_1 _2063_ (.B1(_0135_),
    .Y(_0035_),
    .A1(net331),
    .A2(net322));
 sg13g2_xnor2_1 _2064_ (.Y(_0136_),
    .A(net373),
    .B(_0119_));
 sg13g2_a21oi_1 _2065_ (.A1(_0130_),
    .A2(_0133_),
    .Y(_0137_),
    .B1(_0129_));
 sg13g2_xnor2_1 _2066_ (.Y(_0138_),
    .A(_0136_),
    .B(_0137_));
 sg13g2_nand2_1 _2067_ (.Y(_0139_),
    .A(net322),
    .B(_0138_));
 sg13g2_o21ai_1 _2068_ (.B1(_0139_),
    .Y(_0036_),
    .A1(net329),
    .A2(net322));
 sg13g2_nor2_1 _2069_ (.A(net333),
    .B(net327),
    .Y(_0140_));
 sg13g2_xnor2_1 _2070_ (.Y(_0141_),
    .A(net372),
    .B(net327));
 sg13g2_nand2_1 _2071_ (.Y(_0142_),
    .A(_0130_),
    .B(_0136_));
 sg13g2_o21ai_1 _2072_ (.B1(_0120_),
    .Y(_0143_),
    .A1(net374),
    .A2(net373));
 sg13g2_and2_1 _2073_ (.A(_0131_),
    .B(_0143_),
    .X(_0144_));
 sg13g2_o21ai_1 _2074_ (.B1(_0144_),
    .Y(_0145_),
    .A1(_0132_),
    .A2(_0142_));
 sg13g2_xnor2_1 _2075_ (.Y(_0146_),
    .A(_0141_),
    .B(_0145_));
 sg13g2_nor2_1 _2076_ (.A(net371),
    .B(net324),
    .Y(_0147_));
 sg13g2_a21oi_1 _2077_ (.A1(net324),
    .A2(_0146_),
    .Y(_0037_),
    .B1(_0147_));
 sg13g2_a21oi_1 _2078_ (.A1(_0141_),
    .A2(_0145_),
    .Y(_0148_),
    .B1(_0140_));
 sg13g2_xnor2_1 _2079_ (.Y(_0149_),
    .A(\dog_pos_x[9] ),
    .B(net327));
 sg13g2_xnor2_1 _2080_ (.Y(_0150_),
    .A(_0148_),
    .B(_0149_));
 sg13g2_nand2_1 _2081_ (.Y(_0151_),
    .A(net324),
    .B(_0150_));
 sg13g2_o21ai_1 _2082_ (.B1(_0151_),
    .Y(_0038_),
    .A1(_0341_),
    .A2(net324));
 sg13g2_nand2_1 _2083_ (.Y(_0152_),
    .A(net3),
    .B(\square_y_pos[2] ));
 sg13g2_xor2_1 _2084_ (.B(\square_y_pos[2] ),
    .A(net3),
    .X(_0153_));
 sg13g2_nor2_1 _2085_ (.A(\square_y_pos[1] ),
    .B(net2),
    .Y(_0154_));
 sg13g2_nand2_1 _2086_ (.Y(_0155_),
    .A(\square_y_pos[1] ),
    .B(net2));
 sg13g2_nand2_1 _2087_ (.Y(_0156_),
    .A(net1),
    .B(\square_y_pos[0] ));
 sg13g2_o21ai_1 _2088_ (.B1(_0155_),
    .Y(_0157_),
    .A1(_0154_),
    .A2(_0156_));
 sg13g2_nand2_1 _2089_ (.Y(_0158_),
    .A(_0153_),
    .B(_0157_));
 sg13g2_xnor2_1 _2090_ (.Y(_0159_),
    .A(_0153_),
    .B(_0157_));
 sg13g2_nand2_1 _2091_ (.Y(_0160_),
    .A(net4),
    .B(\square_y_pos[3] ));
 sg13g2_xor2_1 _2092_ (.B(\square_y_pos[3] ),
    .A(net4),
    .X(_0161_));
 sg13g2_xnor2_1 _2093_ (.Y(_0162_),
    .A(net4),
    .B(\square_y_pos[3] ));
 sg13g2_nand2b_1 _2094_ (.Y(_0163_),
    .B(_0161_),
    .A_N(_0152_));
 sg13g2_xnor2_1 _2095_ (.Y(_0164_),
    .A(\square_y_pos[1] ),
    .B(net2));
 sg13g2_a22oi_1 _2096_ (.Y(_0165_),
    .B1(_0164_),
    .B2(_0156_),
    .A2(_0162_),
    .A1(_0152_));
 sg13g2_nand2_1 _2097_ (.Y(_0166_),
    .A(_0163_),
    .B(_0165_));
 sg13g2_nand2_1 _2098_ (.Y(_0167_),
    .A(\square_y_pos[4] ),
    .B(_0160_));
 sg13g2_a21oi_1 _2099_ (.A1(_0353_),
    .A2(_0360_),
    .Y(_0168_),
    .B1(_0164_));
 sg13g2_nand3b_1 _2100_ (.B(_0161_),
    .C(_0153_),
    .Y(_0169_),
    .A_N(_0154_));
 sg13g2_or2_1 _2101_ (.X(_0170_),
    .B(_0160_),
    .A(\square_y_pos[4] ));
 sg13g2_nand3_1 _2102_ (.B(_0169_),
    .C(_0170_),
    .A(_0163_),
    .Y(_0171_));
 sg13g2_nor3_1 _2103_ (.A(_0159_),
    .B(_0166_),
    .C(_0168_),
    .Y(_0172_));
 sg13g2_o21ai_1 _2104_ (.B1(_0167_),
    .Y(_0173_),
    .A1(_0171_),
    .A2(_0172_));
 sg13g2_nor2_1 _2105_ (.A(\square_y_pos[4] ),
    .B(\square_y_pos[5] ),
    .Y(_0174_));
 sg13g2_and2_1 _2106_ (.A(\square_y_pos[4] ),
    .B(\square_y_pos[5] ),
    .X(_0175_));
 sg13g2_nor2_1 _2107_ (.A(_0174_),
    .B(_0175_),
    .Y(_0176_));
 sg13g2_nor3_2 _2108_ (.A(\square_y_pos[4] ),
    .B(\square_y_pos[5] ),
    .C(\square_y_pos[6] ),
    .Y(_0177_));
 sg13g2_and2_1 _2109_ (.A(_0167_),
    .B(_0170_),
    .X(_0178_));
 sg13g2_a221oi_1 _2110_ (.B2(_0172_),
    .C1(_0177_),
    .B1(_0178_),
    .A1(_0173_),
    .Y(_0179_),
    .A2(_0176_));
 sg13g2_o21ai_1 _2111_ (.B1(\square_y_pos[6] ),
    .Y(_0180_),
    .A1(\square_y_pos[4] ),
    .A2(\square_y_pos[5] ));
 sg13g2_o21ai_1 _2112_ (.B1(_0180_),
    .Y(_0181_),
    .A1(_0173_),
    .A2(_0176_));
 sg13g2_or2_1 _2113_ (.X(_0182_),
    .B(_0181_),
    .A(_0179_));
 sg13g2_nand2b_1 _2114_ (.Y(_0183_),
    .B(_0177_),
    .A_N(_0173_));
 sg13g2_nand4_1 _2115_ (.B(\square_y_pos[8] ),
    .C(_0182_),
    .A(\square_y_pos[7] ),
    .Y(_0184_),
    .D(_0183_));
 sg13g2_a21oi_1 _2116_ (.A1(_0348_),
    .A2(_0184_),
    .Y(_0185_),
    .B1(net344));
 sg13g2_nand2b_1 _2117_ (.Y(_0186_),
    .B(\square_y_pos[2] ),
    .A_N(net3));
 sg13g2_nand2_1 _2118_ (.Y(_0187_),
    .A(\square_y_pos[1] ),
    .B(_0347_));
 sg13g2_nand2_1 _2119_ (.Y(_0188_),
    .A(net1),
    .B(_0360_));
 sg13g2_nand2_1 _2120_ (.Y(_0189_),
    .A(_0164_),
    .B(_0188_));
 sg13g2_a21o_1 _2121_ (.A2(_0189_),
    .A1(_0187_),
    .B1(_0153_),
    .X(_0190_));
 sg13g2_and2_1 _2122_ (.A(_0186_),
    .B(_0190_),
    .X(_0191_));
 sg13g2_nor2_1 _2123_ (.A(_0161_),
    .B(_0191_),
    .Y(_0192_));
 sg13g2_a21oi_1 _2124_ (.A1(_0354_),
    .A2(\square_y_pos[3] ),
    .Y(_0193_),
    .B1(_0192_));
 sg13g2_nand2_1 _2125_ (.Y(_0194_),
    .A(_0177_),
    .B(_0193_));
 sg13g2_nor4_1 _2126_ (.A(\square_y_pos[7] ),
    .B(\square_y_pos[8] ),
    .C(\square_y_pos[9] ),
    .D(_0194_),
    .Y(_0195_));
 sg13g2_a21o_2 _2127_ (.A2(_0195_),
    .A1(net344),
    .B1(_0185_),
    .X(_0196_));
 sg13g2_o21ai_1 _2128_ (.B1(net370),
    .Y(_0197_),
    .A1(_0353_),
    .A2(net319));
 sg13g2_nand2b_2 _2129_ (.Y(_0198_),
    .B(net1),
    .A_N(net370));
 sg13g2_o21ai_1 _2130_ (.B1(_0197_),
    .Y(_0039_),
    .A1(net319),
    .A2(_0198_));
 sg13g2_nand2_1 _2131_ (.Y(_0199_),
    .A(net367),
    .B(net316));
 sg13g2_nor2b_2 _2132_ (.A(net343),
    .B_N(net1),
    .Y(_0200_));
 sg13g2_xnor2_1 _2133_ (.Y(_0201_),
    .A(net2),
    .B(_0200_));
 sg13g2_and2_1 _2134_ (.A(net367),
    .B(_0201_),
    .X(_0202_));
 sg13g2_xor2_1 _2135_ (.B(_0201_),
    .A(net367),
    .X(_0203_));
 sg13g2_xnor2_1 _2136_ (.Y(_0204_),
    .A(_0198_),
    .B(_0203_));
 sg13g2_o21ai_1 _2137_ (.B1(_0199_),
    .Y(_0040_),
    .A1(net316),
    .A2(_0204_));
 sg13g2_a21oi_1 _2138_ (.A1(_0347_),
    .A2(_0353_),
    .Y(_0205_),
    .B1(net343));
 sg13g2_xnor2_1 _2139_ (.Y(_0206_),
    .A(net3),
    .B(_0205_));
 sg13g2_and2_1 _2140_ (.A(net363),
    .B(_0206_),
    .X(_0207_));
 sg13g2_xor2_1 _2141_ (.B(_0206_),
    .A(net363),
    .X(_0208_));
 sg13g2_a21o_1 _2142_ (.A2(_0203_),
    .A1(_0198_),
    .B1(_0202_),
    .X(_0209_));
 sg13g2_xnor2_1 _2143_ (.Y(_0210_),
    .A(_0208_),
    .B(_0209_));
 sg13g2_nand2_1 _2144_ (.Y(_0211_),
    .A(net363),
    .B(net316));
 sg13g2_o21ai_1 _2145_ (.B1(_0211_),
    .Y(_0041_),
    .A1(net316),
    .A2(_0210_));
 sg13g2_nor3_1 _2146_ (.A(net2),
    .B(net1),
    .C(net3),
    .Y(_0212_));
 sg13g2_nor2_1 _2147_ (.A(net343),
    .B(_0212_),
    .Y(_0213_));
 sg13g2_xnor2_1 _2148_ (.Y(_0214_),
    .A(net4),
    .B(_0213_));
 sg13g2_nand2_1 _2149_ (.Y(_0215_),
    .A(net359),
    .B(_0214_));
 sg13g2_nor2_1 _2150_ (.A(net359),
    .B(_0214_),
    .Y(_0216_));
 sg13g2_xnor2_1 _2151_ (.Y(_0217_),
    .A(_0318_),
    .B(_0214_));
 sg13g2_a21oi_1 _2152_ (.A1(_0208_),
    .A2(_0209_),
    .Y(_0218_),
    .B1(_0207_));
 sg13g2_xnor2_1 _2153_ (.Y(_0219_),
    .A(_0217_),
    .B(_0218_));
 sg13g2_nor2_1 _2154_ (.A(net315),
    .B(_0219_),
    .Y(_0220_));
 sg13g2_a21oi_1 _2155_ (.A1(_0318_),
    .A2(net315),
    .Y(_0042_),
    .B1(_0220_));
 sg13g2_and2_1 _2156_ (.A(_0354_),
    .B(_0212_),
    .X(_0221_));
 sg13g2_nor2_2 _2157_ (.A(net344),
    .B(_0221_),
    .Y(_0222_));
 sg13g2_or2_1 _2158_ (.X(_0223_),
    .B(_0221_),
    .A(net344));
 sg13g2_xnor2_1 _2159_ (.Y(_0224_),
    .A(net356),
    .B(_0222_));
 sg13g2_o21ai_1 _2160_ (.B1(_0215_),
    .Y(_0225_),
    .A1(_0216_),
    .A2(_0218_));
 sg13g2_and2_1 _2161_ (.A(_0224_),
    .B(_0225_),
    .X(_0226_));
 sg13g2_xor2_1 _2162_ (.B(_0225_),
    .A(_0224_),
    .X(_0227_));
 sg13g2_nor2_1 _2163_ (.A(net315),
    .B(_0227_),
    .Y(_0228_));
 sg13g2_a21oi_1 _2164_ (.A1(net340),
    .A2(net315),
    .Y(_0043_),
    .B1(_0228_));
 sg13g2_xnor2_1 _2165_ (.Y(_0229_),
    .A(net354),
    .B(_0222_));
 sg13g2_a21oi_1 _2166_ (.A1(net356),
    .A2(_0223_),
    .Y(_0230_),
    .B1(_0226_));
 sg13g2_xnor2_1 _2167_ (.Y(_0231_),
    .A(_0229_),
    .B(_0230_));
 sg13g2_nor2_1 _2168_ (.A(net315),
    .B(_0231_),
    .Y(_0232_));
 sg13g2_a21oi_1 _2169_ (.A1(net342),
    .A2(net315),
    .Y(_0044_),
    .B1(_0232_));
 sg13g2_nor2_1 _2170_ (.A(net341),
    .B(_0222_),
    .Y(_0233_));
 sg13g2_xnor2_1 _2171_ (.Y(_0234_),
    .A(net352),
    .B(_0222_));
 sg13g2_nand2_1 _2172_ (.Y(_0235_),
    .A(_0226_),
    .B(_0229_));
 sg13g2_o21ai_1 _2173_ (.B1(_0223_),
    .Y(_0236_),
    .A1(net354),
    .A2(net356));
 sg13g2_nand2_1 _2174_ (.Y(_0237_),
    .A(_0235_),
    .B(_0236_));
 sg13g2_xor2_1 _2175_ (.B(_0237_),
    .A(_0234_),
    .X(_0238_));
 sg13g2_nor2_1 _2176_ (.A(net315),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_a21oi_1 _2177_ (.A1(net341),
    .A2(net315),
    .Y(_0045_),
    .B1(_0239_));
 sg13g2_xnor2_1 _2178_ (.Y(_0240_),
    .A(net351),
    .B(_0222_));
 sg13g2_a21oi_1 _2179_ (.A1(_0234_),
    .A2(_0237_),
    .Y(_0241_),
    .B1(_0233_));
 sg13g2_or2_1 _2180_ (.X(_0242_),
    .B(_0241_),
    .A(_0240_));
 sg13g2_a21oi_1 _2181_ (.A1(_0240_),
    .A2(_0241_),
    .Y(_0243_),
    .B1(net317));
 sg13g2_a22oi_1 _2182_ (.Y(_0046_),
    .B1(_0242_),
    .B2(_0243_),
    .A2(net317),
    .A1(_0328_));
 sg13g2_xnor2_1 _2183_ (.Y(_0244_),
    .A(_0327_),
    .B(_0222_));
 sg13g2_nand4_1 _2184_ (.B(_0229_),
    .C(_0234_),
    .A(_0226_),
    .Y(_0245_),
    .D(_0240_));
 sg13g2_o21ai_1 _2185_ (.B1(_0223_),
    .Y(_0246_),
    .A1(net352),
    .A2(net351));
 sg13g2_and2_1 _2186_ (.A(_0236_),
    .B(_0246_),
    .X(_0247_));
 sg13g2_and3_1 _2187_ (.X(_0248_),
    .A(_0244_),
    .B(_0245_),
    .C(_0247_));
 sg13g2_a21oi_1 _2188_ (.A1(_0245_),
    .A2(_0247_),
    .Y(_0249_),
    .B1(_0244_));
 sg13g2_nor3_1 _2189_ (.A(net317),
    .B(_0248_),
    .C(_0249_),
    .Y(_0250_));
 sg13g2_a21o_1 _2190_ (.A2(net317),
    .A1(net347),
    .B1(_0250_),
    .X(_0047_));
 sg13g2_a21oi_1 _2191_ (.A1(net348),
    .A2(_0223_),
    .Y(_0251_),
    .B1(_0249_));
 sg13g2_xnor2_1 _2192_ (.Y(_0252_),
    .A(\dog_pos_y[9] ),
    .B(_0222_));
 sg13g2_xnor2_1 _2193_ (.Y(_0253_),
    .A(_0251_),
    .B(_0252_));
 sg13g2_mux2_1 _2194_ (.A0(_0253_),
    .A1(\dog_pos_y[9] ),
    .S(net317),
    .X(_0048_));
 sg13g2_nor2b_1 _2195_ (.A(_0082_),
    .B_N(net322),
    .Y(_0254_));
 sg13g2_a21o_1 _2196_ (.A2(_0094_),
    .A1(\square_x_pos[0] ),
    .B1(_0254_),
    .X(_0049_));
 sg13g2_nor2_1 _2197_ (.A(\square_x_pos[1] ),
    .B(net324),
    .Y(_0255_));
 sg13g2_xnor2_1 _2198_ (.Y(_0256_),
    .A(_1114_),
    .B(_0082_));
 sg13g2_xnor2_1 _2199_ (.Y(_0257_),
    .A(_0098_),
    .B(_0256_));
 sg13g2_a21oi_1 _2200_ (.A1(net324),
    .A2(_0257_),
    .Y(_0050_),
    .B1(_0255_));
 sg13g2_nand3_1 _2201_ (.B(_1105_),
    .C(_1113_),
    .A(net328),
    .Y(_0258_));
 sg13g2_nand3_1 _2202_ (.B(_0081_),
    .C(_0083_),
    .A(_1103_),
    .Y(_0259_));
 sg13g2_nand3b_1 _2203_ (.B(_0259_),
    .C(net346),
    .Y(_0260_),
    .A_N(_0084_));
 sg13g2_nand2_1 _2204_ (.Y(_0261_),
    .A(_0258_),
    .B(_0260_));
 sg13g2_mux2_1 _2205_ (.A0(\square_x_pos[2] ),
    .A1(_0261_),
    .S(_0093_),
    .X(_0051_));
 sg13g2_a21oi_1 _2206_ (.A1(net7),
    .A2(\square_x_pos[2] ),
    .Y(_0262_),
    .B1(net346));
 sg13g2_a22oi_1 _2207_ (.Y(_0263_),
    .B1(_0262_),
    .B2(_1105_),
    .A2(_0085_),
    .A1(net346));
 sg13g2_xnor2_1 _2208_ (.Y(_0264_),
    .A(_1098_),
    .B(_0263_));
 sg13g2_nand2_1 _2209_ (.Y(_0265_),
    .A(net323),
    .B(_0264_));
 sg13g2_o21ai_1 _2210_ (.B1(_0265_),
    .Y(_0052_),
    .A1(_0359_),
    .A2(net324));
 sg13g2_o21ai_1 _2211_ (.B1(net328),
    .Y(_0266_),
    .A1(_1107_),
    .A2(_1109_));
 sg13g2_o21ai_1 _2212_ (.B1(_0266_),
    .Y(_0267_),
    .A1(net328),
    .A2(_0087_));
 sg13g2_nand2_1 _2213_ (.Y(_0268_),
    .A(net323),
    .B(_0267_));
 sg13g2_xnor2_1 _2214_ (.Y(_0053_),
    .A(\square_x_pos[4] ),
    .B(_0268_));
 sg13g2_o21ai_1 _2215_ (.B1(\square_x_pos[5] ),
    .Y(_0269_),
    .A1(\square_x_pos[4] ),
    .A2(_0087_));
 sg13g2_a21oi_1 _2216_ (.A1(_0350_),
    .A2(_0088_),
    .Y(_0270_),
    .B1(net328));
 sg13g2_a22oi_1 _2217_ (.Y(_0271_),
    .B1(_0269_),
    .B2(_0270_),
    .A2(_1111_),
    .A1(net328));
 sg13g2_nand2_1 _2218_ (.Y(_0272_),
    .A(net323),
    .B(_0271_));
 sg13g2_o21ai_1 _2219_ (.B1(_0272_),
    .Y(_0054_),
    .A1(_0350_),
    .A2(net323));
 sg13g2_o21ai_1 _2220_ (.B1(_0346_),
    .Y(_0273_),
    .A1(_0350_),
    .A2(_1110_));
 sg13g2_nand3b_1 _2221_ (.B(_0273_),
    .C(net323),
    .Y(_0274_),
    .A_N(_0270_));
 sg13g2_xnor2_1 _2222_ (.Y(_0055_),
    .A(\square_x_pos[6] ),
    .B(_0274_));
 sg13g2_nor3_1 _2223_ (.A(net345),
    .B(_1110_),
    .C(_1124_),
    .Y(_0275_));
 sg13g2_nand3_1 _2224_ (.B(_1095_),
    .C(_0088_),
    .A(net345),
    .Y(_0276_));
 sg13g2_nand2b_1 _2225_ (.Y(_0277_),
    .B(_0276_),
    .A_N(_0275_));
 sg13g2_nand2_1 _2226_ (.Y(_0278_),
    .A(net323),
    .B(_0277_));
 sg13g2_xnor2_1 _2227_ (.Y(_0056_),
    .A(\square_x_pos[7] ),
    .B(_0278_));
 sg13g2_nand2_1 _2228_ (.Y(_0279_),
    .A(\square_x_pos[7] ),
    .B(_0275_));
 sg13g2_a22oi_1 _2229_ (.Y(_0280_),
    .B1(_0275_),
    .B2(\square_x_pos[7] ),
    .A2(_0089_),
    .A1(net346));
 sg13g2_nor2b_1 _2230_ (.A(_0280_),
    .B_N(net323),
    .Y(_0281_));
 sg13g2_xnor2_1 _2231_ (.Y(_0057_),
    .A(_0352_),
    .B(_0281_));
 sg13g2_a22oi_1 _2232_ (.Y(_0282_),
    .B1(_0090_),
    .B2(_0279_),
    .A2(_0352_),
    .A1(net328));
 sg13g2_nand2_1 _2233_ (.Y(_0283_),
    .A(net323),
    .B(_0282_));
 sg13g2_xnor2_1 _2234_ (.Y(_0058_),
    .A(\square_x_pos[9] ),
    .B(_0283_));
 sg13g2_o21ai_1 _2235_ (.B1(\square_y_pos[0] ),
    .Y(_0284_),
    .A1(_0353_),
    .A2(net319));
 sg13g2_o21ai_1 _2236_ (.B1(_0284_),
    .Y(_0059_),
    .A1(_0188_),
    .A2(net319));
 sg13g2_xor2_1 _2237_ (.B(_0188_),
    .A(_0164_),
    .X(_0285_));
 sg13g2_xnor2_1 _2238_ (.Y(_0286_),
    .A(_0200_),
    .B(_0285_));
 sg13g2_nand2_1 _2239_ (.Y(_0287_),
    .A(\square_y_pos[1] ),
    .B(net319));
 sg13g2_o21ai_1 _2240_ (.B1(_0287_),
    .Y(_0060_),
    .A1(net319),
    .A2(_0286_));
 sg13g2_nand3_1 _2241_ (.B(_0187_),
    .C(_0189_),
    .A(_0153_),
    .Y(_0288_));
 sg13g2_nand3_1 _2242_ (.B(_0190_),
    .C(_0288_),
    .A(net343),
    .Y(_0289_));
 sg13g2_o21ai_1 _2243_ (.B1(_0289_),
    .Y(_0290_),
    .A1(net344),
    .A2(_0159_));
 sg13g2_mux2_1 _2244_ (.A0(_0290_),
    .A1(\square_y_pos[2] ),
    .S(net319),
    .X(_0061_));
 sg13g2_a21oi_1 _2245_ (.A1(_0152_),
    .A2(_0158_),
    .Y(_0291_),
    .B1(net344));
 sg13g2_a21oi_1 _2246_ (.A1(net343),
    .A2(_0191_),
    .Y(_0292_),
    .B1(_0291_));
 sg13g2_xnor2_1 _2247_ (.Y(_0293_),
    .A(_0162_),
    .B(_0292_));
 sg13g2_nand2_1 _2248_ (.Y(_0294_),
    .A(\square_y_pos[3] ),
    .B(net318));
 sg13g2_o21ai_1 _2249_ (.B1(_0294_),
    .Y(_0062_),
    .A1(net318),
    .A2(_0293_));
 sg13g2_and2_1 _2250_ (.A(net343),
    .B(_0193_),
    .X(_0295_));
 sg13g2_nand2_1 _2251_ (.Y(_0296_),
    .A(net343),
    .B(_0193_));
 sg13g2_o21ai_1 _2252_ (.B1(_0291_),
    .Y(_0297_),
    .A1(net4),
    .A2(\square_y_pos[3] ));
 sg13g2_o21ai_1 _2253_ (.B1(_0297_),
    .Y(_0298_),
    .A1(net343),
    .A2(_0160_));
 sg13g2_inv_1 _2254_ (.Y(_0299_),
    .A(_0298_));
 sg13g2_a21oi_1 _2255_ (.A1(_0296_),
    .A2(_0299_),
    .Y(_0300_),
    .B1(net318));
 sg13g2_xor2_1 _2256_ (.B(_0300_),
    .A(\square_y_pos[4] ),
    .X(_0063_));
 sg13g2_a21oi_1 _2257_ (.A1(_0175_),
    .A2(_0298_),
    .Y(_0301_),
    .B1(_0295_));
 sg13g2_o21ai_1 _2258_ (.B1(\square_y_pos[5] ),
    .Y(_0302_),
    .A1(net318),
    .A2(_0301_));
 sg13g2_nor2_1 _2259_ (.A(_0176_),
    .B(_0296_),
    .Y(_0303_));
 sg13g2_nor2_1 _2260_ (.A(\square_y_pos[5] ),
    .B(_0299_),
    .Y(_0304_));
 sg13g2_a21oi_1 _2261_ (.A1(\square_y_pos[4] ),
    .A2(_0304_),
    .Y(_0305_),
    .B1(_0303_));
 sg13g2_o21ai_1 _2262_ (.B1(_0302_),
    .Y(_0064_),
    .A1(net318),
    .A2(_0305_));
 sg13g2_nor2_1 _2263_ (.A(_0345_),
    .B(_0174_),
    .Y(_0306_));
 sg13g2_nor3_1 _2264_ (.A(net318),
    .B(_0301_),
    .C(_0306_),
    .Y(_0307_));
 sg13g2_xor2_1 _2265_ (.B(_0307_),
    .A(\square_y_pos[6] ),
    .X(_0065_));
 sg13g2_nand2_1 _2266_ (.Y(_0308_),
    .A(_0177_),
    .B(_0295_));
 sg13g2_nand3_1 _2267_ (.B(_0175_),
    .C(_0298_),
    .A(\square_y_pos[6] ),
    .Y(_0309_));
 sg13g2_a21oi_1 _2268_ (.A1(_0308_),
    .A2(_0309_),
    .Y(_0310_),
    .B1(net318));
 sg13g2_xor2_1 _2269_ (.B(_0310_),
    .A(\square_y_pos[7] ),
    .X(_0066_));
 sg13g2_or2_1 _2270_ (.X(_0311_),
    .B(_0308_),
    .A(\square_y_pos[7] ));
 sg13g2_nand4_1 _2271_ (.B(\square_y_pos[7] ),
    .C(_0175_),
    .A(\square_y_pos[6] ),
    .Y(_0312_),
    .D(_0298_));
 sg13g2_a21oi_1 _2272_ (.A1(_0311_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(net318));
 sg13g2_xor2_1 _2273_ (.B(_0313_),
    .A(\square_y_pos[8] ),
    .X(_0067_));
 sg13g2_nor2_1 _2274_ (.A(\square_y_pos[8] ),
    .B(_0311_),
    .Y(_0314_));
 sg13g2_nor2_1 _2275_ (.A(_0348_),
    .B(_0314_),
    .Y(_0068_));
 sg13g2_nand2b_1 _2276_ (.Y(_0315_),
    .B(_0077_),
    .A_N(_0079_));
 sg13g2_o21ai_1 _2277_ (.B1(_0315_),
    .Y(_0069_),
    .A1(net328),
    .A2(_0091_));
 sg13g2_nand2b_1 _2278_ (.Y(_0316_),
    .B(_0185_),
    .A_N(_0221_));
 sg13g2_o21ai_1 _2279_ (.B1(_0316_),
    .Y(_0070_),
    .A1(_0345_),
    .A2(_0195_));
 sg13g2_dfrbpq_1 _2280_ (.RESET_B(net29),
    .D(net66),
    .Q(hsync),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _2281_ (.RESET_B(net455),
    .D(_0006_),
    .Q(\color_state[0] ),
    .CLK(net427));
 sg13g2_dfrbpq_1 _2282_ (.RESET_B(net456),
    .D(_0007_),
    .Q(\color_state[1] ),
    .CLK(net428));
 sg13g2_dfrbpq_2 _2283_ (.RESET_B(net456),
    .D(_0008_),
    .Q(\color_state[2] ),
    .CLK(\hvsync_gen.vsync ));
 sg13g2_dfrbpq_2 _2284_ (.RESET_B(net45),
    .D(_0009_),
    .Q(\hvsync_gen.vpos[0] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _2285_ (.RESET_B(net44),
    .D(net63),
    .Q(\hvsync_gen.vpos[1] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _2286_ (.RESET_B(net43),
    .D(net55),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _2287_ (.RESET_B(net42),
    .D(_0012_),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _2288_ (.RESET_B(net41),
    .D(_0013_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _2289_ (.RESET_B(net40),
    .D(_0014_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _2290_ (.RESET_B(net39),
    .D(_0015_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _2291_ (.RESET_B(net38),
    .D(_0016_),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _2292_ (.RESET_B(net37),
    .D(_0017_),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _2293_ (.RESET_B(net46),
    .D(net51),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _2294_ (.RESET_B(net36),
    .D(net58),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _2295_ (.RESET_B(net35),
    .D(_0019_),
    .Q(\hvsync_gen.hpos[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _2296_ (.RESET_B(net34),
    .D(_0020_),
    .Q(\hvsync_gen.hpos[1] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _2297_ (.RESET_B(net33),
    .D(_0021_),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _2298_ (.RESET_B(net32),
    .D(_0022_),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _2299_ (.RESET_B(net31),
    .D(_0023_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _2300_ (.RESET_B(net30),
    .D(_0024_),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _2301_ (.RESET_B(net28),
    .D(_0025_),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _2302_ (.RESET_B(net27),
    .D(_0026_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _2303_ (.RESET_B(net26),
    .D(_0027_),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _2304_ (.RESET_B(net25),
    .D(_0028_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _2305_ (.RESET_B(net455),
    .D(_0029_),
    .Q(\dog_pos_x[0] ),
    .CLK(net427));
 sg13g2_dfrbpq_1 _2306_ (.RESET_B(net454),
    .D(_0030_),
    .Q(\dog_pos_x[1] ),
    .CLK(net426));
 sg13g2_dfrbpq_1 _2307_ (.RESET_B(net454),
    .D(_0031_),
    .Q(\dog_pos_x[2] ),
    .CLK(net426));
 sg13g2_dfrbpq_1 _2308_ (.RESET_B(net454),
    .D(_0032_),
    .Q(\dog_pos_x[3] ),
    .CLK(net426));
 sg13g2_dfrbpq_1 _2309_ (.RESET_B(net455),
    .D(_0033_),
    .Q(\dog_pos_x[4] ),
    .CLK(net427));
 sg13g2_dfrbpq_2 _2310_ (.RESET_B(net455),
    .D(_0034_),
    .Q(\dog_pos_x[5] ),
    .CLK(net427));
 sg13g2_dfrbpq_2 _2311_ (.RESET_B(net455),
    .D(_0035_),
    .Q(\dog_pos_x[6] ),
    .CLK(net427));
 sg13g2_dfrbpq_2 _2312_ (.RESET_B(net456),
    .D(_0036_),
    .Q(\dog_pos_x[7] ),
    .CLK(net428));
 sg13g2_dfrbpq_2 _2313_ (.RESET_B(net457),
    .D(_0037_),
    .Q(\dog_pos_x[8] ),
    .CLK(net428));
 sg13g2_dfrbpq_2 _2314_ (.RESET_B(net456),
    .D(_0038_),
    .Q(\dog_pos_x[9] ),
    .CLK(net428));
 sg13g2_dfrbpq_1 _2315_ (.RESET_B(net460),
    .D(_0039_),
    .Q(\dog_pos_y[0] ),
    .CLK(net433));
 sg13g2_dfrbpq_1 _2316_ (.RESET_B(net460),
    .D(_0040_),
    .Q(\dog_pos_y[1] ),
    .CLK(net431));
 sg13g2_dfrbpq_1 _2317_ (.RESET_B(net460),
    .D(_0041_),
    .Q(\dog_pos_y[2] ),
    .CLK(net431));
 sg13g2_dfrbpq_1 _2318_ (.RESET_B(net461),
    .D(_0042_),
    .Q(\dog_pos_y[3] ),
    .CLK(net431));
 sg13g2_dfrbpq_2 _2319_ (.RESET_B(net462),
    .D(_0043_),
    .Q(\dog_pos_y[4] ),
    .CLK(net432));
 sg13g2_dfrbpq_1 _2320_ (.RESET_B(net462),
    .D(_0044_),
    .Q(\dog_pos_y[5] ),
    .CLK(net432));
 sg13g2_dfrbpq_1 _2321_ (.RESET_B(net462),
    .D(_0045_),
    .Q(\dog_pos_y[6] ),
    .CLK(net431));
 sg13g2_dfrbpq_1 _2322_ (.RESET_B(net460),
    .D(_0046_),
    .Q(\dog_pos_y[7] ),
    .CLK(net431));
 sg13g2_dfrbpq_2 _2323_ (.RESET_B(net458),
    .D(_0047_),
    .Q(\dog_pos_y[8] ),
    .CLK(net429));
 sg13g2_dfrbpq_2 _2324_ (.RESET_B(net458),
    .D(_0048_),
    .Q(\dog_pos_y[9] ),
    .CLK(net429));
 sg13g2_dfrbpq_2 _2325_ (.RESET_B(net454),
    .D(_0049_),
    .Q(\square_x_pos[0] ),
    .CLK(net426));
 sg13g2_dfrbpq_2 _2326_ (.RESET_B(net456),
    .D(_0050_),
    .Q(\square_x_pos[1] ),
    .CLK(net428));
 sg13g2_dfrbpq_2 _2327_ (.RESET_B(net459),
    .D(_0051_),
    .Q(\square_x_pos[2] ),
    .CLK(net430));
 sg13g2_dfrbpq_1 _2328_ (.RESET_B(net459),
    .D(_0052_),
    .Q(\square_x_pos[3] ),
    .CLK(net430));
 sg13g2_dfrbpq_2 _2329_ (.RESET_B(net458),
    .D(_0053_),
    .Q(\square_x_pos[4] ),
    .CLK(net429));
 sg13g2_dfrbpq_2 _2330_ (.RESET_B(net459),
    .D(_0054_),
    .Q(\square_x_pos[5] ),
    .CLK(net430));
 sg13g2_dfrbpq_2 _2331_ (.RESET_B(net458),
    .D(_0055_),
    .Q(\square_x_pos[6] ),
    .CLK(net429));
 sg13g2_dfrbpq_2 _2332_ (.RESET_B(net458),
    .D(_0056_),
    .Q(\square_x_pos[7] ),
    .CLK(net429));
 sg13g2_dfrbpq_1 _2333_ (.RESET_B(net458),
    .D(_0057_),
    .Q(\square_x_pos[8] ),
    .CLK(net429));
 sg13g2_dfrbpq_1 _2334_ (.RESET_B(net456),
    .D(_0058_),
    .Q(\square_x_pos[9] ),
    .CLK(net428));
 sg13g2_dfrbpq_1 _2335_ (.RESET_B(net461),
    .D(_0059_),
    .Q(\square_y_pos[0] ),
    .CLK(net432));
 sg13g2_dfrbpq_2 _2336_ (.RESET_B(net461),
    .D(_0060_),
    .Q(\square_y_pos[1] ),
    .CLK(net432));
 sg13g2_dfrbpq_2 _2337_ (.RESET_B(net461),
    .D(_0061_),
    .Q(\square_y_pos[2] ),
    .CLK(net432));
 sg13g2_dfrbpq_2 _2338_ (.RESET_B(net461),
    .D(_0062_),
    .Q(\square_y_pos[3] ),
    .CLK(net432));
 sg13g2_dfrbpq_2 _2339_ (.RESET_B(net459),
    .D(_0063_),
    .Q(\square_y_pos[4] ),
    .CLK(net429));
 sg13g2_dfrbpq_2 _2340_ (.RESET_B(net458),
    .D(_0064_),
    .Q(\square_y_pos[5] ),
    .CLK(net429));
 sg13g2_dfrbpq_2 _2341_ (.RESET_B(net458),
    .D(_0065_),
    .Q(\square_y_pos[6] ),
    .CLK(net430));
 sg13g2_dfrbpq_2 _2342_ (.RESET_B(net460),
    .D(_0066_),
    .Q(\square_y_pos[7] ),
    .CLK(net432));
 sg13g2_dfrbpq_2 _2343_ (.RESET_B(net460),
    .D(_0067_),
    .Q(\square_y_pos[8] ),
    .CLK(net431));
 sg13g2_dfrbpq_1 _2344_ (.RESET_B(net460),
    .D(_0068_),
    .Q(\square_y_pos[9] ),
    .CLK(net431));
 sg13g2_dfrbpq_1 _2345_ (.RESET_B(net456),
    .D(_0069_),
    .Q(horz_dir),
    .CLK(net428));
 sg13g2_dfrbpq_2 _2346_ (.RESET_B(net454),
    .D(_0000_),
    .Q(\tick_count[0] ),
    .CLK(net426));
 sg13g2_dfrbpq_2 _2347_ (.RESET_B(net454),
    .D(_0001_),
    .Q(\tick_count[1] ),
    .CLK(net426));
 sg13g2_dfrbpq_1 _2348_ (.RESET_B(net454),
    .D(_0002_),
    .Q(\tick_count[2] ),
    .CLK(net426));
 sg13g2_dfrbpq_1 _2349_ (.RESET_B(net454),
    .D(_0003_),
    .Q(\tick_count[3] ),
    .CLK(net426));
 sg13g2_dfrbpq_1 _2350_ (.RESET_B(net460),
    .D(_0070_),
    .Q(vert_dir),
    .CLK(net431));
 sg13g2_tiehi _2303__26 (.L_HI(net26));
 sg13g2_tiehi _2302__27 (.L_HI(net27));
 sg13g2_tiehi _2301__28 (.L_HI(net28));
 sg13g2_tiehi _2280__29 (.L_HI(net29));
 sg13g2_tiehi _2300__30 (.L_HI(net30));
 sg13g2_tiehi _2299__31 (.L_HI(net31));
 sg13g2_tiehi _2298__32 (.L_HI(net32));
 sg13g2_tiehi _2297__33 (.L_HI(net33));
 sg13g2_tiehi _2296__34 (.L_HI(net34));
 sg13g2_tiehi _2295__35 (.L_HI(net35));
 sg13g2_tiehi _2294__36 (.L_HI(net36));
 sg13g2_tiehi _2292__37 (.L_HI(net37));
 sg13g2_tiehi _2291__38 (.L_HI(net38));
 sg13g2_tiehi _2290__39 (.L_HI(net39));
 sg13g2_tiehi _2289__40 (.L_HI(net40));
 sg13g2_tiehi _2288__41 (.L_HI(net41));
 sg13g2_tiehi _2287__42 (.L_HI(net42));
 sg13g2_tiehi _2286__43 (.L_HI(net43));
 sg13g2_tiehi _2285__44 (.L_HI(net44));
 sg13g2_tiehi _2284__45 (.L_HI(net45));
 sg13g2_tiehi _2293__46 (.L_HI(net46));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_vga_example_10 (.L_LO(net10));
 sg13g2_tielo tt_um_vga_example_11 (.L_LO(net11));
 sg13g2_tielo tt_um_vga_example_12 (.L_LO(net12));
 sg13g2_tielo tt_um_vga_example_13 (.L_LO(net13));
 sg13g2_tielo tt_um_vga_example_14 (.L_LO(net14));
 sg13g2_tielo tt_um_vga_example_15 (.L_LO(net15));
 sg13g2_tielo tt_um_vga_example_16 (.L_LO(net16));
 sg13g2_tielo tt_um_vga_example_17 (.L_LO(net17));
 sg13g2_tielo tt_um_vga_example_18 (.L_LO(net18));
 sg13g2_tielo tt_um_vga_example_19 (.L_LO(net19));
 sg13g2_tielo tt_um_vga_example_20 (.L_LO(net20));
 sg13g2_tielo tt_um_vga_example_21 (.L_LO(net21));
 sg13g2_tielo tt_um_vga_example_22 (.L_LO(net22));
 sg13g2_tielo tt_um_vga_example_23 (.L_LO(net23));
 sg13g2_tielo tt_um_vga_example_24 (.L_LO(net24));
 sg13g2_tiehi _2304__25 (.L_HI(net25));
 sg13g2_buf_1 _2389_ (.A(net430),
    .X(uo_out[3]));
 sg13g2_buf_1 _2390_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout315 (.A(net317),
    .X(net315));
 sg13g2_buf_1 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_8 fanout317 (.A(_0196_),
    .X(net317));
 sg13g2_buf_8 fanout318 (.A(_0196_),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(_0196_),
    .X(net319));
 sg13g2_buf_8 fanout320 (.A(net322),
    .X(net320));
 sg13g2_buf_1 fanout321 (.A(net322),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(_0093_),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(net324),
    .X(net323));
 sg13g2_buf_8 fanout324 (.A(_0093_),
    .X(net324));
 sg13g2_buf_8 fanout325 (.A(_1059_),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(_1056_),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(_0119_),
    .X(net327));
 sg13g2_buf_8 fanout328 (.A(_0346_),
    .X(net328));
 sg13g2_buf_8 fanout329 (.A(_0342_),
    .X(net329));
 sg13g2_buf_8 fanout330 (.A(_0335_),
    .X(net330));
 sg13g2_buf_8 fanout331 (.A(_0335_),
    .X(net331));
 sg13g2_buf_8 fanout332 (.A(_0333_),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(_0333_),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(_0332_),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(_0331_),
    .X(net335));
 sg13g2_buf_8 fanout336 (.A(_0331_),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_8 fanout338 (.A(_0330_),
    .X(net338));
 sg13g2_buf_1 fanout339 (.A(_0330_),
    .X(net339));
 sg13g2_buf_8 fanout340 (.A(_0322_),
    .X(net340));
 sg13g2_buf_8 fanout341 (.A(_0321_),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(_0320_),
    .X(net342));
 sg13g2_buf_8 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_8 fanout344 (.A(vert_dir),
    .X(net344));
 sg13g2_buf_8 fanout345 (.A(horz_dir),
    .X(net345));
 sg13g2_buf_1 fanout346 (.A(horz_dir),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(\dog_pos_y[8] ),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(\dog_pos_y[8] ),
    .X(net348));
 sg13g2_buf_8 fanout349 (.A(net350),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_8 fanout351 (.A(\dog_pos_y[7] ),
    .X(net351));
 sg13g2_buf_8 fanout352 (.A(\dog_pos_y[6] ),
    .X(net352));
 sg13g2_buf_8 fanout353 (.A(\dog_pos_y[5] ),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(\dog_pos_y[5] ),
    .X(net354));
 sg13g2_buf_8 fanout355 (.A(\dog_pos_y[4] ),
    .X(net355));
 sg13g2_buf_8 fanout356 (.A(\dog_pos_y[4] ),
    .X(net356));
 sg13g2_buf_8 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_8 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_8 fanout359 (.A(\dog_pos_y[3] ),
    .X(net359));
 sg13g2_buf_8 fanout360 (.A(net362),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_8 fanout362 (.A(net363),
    .X(net362));
 sg13g2_buf_8 fanout363 (.A(\dog_pos_y[2] ),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net365),
    .X(net364));
 sg13g2_buf_8 fanout365 (.A(net366),
    .X(net365));
 sg13g2_buf_1 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(\dog_pos_y[1] ),
    .X(net367));
 sg13g2_buf_8 fanout368 (.A(net370),
    .X(net368));
 sg13g2_buf_1 fanout369 (.A(net370),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(\dog_pos_y[0] ),
    .X(net370));
 sg13g2_buf_8 fanout371 (.A(\dog_pos_x[8] ),
    .X(net371));
 sg13g2_buf_8 fanout372 (.A(\dog_pos_x[8] ),
    .X(net372));
 sg13g2_buf_8 fanout373 (.A(\dog_pos_x[7] ),
    .X(net373));
 sg13g2_buf_8 fanout374 (.A(\dog_pos_x[6] ),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(\dog_pos_x[6] ),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(\dog_pos_x[5] ),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(\dog_pos_x[5] ),
    .X(net378));
 sg13g2_buf_8 fanout379 (.A(net381),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(net381),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(\dog_pos_x[4] ),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(net385),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(net385),
    .X(net383));
 sg13g2_buf_8 fanout384 (.A(net385),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(\dog_pos_x[3] ),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(net387),
    .X(net386));
 sg13g2_buf_8 fanout387 (.A(net389),
    .X(net387));
 sg13g2_buf_8 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_8 fanout389 (.A(\dog_pos_x[2] ),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(net391),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(net394),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(net394),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(\dog_pos_x[1] ),
    .X(net394));
 sg13g2_buf_8 fanout395 (.A(net396),
    .X(net395));
 sg13g2_buf_1 fanout396 (.A(net397),
    .X(net396));
 sg13g2_buf_1 fanout397 (.A(\dog_pos_x[0] ),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(_0340_),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(_0339_),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(_0338_),
    .X(net400));
 sg13g2_buf_8 fanout401 (.A(_0337_),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(_0326_),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(_0324_),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(net406),
    .X(net404));
 sg13g2_buf_8 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_8 fanout406 (.A(net59),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(net409),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(net69),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net412),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(net412),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(net65),
    .X(net412));
 sg13g2_buf_8 fanout413 (.A(\hvsync_gen.hpos[6] ),
    .X(net413));
 sg13g2_buf_8 fanout414 (.A(net60),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(net417),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(\hvsync_gen.hpos[5] ),
    .X(net417));
 sg13g2_buf_8 fanout418 (.A(net419),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(\hvsync_gen.hpos[4] ),
    .X(net419));
 sg13g2_buf_8 fanout420 (.A(net421),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net67),
    .X(net421));
 sg13g2_buf_8 fanout422 (.A(net423),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(net64),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(net49),
    .X(net424));
 sg13g2_buf_1 fanout425 (.A(\hvsync_gen.hpos[1] ),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_8 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(\hvsync_gen.vsync ),
    .X(net428));
 sg13g2_buf_8 fanout429 (.A(net433),
    .X(net429));
 sg13g2_buf_1 fanout430 (.A(net433),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net432),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(net433),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(\hvsync_gen.vsync ),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(net437),
    .X(net434));
 sg13g2_buf_8 fanout435 (.A(net437),
    .X(net435));
 sg13g2_buf_1 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(net70),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(net439),
    .X(net438));
 sg13g2_buf_8 fanout439 (.A(net440),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(net52),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(net442),
    .X(net441));
 sg13g2_buf_8 fanout442 (.A(\hvsync_gen.vpos[6] ),
    .X(net442));
 sg13g2_buf_8 fanout443 (.A(net445),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net445),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(net68),
    .X(net445));
 sg13g2_buf_8 fanout446 (.A(net53),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(\hvsync_gen.vpos[4] ),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(\hvsync_gen.vpos[3] ),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(net56),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(net54),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(\hvsync_gen.vpos[2] ),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(net62),
    .X(net452));
 sg13g2_buf_8 fanout453 (.A(net5),
    .X(net453));
 sg13g2_buf_8 fanout454 (.A(net455),
    .X(net454));
 sg13g2_buf_8 fanout455 (.A(net456),
    .X(net455));
 sg13g2_buf_8 fanout456 (.A(net457),
    .X(net456));
 sg13g2_buf_8 fanout457 (.A(rst_n),
    .X(net457));
 sg13g2_buf_8 fanout458 (.A(net462),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(net462),
    .X(net459));
 sg13g2_buf_8 fanout460 (.A(net461),
    .X(net460));
 sg13g2_buf_8 fanout461 (.A(net462),
    .X(net461));
 sg13g2_buf_8 fanout462 (.A(rst_n),
    .X(net462));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_vga_example_9 (.L_LO(net9));
 sg13g2_buf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_2_2__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hvsync_gen.hpos[0] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold2 (.A(\hvsync_gen.vpos[0] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold3 (.A(\hvsync_gen.hpos[1] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.vpos[9] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0018_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold6 (.A(\hvsync_gen.vpos[7] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold7 (.A(\hvsync_gen.vpos[4] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold8 (.A(\hvsync_gen.vpos[2] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0011_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold10 (.A(\hvsync_gen.vpos[3] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold11 (.A(_1045_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0005_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hvsync_gen.hpos[9] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold14 (.A(\hvsync_gen.hpos[6] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold15 (.A(_1088_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold16 (.A(\hvsync_gen.vpos[1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0010_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold18 (.A(\hvsync_gen.hpos[2] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hvsync_gen.hpos[7] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0004_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hvsync_gen.hpos[3] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hvsync_gen.vpos[5] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.hpos[8] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.vpos[8] ),
    .X(net70));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_4 FILLER_2_70 ();
 sg13g2_fill_1 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_79 ();
 sg13g2_decap_8 FILLER_2_86 ();
 sg13g2_decap_8 FILLER_2_93 ();
 sg13g2_decap_8 FILLER_2_100 ();
 sg13g2_decap_8 FILLER_2_107 ();
 sg13g2_decap_8 FILLER_2_114 ();
 sg13g2_decap_8 FILLER_2_121 ();
 sg13g2_decap_8 FILLER_2_128 ();
 sg13g2_decap_8 FILLER_2_135 ();
 sg13g2_decap_8 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_156 ();
 sg13g2_decap_8 FILLER_2_163 ();
 sg13g2_decap_8 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_8 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_decap_8 FILLER_2_212 ();
 sg13g2_decap_8 FILLER_2_219 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_7 ();
 sg13g2_decap_4 FILLER_3_12 ();
 sg13g2_fill_2 FILLER_3_16 ();
 sg13g2_fill_1 FILLER_3_22 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_fill_2 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_fill_2 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_fill_2 FILLER_3_130 ();
 sg13g2_fill_1 FILLER_3_132 ();
 sg13g2_decap_8 FILLER_3_146 ();
 sg13g2_decap_4 FILLER_3_153 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_4 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_172 ();
 sg13g2_fill_2 FILLER_3_186 ();
 sg13g2_fill_1 FILLER_3_188 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_4 FILLER_3_403 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_61 ();
 sg13g2_fill_2 FILLER_4_68 ();
 sg13g2_fill_1 FILLER_4_70 ();
 sg13g2_decap_4 FILLER_4_84 ();
 sg13g2_fill_2 FILLER_4_88 ();
 sg13g2_fill_2 FILLER_4_145 ();
 sg13g2_fill_1 FILLER_4_147 ();
 sg13g2_decap_4 FILLER_4_179 ();
 sg13g2_fill_2 FILLER_4_183 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_8 FILLER_4_223 ();
 sg13g2_decap_8 FILLER_4_230 ();
 sg13g2_decap_8 FILLER_4_237 ();
 sg13g2_decap_8 FILLER_4_244 ();
 sg13g2_decap_8 FILLER_4_251 ();
 sg13g2_decap_8 FILLER_4_258 ();
 sg13g2_decap_8 FILLER_4_265 ();
 sg13g2_decap_8 FILLER_4_272 ();
 sg13g2_decap_8 FILLER_4_279 ();
 sg13g2_decap_8 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_293 ();
 sg13g2_decap_8 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_decap_8 FILLER_4_314 ();
 sg13g2_fill_1 FILLER_4_321 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_decap_8 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_386 ();
 sg13g2_decap_8 FILLER_4_393 ();
 sg13g2_decap_8 FILLER_4_400 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_4 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_9 ();
 sg13g2_decap_8 FILLER_5_16 ();
 sg13g2_decap_4 FILLER_5_23 ();
 sg13g2_decap_4 FILLER_5_31 ();
 sg13g2_fill_2 FILLER_5_39 ();
 sg13g2_fill_1 FILLER_5_41 ();
 sg13g2_fill_2 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_52 ();
 sg13g2_fill_2 FILLER_5_59 ();
 sg13g2_fill_1 FILLER_5_61 ();
 sg13g2_fill_2 FILLER_5_67 ();
 sg13g2_fill_1 FILLER_5_120 ();
 sg13g2_decap_4 FILLER_5_134 ();
 sg13g2_fill_1 FILLER_5_138 ();
 sg13g2_decap_4 FILLER_5_160 ();
 sg13g2_fill_1 FILLER_5_175 ();
 sg13g2_fill_2 FILLER_5_190 ();
 sg13g2_fill_1 FILLER_5_192 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_4 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_4 FILLER_5_306 ();
 sg13g2_fill_2 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_fill_1 FILLER_5_351 ();
 sg13g2_decap_4 FILLER_5_357 ();
 sg13g2_fill_1 FILLER_5_361 ();
 sg13g2_fill_2 FILLER_5_366 ();
 sg13g2_fill_1 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_fill_2 FILLER_6_57 ();
 sg13g2_fill_2 FILLER_6_72 ();
 sg13g2_fill_2 FILLER_6_79 ();
 sg13g2_fill_1 FILLER_6_81 ();
 sg13g2_fill_2 FILLER_6_100 ();
 sg13g2_fill_1 FILLER_6_102 ();
 sg13g2_decap_4 FILLER_6_143 ();
 sg13g2_fill_2 FILLER_6_147 ();
 sg13g2_fill_2 FILLER_6_158 ();
 sg13g2_fill_1 FILLER_6_160 ();
 sg13g2_fill_2 FILLER_6_212 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_fill_2 FILLER_6_280 ();
 sg13g2_fill_2 FILLER_6_331 ();
 sg13g2_fill_2 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_fill_1 FILLER_6_399 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_24 ();
 sg13g2_decap_8 FILLER_7_31 ();
 sg13g2_fill_1 FILLER_7_44 ();
 sg13g2_decap_4 FILLER_7_50 ();
 sg13g2_fill_1 FILLER_7_54 ();
 sg13g2_decap_4 FILLER_7_63 ();
 sg13g2_decap_4 FILLER_7_73 ();
 sg13g2_fill_2 FILLER_7_86 ();
 sg13g2_fill_2 FILLER_7_101 ();
 sg13g2_fill_1 FILLER_7_112 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_decap_4 FILLER_7_141 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_decap_4 FILLER_7_166 ();
 sg13g2_decap_4 FILLER_7_242 ();
 sg13g2_decap_8 FILLER_7_250 ();
 sg13g2_fill_1 FILLER_7_257 ();
 sg13g2_decap_8 FILLER_7_262 ();
 sg13g2_decap_4 FILLER_7_269 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_fill_2 FILLER_7_298 ();
 sg13g2_fill_1 FILLER_7_300 ();
 sg13g2_fill_2 FILLER_7_319 ();
 sg13g2_fill_1 FILLER_7_352 ();
 sg13g2_fill_1 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_392 ();
 sg13g2_fill_1 FILLER_7_394 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_24 ();
 sg13g2_fill_1 FILLER_8_31 ();
 sg13g2_decap_4 FILLER_8_72 ();
 sg13g2_fill_1 FILLER_8_76 ();
 sg13g2_fill_1 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_90 ();
 sg13g2_fill_1 FILLER_8_92 ();
 sg13g2_fill_1 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_118 ();
 sg13g2_decap_4 FILLER_8_129 ();
 sg13g2_fill_1 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_1 FILLER_8_147 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_decap_4 FILLER_8_158 ();
 sg13g2_fill_1 FILLER_8_162 ();
 sg13g2_decap_4 FILLER_8_167 ();
 sg13g2_fill_2 FILLER_8_171 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_4 FILLER_8_188 ();
 sg13g2_fill_2 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_202 ();
 sg13g2_fill_2 FILLER_8_216 ();
 sg13g2_fill_1 FILLER_8_218 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_fill_1 FILLER_8_293 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_fill_2 FILLER_8_311 ();
 sg13g2_fill_2 FILLER_8_334 ();
 sg13g2_fill_1 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_fill_1 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_24 ();
 sg13g2_decap_8 FILLER_9_31 ();
 sg13g2_fill_1 FILLER_9_38 ();
 sg13g2_decap_8 FILLER_9_54 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_fill_2 FILLER_9_124 ();
 sg13g2_fill_2 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_159 ();
 sg13g2_decap_4 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_206 ();
 sg13g2_fill_1 FILLER_9_208 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_fill_2 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_292 ();
 sg13g2_fill_1 FILLER_9_299 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_fill_1 FILLER_9_354 ();
 sg13g2_decap_4 FILLER_9_360 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_4 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_17 ();
 sg13g2_decap_8 FILLER_10_33 ();
 sg13g2_fill_1 FILLER_10_40 ();
 sg13g2_decap_4 FILLER_10_54 ();
 sg13g2_fill_1 FILLER_10_58 ();
 sg13g2_fill_2 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_73 ();
 sg13g2_decap_8 FILLER_10_80 ();
 sg13g2_fill_2 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_103 ();
 sg13g2_decap_8 FILLER_10_111 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_139 ();
 sg13g2_decap_8 FILLER_10_155 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_fill_1 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_fill_2 FILLER_10_217 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_decap_4 FILLER_10_248 ();
 sg13g2_fill_2 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_decap_4 FILLER_10_269 ();
 sg13g2_fill_2 FILLER_10_273 ();
 sg13g2_fill_2 FILLER_10_376 ();
 sg13g2_fill_1 FILLER_10_378 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_decap_4 FILLER_11_21 ();
 sg13g2_fill_1 FILLER_11_25 ();
 sg13g2_fill_1 FILLER_11_78 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_fill_1 FILLER_11_99 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_fill_1 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_129 ();
 sg13g2_fill_2 FILLER_11_151 ();
 sg13g2_fill_1 FILLER_11_157 ();
 sg13g2_decap_4 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_190 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_fill_1 FILLER_11_204 ();
 sg13g2_decap_4 FILLER_11_228 ();
 sg13g2_fill_2 FILLER_11_264 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_fill_2 FILLER_11_301 ();
 sg13g2_fill_1 FILLER_11_309 ();
 sg13g2_fill_2 FILLER_11_315 ();
 sg13g2_decap_4 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_4 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_fill_1 FILLER_11_366 ();
 sg13g2_fill_2 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_25 ();
 sg13g2_fill_1 FILLER_12_27 ();
 sg13g2_fill_2 FILLER_12_38 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_decap_8 FILLER_12_52 ();
 sg13g2_decap_4 FILLER_12_59 ();
 sg13g2_fill_1 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_76 ();
 sg13g2_fill_2 FILLER_12_87 ();
 sg13g2_fill_2 FILLER_12_94 ();
 sg13g2_fill_1 FILLER_12_96 ();
 sg13g2_fill_2 FILLER_12_102 ();
 sg13g2_fill_1 FILLER_12_104 ();
 sg13g2_decap_4 FILLER_12_121 ();
 sg13g2_fill_2 FILLER_12_130 ();
 sg13g2_fill_1 FILLER_12_132 ();
 sg13g2_fill_2 FILLER_12_138 ();
 sg13g2_fill_2 FILLER_12_158 ();
 sg13g2_decap_4 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_fill_2 FILLER_12_234 ();
 sg13g2_decap_8 FILLER_12_248 ();
 sg13g2_fill_1 FILLER_12_259 ();
 sg13g2_fill_1 FILLER_12_273 ();
 sg13g2_fill_2 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_fill_2 FILLER_12_364 ();
 sg13g2_fill_1 FILLER_12_366 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_fill_2 FILLER_12_379 ();
 sg13g2_fill_2 FILLER_12_389 ();
 sg13g2_fill_1 FILLER_12_391 ();
 sg13g2_decap_4 FILLER_12_396 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_22 ();
 sg13g2_fill_1 FILLER_13_31 ();
 sg13g2_fill_2 FILLER_13_52 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_fill_2 FILLER_13_78 ();
 sg13g2_fill_1 FILLER_13_80 ();
 sg13g2_fill_2 FILLER_13_89 ();
 sg13g2_fill_1 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_108 ();
 sg13g2_fill_2 FILLER_13_126 ();
 sg13g2_fill_1 FILLER_13_148 ();
 sg13g2_fill_2 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_176 ();
 sg13g2_decap_4 FILLER_13_192 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_decap_4 FILLER_13_221 ();
 sg13g2_fill_1 FILLER_13_255 ();
 sg13g2_fill_2 FILLER_13_268 ();
 sg13g2_fill_1 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_289 ();
 sg13g2_fill_1 FILLER_13_308 ();
 sg13g2_decap_4 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_324 ();
 sg13g2_fill_1 FILLER_13_338 ();
 sg13g2_fill_2 FILLER_13_343 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_fill_2 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_4 FILLER_14_20 ();
 sg13g2_decap_8 FILLER_14_34 ();
 sg13g2_fill_1 FILLER_14_41 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_55 ();
 sg13g2_fill_1 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_75 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_decap_8 FILLER_14_97 ();
 sg13g2_fill_2 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_fill_2 FILLER_14_131 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_fill_1 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_146 ();
 sg13g2_decap_4 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_4 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_8 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_205 ();
 sg13g2_fill_1 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_decap_4 FILLER_14_248 ();
 sg13g2_fill_1 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_fill_2 FILLER_14_270 ();
 sg13g2_fill_1 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_290 ();
 sg13g2_fill_1 FILLER_14_311 ();
 sg13g2_fill_2 FILLER_14_317 ();
 sg13g2_fill_2 FILLER_14_328 ();
 sg13g2_fill_2 FILLER_14_338 ();
 sg13g2_decap_4 FILLER_14_350 ();
 sg13g2_decap_4 FILLER_14_359 ();
 sg13g2_decap_8 FILLER_14_373 ();
 sg13g2_decap_4 FILLER_14_380 ();
 sg13g2_fill_1 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_4 ();
 sg13g2_fill_2 FILLER_15_41 ();
 sg13g2_fill_1 FILLER_15_43 ();
 sg13g2_decap_4 FILLER_15_82 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_98 ();
 sg13g2_fill_1 FILLER_15_105 ();
 sg13g2_fill_1 FILLER_15_112 ();
 sg13g2_decap_4 FILLER_15_121 ();
 sg13g2_fill_2 FILLER_15_144 ();
 sg13g2_fill_1 FILLER_15_146 ();
 sg13g2_decap_4 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_177 ();
 sg13g2_decap_8 FILLER_15_184 ();
 sg13g2_fill_2 FILLER_15_198 ();
 sg13g2_fill_1 FILLER_15_200 ();
 sg13g2_decap_4 FILLER_15_215 ();
 sg13g2_fill_2 FILLER_15_219 ();
 sg13g2_fill_1 FILLER_15_245 ();
 sg13g2_fill_2 FILLER_15_253 ();
 sg13g2_fill_2 FILLER_15_277 ();
 sg13g2_decap_4 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_4 FILLER_15_315 ();
 sg13g2_fill_1 FILLER_15_319 ();
 sg13g2_fill_2 FILLER_15_338 ();
 sg13g2_fill_2 FILLER_15_362 ();
 sg13g2_fill_1 FILLER_15_364 ();
 sg13g2_fill_2 FILLER_15_380 ();
 sg13g2_fill_1 FILLER_15_382 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_2 FILLER_16_33 ();
 sg13g2_fill_1 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_fill_2 FILLER_16_67 ();
 sg13g2_fill_1 FILLER_16_69 ();
 sg13g2_fill_2 FILLER_16_83 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_107 ();
 sg13g2_decap_4 FILLER_16_138 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_1 FILLER_16_155 ();
 sg13g2_fill_2 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_178 ();
 sg13g2_fill_1 FILLER_16_180 ();
 sg13g2_decap_4 FILLER_16_199 ();
 sg13g2_fill_1 FILLER_16_203 ();
 sg13g2_fill_2 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_211 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_251 ();
 sg13g2_decap_4 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_283 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_4 FILLER_16_296 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_341 ();
 sg13g2_decap_4 FILLER_16_347 ();
 sg13g2_fill_1 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_369 ();
 sg13g2_fill_1 FILLER_16_376 ();
 sg13g2_decap_4 FILLER_16_403 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_2 FILLER_17_83 ();
 sg13g2_fill_1 FILLER_17_85 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_110 ();
 sg13g2_fill_2 FILLER_17_125 ();
 sg13g2_fill_2 FILLER_17_140 ();
 sg13g2_decap_4 FILLER_17_155 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_fill_2 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_decap_4 FILLER_17_209 ();
 sg13g2_decap_8 FILLER_17_225 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_264 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_decap_4 FILLER_17_288 ();
 sg13g2_fill_2 FILLER_17_302 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_4 FILLER_17_330 ();
 sg13g2_fill_1 FILLER_17_344 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_decap_4 FILLER_17_373 ();
 sg13g2_fill_1 FILLER_17_377 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_19 ();
 sg13g2_decap_8 FILLER_18_26 ();
 sg13g2_decap_8 FILLER_18_33 ();
 sg13g2_fill_1 FILLER_18_40 ();
 sg13g2_decap_4 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_57 ();
 sg13g2_decap_8 FILLER_18_80 ();
 sg13g2_fill_2 FILLER_18_87 ();
 sg13g2_fill_1 FILLER_18_89 ();
 sg13g2_decap_4 FILLER_18_102 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_163 ();
 sg13g2_fill_2 FILLER_18_171 ();
 sg13g2_fill_1 FILLER_18_181 ();
 sg13g2_fill_2 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_fill_2 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_4 FILLER_18_237 ();
 sg13g2_fill_1 FILLER_18_241 ();
 sg13g2_fill_2 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_fill_2 FILLER_18_272 ();
 sg13g2_decap_4 FILLER_18_285 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_fill_1 FILLER_18_303 ();
 sg13g2_decap_4 FILLER_18_309 ();
 sg13g2_decap_4 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_321 ();
 sg13g2_fill_2 FILLER_18_328 ();
 sg13g2_fill_2 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_339 ();
 sg13g2_decap_4 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_decap_4 FILLER_18_377 ();
 sg13g2_fill_1 FILLER_18_381 ();
 sg13g2_decap_4 FILLER_18_404 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_20 ();
 sg13g2_decap_4 FILLER_19_34 ();
 sg13g2_decap_4 FILLER_19_58 ();
 sg13g2_fill_1 FILLER_19_62 ();
 sg13g2_fill_2 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_fill_2 FILLER_19_127 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_decap_4 FILLER_19_135 ();
 sg13g2_fill_2 FILLER_19_139 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_4 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_179 ();
 sg13g2_fill_1 FILLER_19_184 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_251 ();
 sg13g2_decap_4 FILLER_19_262 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_2 FILLER_19_293 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_fill_1 FILLER_19_303 ();
 sg13g2_fill_1 FILLER_19_340 ();
 sg13g2_fill_2 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_363 ();
 sg13g2_fill_2 FILLER_19_385 ();
 sg13g2_fill_1 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_31 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_54 ();
 sg13g2_decap_4 FILLER_20_87 ();
 sg13g2_fill_1 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_104 ();
 sg13g2_fill_2 FILLER_20_111 ();
 sg13g2_fill_2 FILLER_20_118 ();
 sg13g2_fill_1 FILLER_20_120 ();
 sg13g2_decap_4 FILLER_20_188 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_232 ();
 sg13g2_fill_1 FILLER_20_243 ();
 sg13g2_fill_1 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_258 ();
 sg13g2_fill_1 FILLER_20_260 ();
 sg13g2_decap_4 FILLER_20_269 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_fill_2 FILLER_20_343 ();
 sg13g2_fill_1 FILLER_20_345 ();
 sg13g2_fill_2 FILLER_20_355 ();
 sg13g2_fill_1 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_363 ();
 sg13g2_decap_4 FILLER_20_370 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_decap_4 FILLER_20_385 ();
 sg13g2_fill_1 FILLER_20_389 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_4 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_decap_4 FILLER_21_57 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_72 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_99 ();
 sg13g2_fill_1 FILLER_21_101 ();
 sg13g2_fill_2 FILLER_21_114 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_decap_4 FILLER_21_132 ();
 sg13g2_fill_1 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_157 ();
 sg13g2_fill_1 FILLER_21_159 ();
 sg13g2_decap_4 FILLER_21_164 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_fill_2 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_fill_2 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_decap_8 FILLER_21_317 ();
 sg13g2_decap_4 FILLER_21_324 ();
 sg13g2_decap_4 FILLER_21_346 ();
 sg13g2_fill_1 FILLER_21_391 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_41 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_decap_4 FILLER_22_73 ();
 sg13g2_decap_4 FILLER_22_90 ();
 sg13g2_fill_1 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_fill_2 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_135 ();
 sg13g2_decap_8 FILLER_22_170 ();
 sg13g2_fill_2 FILLER_22_177 ();
 sg13g2_fill_1 FILLER_22_179 ();
 sg13g2_fill_2 FILLER_22_188 ();
 sg13g2_fill_1 FILLER_22_190 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_decap_8 FILLER_22_223 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_fill_1 FILLER_22_232 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_268 ();
 sg13g2_fill_1 FILLER_22_270 ();
 sg13g2_decap_4 FILLER_22_284 ();
 sg13g2_decap_4 FILLER_22_292 ();
 sg13g2_decap_4 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_319 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_decap_4 FILLER_22_336 ();
 sg13g2_decap_4 FILLER_22_346 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_4 FILLER_22_377 ();
 sg13g2_fill_1 FILLER_22_385 ();
 sg13g2_fill_1 FILLER_22_394 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_20 ();
 sg13g2_decap_8 FILLER_23_34 ();
 sg13g2_fill_1 FILLER_23_41 ();
 sg13g2_decap_4 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_decap_4 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_fill_1 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_4 FILLER_23_165 ();
 sg13g2_decap_4 FILLER_23_179 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_198 ();
 sg13g2_decap_4 FILLER_23_205 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_fill_2 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_fill_2 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_261 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_277 ();
 sg13g2_fill_2 FILLER_23_285 ();
 sg13g2_fill_2 FILLER_23_300 ();
 sg13g2_fill_1 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_fill_2 FILLER_23_346 ();
 sg13g2_decap_4 FILLER_23_365 ();
 sg13g2_fill_2 FILLER_23_369 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_fill_2 FILLER_24_30 ();
 sg13g2_fill_1 FILLER_24_32 ();
 sg13g2_fill_2 FILLER_24_45 ();
 sg13g2_fill_1 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_56 ();
 sg13g2_fill_1 FILLER_24_58 ();
 sg13g2_fill_2 FILLER_24_67 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_decap_4 FILLER_24_75 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_fill_2 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_110 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_fill_1 FILLER_24_141 ();
 sg13g2_decap_4 FILLER_24_159 ();
 sg13g2_fill_1 FILLER_24_163 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_210 ();
 sg13g2_decap_4 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_257 ();
 sg13g2_fill_2 FILLER_24_308 ();
 sg13g2_fill_1 FILLER_24_310 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_334 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_fill_1 FILLER_24_342 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_fill_2 FILLER_25_32 ();
 sg13g2_decap_4 FILLER_25_71 ();
 sg13g2_fill_2 FILLER_25_108 ();
 sg13g2_decap_8 FILLER_25_136 ();
 sg13g2_decap_8 FILLER_25_143 ();
 sg13g2_decap_4 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_decap_4 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_242 ();
 sg13g2_fill_1 FILLER_25_249 ();
 sg13g2_decap_4 FILLER_25_262 ();
 sg13g2_decap_8 FILLER_25_271 ();
 sg13g2_decap_4 FILLER_25_278 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_decap_4 FILLER_25_294 ();
 sg13g2_fill_2 FILLER_25_305 ();
 sg13g2_fill_2 FILLER_25_318 ();
 sg13g2_fill_1 FILLER_25_336 ();
 sg13g2_decap_4 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_4 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_47 ();
 sg13g2_fill_2 FILLER_26_54 ();
 sg13g2_fill_1 FILLER_26_56 ();
 sg13g2_fill_1 FILLER_26_62 ();
 sg13g2_decap_8 FILLER_26_68 ();
 sg13g2_fill_2 FILLER_26_75 ();
 sg13g2_fill_1 FILLER_26_77 ();
 sg13g2_fill_2 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_decap_8 FILLER_26_212 ();
 sg13g2_decap_4 FILLER_26_219 ();
 sg13g2_fill_2 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_254 ();
 sg13g2_fill_2 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_decap_4 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_4 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_4 FILLER_26_309 ();
 sg13g2_fill_1 FILLER_26_313 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_fill_2 FILLER_26_392 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_27 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_1 FILLER_27_71 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_fill_2 FILLER_27_98 ();
 sg13g2_fill_2 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_118 ();
 sg13g2_decap_8 FILLER_27_127 ();
 sg13g2_decap_4 FILLER_27_138 ();
 sg13g2_fill_1 FILLER_27_142 ();
 sg13g2_decap_4 FILLER_27_147 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_decap_8 FILLER_27_160 ();
 sg13g2_decap_8 FILLER_27_194 ();
 sg13g2_decap_4 FILLER_27_201 ();
 sg13g2_decap_4 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_245 ();
 sg13g2_decap_4 FILLER_27_263 ();
 sg13g2_decap_4 FILLER_27_290 ();
 sg13g2_fill_2 FILLER_27_294 ();
 sg13g2_decap_4 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_325 ();
 sg13g2_fill_2 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_341 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_2 ();
 sg13g2_fill_2 FILLER_28_29 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_4 FILLER_28_56 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_187 ();
 sg13g2_decap_8 FILLER_28_194 ();
 sg13g2_decap_8 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_fill_2 FILLER_28_237 ();
 sg13g2_fill_1 FILLER_28_239 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_305 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_317 ();
 sg13g2_decap_4 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_2 FILLER_28_375 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_4 FILLER_29_27 ();
 sg13g2_fill_1 FILLER_29_31 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_4 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_73 ();
 sg13g2_fill_1 FILLER_29_75 ();
 sg13g2_decap_8 FILLER_29_83 ();
 sg13g2_decap_4 FILLER_29_90 ();
 sg13g2_fill_1 FILLER_29_94 ();
 sg13g2_decap_4 FILLER_29_108 ();
 sg13g2_decap_4 FILLER_29_122 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_fill_2 FILLER_29_147 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_1 FILLER_29_171 ();
 sg13g2_fill_2 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_decap_8 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_decap_4 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_267 ();
 sg13g2_fill_2 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_343 ();
 sg13g2_fill_1 FILLER_29_345 ();
 sg13g2_decap_4 FILLER_29_363 ();
 sg13g2_fill_1 FILLER_29_367 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_384 ();
 sg13g2_decap_4 FILLER_29_391 ();
 sg13g2_fill_1 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_4 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_11 ();
 sg13g2_decap_8 FILLER_30_55 ();
 sg13g2_fill_2 FILLER_30_62 ();
 sg13g2_decap_8 FILLER_30_71 ();
 sg13g2_decap_4 FILLER_30_78 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_fill_2 FILLER_30_92 ();
 sg13g2_fill_1 FILLER_30_94 ();
 sg13g2_decap_4 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_124 ();
 sg13g2_fill_1 FILLER_30_150 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_177 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_decap_4 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_decap_8 FILLER_30_239 ();
 sg13g2_decap_4 FILLER_30_246 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_fill_1 FILLER_30_358 ();
 sg13g2_fill_2 FILLER_30_367 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_decap_4 FILLER_30_403 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_40 ();
 sg13g2_fill_2 FILLER_31_47 ();
 sg13g2_fill_1 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_58 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_decap_4 FILLER_31_99 ();
 sg13g2_decap_8 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_121 ();
 sg13g2_fill_1 FILLER_31_123 ();
 sg13g2_decap_4 FILLER_31_129 ();
 sg13g2_fill_2 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_31_143 ();
 sg13g2_fill_1 FILLER_31_145 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_decap_8 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_decap_8 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_292 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_decap_4 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_335 ();
 sg13g2_decap_4 FILLER_31_342 ();
 sg13g2_fill_1 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_370 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_4 FILLER_32_27 ();
 sg13g2_fill_2 FILLER_32_72 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_fill_2 FILLER_32_128 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_fill_2 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_177 ();
 sg13g2_fill_2 FILLER_32_188 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_fill_2 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_32_201 ();
 sg13g2_fill_2 FILLER_32_230 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_288 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_299 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_fill_2 FILLER_32_376 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_29 ();
 sg13g2_decap_4 FILLER_33_36 ();
 sg13g2_fill_2 FILLER_33_40 ();
 sg13g2_fill_2 FILLER_33_55 ();
 sg13g2_fill_1 FILLER_33_86 ();
 sg13g2_fill_2 FILLER_33_94 ();
 sg13g2_decap_4 FILLER_33_107 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_fill_2 FILLER_33_134 ();
 sg13g2_decap_4 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_decap_4 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_358 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_11 ();
 sg13g2_fill_1 FILLER_34_18 ();
 sg13g2_fill_2 FILLER_34_55 ();
 sg13g2_fill_1 FILLER_34_57 ();
 sg13g2_decap_8 FILLER_34_80 ();
 sg13g2_decap_4 FILLER_34_106 ();
 sg13g2_fill_2 FILLER_34_110 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_163 ();
 sg13g2_decap_8 FILLER_34_168 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_fill_2 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_decap_4 FILLER_34_204 ();
 sg13g2_fill_2 FILLER_34_212 ();
 sg13g2_decap_4 FILLER_34_227 ();
 sg13g2_fill_1 FILLER_34_231 ();
 sg13g2_decap_8 FILLER_34_248 ();
 sg13g2_decap_8 FILLER_34_255 ();
 sg13g2_decap_8 FILLER_34_262 ();
 sg13g2_decap_4 FILLER_34_269 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_decap_4 FILLER_34_286 ();
 sg13g2_fill_1 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_294 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_308 ();
 sg13g2_fill_2 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_323 ();
 sg13g2_fill_1 FILLER_34_342 ();
 sg13g2_decap_4 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_fill_2 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_fill_2 FILLER_34_385 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_36 ();
 sg13g2_decap_8 FILLER_35_43 ();
 sg13g2_fill_1 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_64 ();
 sg13g2_fill_2 FILLER_35_93 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_decap_4 FILLER_35_139 ();
 sg13g2_fill_1 FILLER_35_143 ();
 sg13g2_decap_4 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_fill_2 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_4 FILLER_35_315 ();
 sg13g2_fill_2 FILLER_35_319 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_decap_4 FILLER_35_367 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_36_62 ();
 sg13g2_decap_8 FILLER_36_69 ();
 sg13g2_fill_2 FILLER_36_76 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_110 ();
 sg13g2_decap_8 FILLER_36_117 ();
 sg13g2_fill_2 FILLER_36_124 ();
 sg13g2_fill_1 FILLER_36_126 ();
 sg13g2_fill_2 FILLER_36_141 ();
 sg13g2_decap_8 FILLER_36_148 ();
 sg13g2_decap_4 FILLER_36_155 ();
 sg13g2_fill_2 FILLER_36_159 ();
 sg13g2_decap_8 FILLER_36_170 ();
 sg13g2_decap_4 FILLER_36_177 ();
 sg13g2_fill_2 FILLER_36_181 ();
 sg13g2_decap_4 FILLER_36_188 ();
 sg13g2_fill_1 FILLER_36_192 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_decap_8 FILLER_36_220 ();
 sg13g2_fill_2 FILLER_36_240 ();
 sg13g2_decap_4 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_321 ();
 sg13g2_fill_1 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_335 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_1 FILLER_37_18 ();
 sg13g2_decap_8 FILLER_37_29 ();
 sg13g2_decap_8 FILLER_37_36 ();
 sg13g2_decap_8 FILLER_37_43 ();
 sg13g2_decap_8 FILLER_37_50 ();
 sg13g2_decap_4 FILLER_37_57 ();
 sg13g2_fill_1 FILLER_37_61 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_331 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_370 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_139 ();
 sg13g2_fill_1 FILLER_38_141 ();
 sg13g2_fill_2 FILLER_38_150 ();
 sg13g2_fill_2 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_209 ();
 sg13g2_decap_8 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_223 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_240 ();
 sg13g2_decap_8 FILLER_38_248 ();
 sg13g2_decap_8 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_262 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_325 ();
 sg13g2_fill_1 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_333 ();
 sg13g2_fill_1 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_359 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
