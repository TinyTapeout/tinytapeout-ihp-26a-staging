module tt_um_techhu_rv32_trial (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire clk_regs;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire \addr[0] ;
 wire \addr[10] ;
 wire \addr[11] ;
 wire \addr[12] ;
 wire \addr[13] ;
 wire \addr[14] ;
 wire \addr[15] ;
 wire \addr[16] ;
 wire \addr[17] ;
 wire \addr[18] ;
 wire \addr[19] ;
 wire \addr[1] ;
 wire \addr[20] ;
 wire \addr[21] ;
 wire \addr[22] ;
 wire \addr[23] ;
 wire \addr[24] ;
 wire \addr[25] ;
 wire \addr[26] ;
 wire \addr[27] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire combined_rst_n;
 wire \crc16_read[0] ;
 wire \crc16_read[10] ;
 wire \crc16_read[11] ;
 wire \crc16_read[12] ;
 wire \crc16_read[13] ;
 wire \crc16_read[14] ;
 wire \crc16_read[15] ;
 wire \crc16_read[1] ;
 wire \crc16_read[2] ;
 wire \crc16_read[3] ;
 wire \crc16_read[4] ;
 wire \crc16_read[5] ;
 wire \crc16_read[6] ;
 wire \crc16_read[7] ;
 wire \crc16_read[8] ;
 wire \crc16_read[9] ;
 wire \crc_peri_data[0] ;
 wire \crc_peri_data[1] ;
 wire \crc_peri_data[2] ;
 wire \crc_peri_data[3] ;
 wire \crc_peri_data[4] ;
 wire \crc_peri_data[5] ;
 wire \crc_peri_data[6] ;
 wire \crc_peri_data[7] ;
 wire \data_to_write[10] ;
 wire \data_to_write[11] ;
 wire \data_to_write[12] ;
 wire \data_to_write[13] ;
 wire \data_to_write[14] ;
 wire \data_to_write[15] ;
 wire \data_to_write[16] ;
 wire \data_to_write[17] ;
 wire \data_to_write[18] ;
 wire \data_to_write[19] ;
 wire \data_to_write[20] ;
 wire \data_to_write[21] ;
 wire \data_to_write[22] ;
 wire \data_to_write[23] ;
 wire \data_to_write[24] ;
 wire \data_to_write[25] ;
 wire \data_to_write[26] ;
 wire \data_to_write[27] ;
 wire \data_to_write[28] ;
 wire \data_to_write[29] ;
 wire \data_to_write[30] ;
 wire \data_to_write[31] ;
 wire \data_to_write[8] ;
 wire \data_to_write[9] ;
 wire debug_data_continue;
 wire debug_instr_valid;
 wire \dio1_sync[0] ;
 wire \dio1_sync[1] ;
 wire \gpio_out[0] ;
 wire \gpio_out[1] ;
 wire \gpio_out[2] ;
 wire \gpio_out[3] ;
 wire \gpio_out[4] ;
 wire \gpio_out[5] ;
 wire \gpio_out[6] ;
 wire \gpio_out[7] ;
 wire \gpio_out_sel[0] ;
 wire \gpio_out_sel[1] ;
 wire \gpio_out_sel[2] ;
 wire \gpio_out_sel[3] ;
 wire \gpio_out_sel[4] ;
 wire \gpio_out_sel[5] ;
 wire \gpio_out_sel[6] ;
 wire \gpio_out_sel[7] ;
 wire \i2c_config_out[0] ;
 wire \i2c_config_out[10] ;
 wire \i2c_config_out[11] ;
 wire \i2c_config_out[12] ;
 wire \i2c_config_out[13] ;
 wire \i2c_config_out[14] ;
 wire \i2c_config_out[15] ;
 wire \i2c_config_out[1] ;
 wire \i2c_config_out[2] ;
 wire \i2c_config_out[3] ;
 wire \i2c_config_out[4] ;
 wire \i2c_config_out[5] ;
 wire \i2c_config_out[6] ;
 wire \i2c_config_out[7] ;
 wire \i2c_config_out[8] ;
 wire \i2c_config_out[9] ;
 wire \i2c_data_out[0] ;
 wire \i2c_data_out[1] ;
 wire \i2c_data_out[2] ;
 wire \i2c_data_out[3] ;
 wire \i2c_data_out[4] ;
 wire \i2c_data_out[5] ;
 wire \i2c_data_out[6] ;
 wire \i2c_data_out[7] ;
 wire \i2c_data_out[8] ;
 wire \i_crc16.bit_cnt[0] ;
 wire \i_crc16.bit_cnt[1] ;
 wire \i_crc16.bit_cnt[2] ;
 wire \i_crc16.bit_cnt[3] ;
 wire \i_crc16.rst_n ;
 wire \i_i2c_peri.addr_latch[0] ;
 wire \i_i2c_peri.addr_latch[1] ;
 wire \i_i2c_peri.addr_latch[2] ;
 wire \i_i2c_peri.addr_latch[3] ;
 wire \i_i2c_peri.addr_latch[4] ;
 wire \i_i2c_peri.addr_latch[5] ;
 wire \i_i2c_peri.addr_latch[6] ;
 wire \i_i2c_peri.cmd_addr_reg[0] ;
 wire \i_i2c_peri.cmd_addr_reg[1] ;
 wire \i_i2c_peri.cmd_addr_reg[2] ;
 wire \i_i2c_peri.cmd_addr_reg[3] ;
 wire \i_i2c_peri.cmd_addr_reg[4] ;
 wire \i_i2c_peri.cmd_addr_reg[5] ;
 wire \i_i2c_peri.cmd_addr_reg[6] ;
 wire \i_i2c_peri.cmd_pending ;
 wire \i_i2c_peri.cmd_read_reg ;
 wire \i_i2c_peri.cmd_start_reg ;
 wire \i_i2c_peri.cmd_stop_reg ;
 wire \i_i2c_peri.cmd_write_m_reg ;
 wire \i_i2c_peri.i_i2c.addr_reg[0] ;
 wire \i_i2c_peri.i_i2c.addr_reg[1] ;
 wire \i_i2c_peri.i_i2c.addr_reg[2] ;
 wire \i_i2c_peri.i_i2c.addr_reg[3] ;
 wire \i_i2c_peri.i_i2c.addr_reg[4] ;
 wire \i_i2c_peri.i_i2c.addr_reg[5] ;
 wire \i_i2c_peri.i_i2c.addr_reg[6] ;
 wire \i_i2c_peri.i_i2c.bit_count_reg[0] ;
 wire \i_i2c_peri.i_i2c.bit_count_reg[1] ;
 wire \i_i2c_peri.i_i2c.bit_count_reg[2] ;
 wire \i_i2c_peri.i_i2c.bit_count_reg[3] ;
 wire \i_i2c_peri.i_i2c.bus_active_reg ;
 wire \i_i2c_peri.i_i2c.busy_reg ;
 wire \i_i2c_peri.i_i2c.data_reg[0] ;
 wire \i_i2c_peri.i_i2c.data_reg[1] ;
 wire \i_i2c_peri.i_i2c.data_reg[2] ;
 wire \i_i2c_peri.i_i2c.data_reg[3] ;
 wire \i_i2c_peri.i_i2c.data_reg[4] ;
 wire \i_i2c_peri.i_i2c.data_reg[5] ;
 wire \i_i2c_peri.i_i2c.data_reg[6] ;
 wire \i_i2c_peri.i_i2c.data_reg[7] ;
 wire \i_i2c_peri.i_i2c.delay_reg[0] ;
 wire \i_i2c_peri.i_i2c.delay_reg[10] ;
 wire \i_i2c_peri.i_i2c.delay_reg[11] ;
 wire \i_i2c_peri.i_i2c.delay_reg[12] ;
 wire \i_i2c_peri.i_i2c.delay_reg[13] ;
 wire \i_i2c_peri.i_i2c.delay_reg[14] ;
 wire \i_i2c_peri.i_i2c.delay_reg[15] ;
 wire \i_i2c_peri.i_i2c.delay_reg[16] ;
 wire \i_i2c_peri.i_i2c.delay_reg[1] ;
 wire \i_i2c_peri.i_i2c.delay_reg[2] ;
 wire \i_i2c_peri.i_i2c.delay_reg[3] ;
 wire \i_i2c_peri.i_i2c.delay_reg[4] ;
 wire \i_i2c_peri.i_i2c.delay_reg[5] ;
 wire \i_i2c_peri.i_i2c.delay_reg[6] ;
 wire \i_i2c_peri.i_i2c.delay_reg[7] ;
 wire \i_i2c_peri.i_i2c.delay_reg[8] ;
 wire \i_i2c_peri.i_i2c.delay_reg[9] ;
 wire \i_i2c_peri.i_i2c.delay_scl_reg ;
 wire \i_i2c_peri.i_i2c.delay_sda_reg ;
 wire \i_i2c_peri.i_i2c.last_reg ;
 wire \i_i2c_peri.i_i2c.last_sda_i_reg ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[0] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[1] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[2] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[3] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[4] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[5] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[6] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tdata_reg[7] ;
 wire \i_i2c_peri.i_i2c.m_axis_data_tvalid_reg ;
 wire \i_i2c_peri.i_i2c.missed_ack_reg ;
 wire \i_i2c_peri.i_i2c.mode_read_reg ;
 wire \i_i2c_peri.i_i2c.mode_stop_reg ;
 wire \i_i2c_peri.i_i2c.mode_write_multiple_reg ;
 wire \i_i2c_peri.i_i2c.phy_rx_data_reg ;
 wire \i_i2c_peri.i_i2c.phy_state_reg[0] ;
 wire \i_i2c_peri.i_i2c.phy_state_reg[1] ;
 wire \i_i2c_peri.i_i2c.phy_state_reg[2] ;
 wire \i_i2c_peri.i_i2c.phy_state_reg[3] ;
 wire \i_i2c_peri.i_i2c.s_axis_cmd_ready_reg ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[0] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[1] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[2] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[3] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[4] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[5] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[6] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tdata[7] ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tlast ;
 wire \i_i2c_peri.i_i2c.s_axis_data_tready_reg ;
 wire \i_i2c_peri.i_i2c.scl_o_reg ;
 wire \i_i2c_peri.i_i2c.sda_i ;
 wire \i_i2c_peri.i_i2c.sda_i_reg ;
 wire \i_i2c_peri.i_i2c.sda_o_reg ;
 wire \i_i2c_peri.i_i2c.state_reg[0] ;
 wire \i_i2c_peri.i_i2c.state_reg[1] ;
 wire \i_i2c_peri.i_i2c.state_reg[2] ;
 wire \i_i2c_peri.i_i2c.state_reg[3] ;
 wire \i_i2c_peri.rx_has_data ;
 wire \i_i2c_peri.sda_sync[0] ;
 wire \i_i2c_peri.tx_pending ;
 wire \i_latch_mem.cycle[0] ;
 wire \i_latch_mem.cycle[1] ;
 wire \i_latch_mem.data_out[0] ;
 wire \i_latch_mem.data_out[10] ;
 wire \i_latch_mem.data_out[11] ;
 wire \i_latch_mem.data_out[12] ;
 wire \i_latch_mem.data_out[13] ;
 wire \i_latch_mem.data_out[14] ;
 wire \i_latch_mem.data_out[15] ;
 wire \i_latch_mem.data_out[16] ;
 wire \i_latch_mem.data_out[17] ;
 wire \i_latch_mem.data_out[18] ;
 wire \i_latch_mem.data_out[19] ;
 wire \i_latch_mem.data_out[1] ;
 wire \i_latch_mem.data_out[20] ;
 wire \i_latch_mem.data_out[21] ;
 wire \i_latch_mem.data_out[22] ;
 wire \i_latch_mem.data_out[23] ;
 wire \i_latch_mem.data_out[24] ;
 wire \i_latch_mem.data_out[25] ;
 wire \i_latch_mem.data_out[26] ;
 wire \i_latch_mem.data_out[27] ;
 wire \i_latch_mem.data_out[28] ;
 wire \i_latch_mem.data_out[29] ;
 wire \i_latch_mem.data_out[2] ;
 wire \i_latch_mem.data_out[30] ;
 wire \i_latch_mem.data_out[31] ;
 wire \i_latch_mem.data_out[3] ;
 wire \i_latch_mem.data_out[4] ;
 wire \i_latch_mem.data_out[5] ;
 wire \i_latch_mem.data_out[6] ;
 wire \i_latch_mem.data_out[7] ;
 wire \i_latch_mem.data_out[8] ;
 wire \i_latch_mem.data_out[9] ;
 wire \i_latch_mem.data_ready ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[0].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[10].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[11].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[12].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[13].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[14].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[15].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[16].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[17].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[18].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[19].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[1].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[20].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[21].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[22].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[23].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[24].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[25].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[26].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[27].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[28].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[29].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[2].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[30].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[31].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[3].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[4].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[5].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[6].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[7].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[8].l_ram.data_out[7] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[0] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[1] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[2] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[3] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[4] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[5] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[6] ;
 wire \i_latch_mem.genblk1[9].l_ram.data_out[7] ;
 wire \i_rtc.seconds_out[0] ;
 wire \i_rtc.seconds_out[10] ;
 wire \i_rtc.seconds_out[11] ;
 wire \i_rtc.seconds_out[12] ;
 wire \i_rtc.seconds_out[13] ;
 wire \i_rtc.seconds_out[14] ;
 wire \i_rtc.seconds_out[15] ;
 wire \i_rtc.seconds_out[16] ;
 wire \i_rtc.seconds_out[17] ;
 wire \i_rtc.seconds_out[18] ;
 wire \i_rtc.seconds_out[19] ;
 wire \i_rtc.seconds_out[1] ;
 wire \i_rtc.seconds_out[20] ;
 wire \i_rtc.seconds_out[21] ;
 wire \i_rtc.seconds_out[22] ;
 wire \i_rtc.seconds_out[23] ;
 wire \i_rtc.seconds_out[24] ;
 wire \i_rtc.seconds_out[25] ;
 wire \i_rtc.seconds_out[26] ;
 wire \i_rtc.seconds_out[27] ;
 wire \i_rtc.seconds_out[28] ;
 wire \i_rtc.seconds_out[29] ;
 wire \i_rtc.seconds_out[2] ;
 wire \i_rtc.seconds_out[30] ;
 wire \i_rtc.seconds_out[31] ;
 wire \i_rtc.seconds_out[3] ;
 wire \i_rtc.seconds_out[4] ;
 wire \i_rtc.seconds_out[5] ;
 wire \i_rtc.seconds_out[6] ;
 wire \i_rtc.seconds_out[7] ;
 wire \i_rtc.seconds_out[8] ;
 wire \i_rtc.seconds_out[9] ;
 wire \i_rtc.us_count[0] ;
 wire \i_rtc.us_count[10] ;
 wire \i_rtc.us_count[11] ;
 wire \i_rtc.us_count[12] ;
 wire \i_rtc.us_count[13] ;
 wire \i_rtc.us_count[14] ;
 wire \i_rtc.us_count[15] ;
 wire \i_rtc.us_count[16] ;
 wire \i_rtc.us_count[17] ;
 wire \i_rtc.us_count[18] ;
 wire \i_rtc.us_count[19] ;
 wire \i_rtc.us_count[1] ;
 wire \i_rtc.us_count[2] ;
 wire \i_rtc.us_count[3] ;
 wire \i_rtc.us_count[4] ;
 wire \i_rtc.us_count[5] ;
 wire \i_rtc.us_count[6] ;
 wire \i_rtc.us_count[7] ;
 wire \i_rtc.us_count[8] ;
 wire \i_rtc.us_count[9] ;
 wire \i_seal.byte_idx[0] ;
 wire \i_seal.byte_idx[1] ;
 wire \i_seal.byte_idx[2] ;
 wire \i_seal.byte_idx[3] ;
 wire \i_seal.byte_sent ;
 wire \i_seal.commit_dropped ;
 wire \i_seal.crc_byte[0] ;
 wire \i_seal.crc_byte[1] ;
 wire \i_seal.crc_byte[2] ;
 wire \i_seal.crc_byte[3] ;
 wire \i_seal.crc_byte[4] ;
 wire \i_seal.crc_byte[5] ;
 wire \i_seal.crc_byte[6] ;
 wire \i_seal.crc_byte[7] ;
 wire \i_seal.crc_feed ;
 wire \i_seal.crc_init ;
 wire \i_seal.cur_mono[0] ;
 wire \i_seal.cur_mono[10] ;
 wire \i_seal.cur_mono[11] ;
 wire \i_seal.cur_mono[12] ;
 wire \i_seal.cur_mono[13] ;
 wire \i_seal.cur_mono[14] ;
 wire \i_seal.cur_mono[15] ;
 wire \i_seal.cur_mono[16] ;
 wire \i_seal.cur_mono[17] ;
 wire \i_seal.cur_mono[18] ;
 wire \i_seal.cur_mono[19] ;
 wire \i_seal.cur_mono[1] ;
 wire \i_seal.cur_mono[20] ;
 wire \i_seal.cur_mono[21] ;
 wire \i_seal.cur_mono[22] ;
 wire \i_seal.cur_mono[23] ;
 wire \i_seal.cur_mono[24] ;
 wire \i_seal.cur_mono[25] ;
 wire \i_seal.cur_mono[26] ;
 wire \i_seal.cur_mono[27] ;
 wire \i_seal.cur_mono[28] ;
 wire \i_seal.cur_mono[29] ;
 wire \i_seal.cur_mono[2] ;
 wire \i_seal.cur_mono[30] ;
 wire \i_seal.cur_mono[31] ;
 wire \i_seal.cur_mono[3] ;
 wire \i_seal.cur_mono[4] ;
 wire \i_seal.cur_mono[5] ;
 wire \i_seal.cur_mono[6] ;
 wire \i_seal.cur_mono[7] ;
 wire \i_seal.cur_mono[8] ;
 wire \i_seal.cur_mono[9] ;
 wire \i_seal.mono_count[0] ;
 wire \i_seal.mono_count[10] ;
 wire \i_seal.mono_count[11] ;
 wire \i_seal.mono_count[12] ;
 wire \i_seal.mono_count[13] ;
 wire \i_seal.mono_count[14] ;
 wire \i_seal.mono_count[15] ;
 wire \i_seal.mono_count[16] ;
 wire \i_seal.mono_count[17] ;
 wire \i_seal.mono_count[18] ;
 wire \i_seal.mono_count[19] ;
 wire \i_seal.mono_count[1] ;
 wire \i_seal.mono_count[20] ;
 wire \i_seal.mono_count[21] ;
 wire \i_seal.mono_count[22] ;
 wire \i_seal.mono_count[23] ;
 wire \i_seal.mono_count[24] ;
 wire \i_seal.mono_count[25] ;
 wire \i_seal.mono_count[26] ;
 wire \i_seal.mono_count[27] ;
 wire \i_seal.mono_count[28] ;
 wire \i_seal.mono_count[29] ;
 wire \i_seal.mono_count[2] ;
 wire \i_seal.mono_count[30] ;
 wire \i_seal.mono_count[31] ;
 wire \i_seal.mono_count[3] ;
 wire \i_seal.mono_count[4] ;
 wire \i_seal.mono_count[5] ;
 wire \i_seal.mono_count[6] ;
 wire \i_seal.mono_count[7] ;
 wire \i_seal.mono_count[8] ;
 wire \i_seal.mono_count[9] ;
 wire \i_seal.read_seq[0] ;
 wire \i_seal.read_seq[1] ;
 wire \i_seal.sealed_crc[0] ;
 wire \i_seal.sealed_crc[10] ;
 wire \i_seal.sealed_crc[11] ;
 wire \i_seal.sealed_crc[12] ;
 wire \i_seal.sealed_crc[13] ;
 wire \i_seal.sealed_crc[14] ;
 wire \i_seal.sealed_crc[15] ;
 wire \i_seal.sealed_crc[1] ;
 wire \i_seal.sealed_crc[2] ;
 wire \i_seal.sealed_crc[3] ;
 wire \i_seal.sealed_crc[4] ;
 wire \i_seal.sealed_crc[5] ;
 wire \i_seal.sealed_crc[6] ;
 wire \i_seal.sealed_crc[7] ;
 wire \i_seal.sealed_crc[8] ;
 wire \i_seal.sealed_crc[9] ;
 wire \i_seal.sealed_mono[0] ;
 wire \i_seal.sealed_mono[10] ;
 wire \i_seal.sealed_mono[11] ;
 wire \i_seal.sealed_mono[12] ;
 wire \i_seal.sealed_mono[13] ;
 wire \i_seal.sealed_mono[14] ;
 wire \i_seal.sealed_mono[15] ;
 wire \i_seal.sealed_mono[16] ;
 wire \i_seal.sealed_mono[17] ;
 wire \i_seal.sealed_mono[18] ;
 wire \i_seal.sealed_mono[19] ;
 wire \i_seal.sealed_mono[1] ;
 wire \i_seal.sealed_mono[20] ;
 wire \i_seal.sealed_mono[21] ;
 wire \i_seal.sealed_mono[22] ;
 wire \i_seal.sealed_mono[23] ;
 wire \i_seal.sealed_mono[24] ;
 wire \i_seal.sealed_mono[25] ;
 wire \i_seal.sealed_mono[26] ;
 wire \i_seal.sealed_mono[27] ;
 wire \i_seal.sealed_mono[28] ;
 wire \i_seal.sealed_mono[29] ;
 wire \i_seal.sealed_mono[2] ;
 wire \i_seal.sealed_mono[30] ;
 wire \i_seal.sealed_mono[31] ;
 wire \i_seal.sealed_mono[3] ;
 wire \i_seal.sealed_mono[4] ;
 wire \i_seal.sealed_mono[5] ;
 wire \i_seal.sealed_mono[6] ;
 wire \i_seal.sealed_mono[7] ;
 wire \i_seal.sealed_mono[8] ;
 wire \i_seal.sealed_mono[9] ;
 wire \i_seal.sealed_sid[0] ;
 wire \i_seal.sealed_sid[1] ;
 wire \i_seal.sealed_sid[2] ;
 wire \i_seal.sealed_sid[3] ;
 wire \i_seal.sealed_sid[4] ;
 wire \i_seal.sealed_sid[5] ;
 wire \i_seal.sealed_sid[6] ;
 wire \i_seal.sealed_sid[7] ;
 wire \i_seal.sealed_value[0] ;
 wire \i_seal.sealed_value[10] ;
 wire \i_seal.sealed_value[11] ;
 wire \i_seal.sealed_value[12] ;
 wire \i_seal.sealed_value[13] ;
 wire \i_seal.sealed_value[14] ;
 wire \i_seal.sealed_value[15] ;
 wire \i_seal.sealed_value[16] ;
 wire \i_seal.sealed_value[17] ;
 wire \i_seal.sealed_value[18] ;
 wire \i_seal.sealed_value[19] ;
 wire \i_seal.sealed_value[1] ;
 wire \i_seal.sealed_value[20] ;
 wire \i_seal.sealed_value[21] ;
 wire \i_seal.sealed_value[22] ;
 wire \i_seal.sealed_value[23] ;
 wire \i_seal.sealed_value[24] ;
 wire \i_seal.sealed_value[25] ;
 wire \i_seal.sealed_value[26] ;
 wire \i_seal.sealed_value[27] ;
 wire \i_seal.sealed_value[28] ;
 wire \i_seal.sealed_value[29] ;
 wire \i_seal.sealed_value[2] ;
 wire \i_seal.sealed_value[30] ;
 wire \i_seal.sealed_value[31] ;
 wire \i_seal.sealed_value[3] ;
 wire \i_seal.sealed_value[4] ;
 wire \i_seal.sealed_value[5] ;
 wire \i_seal.sealed_value[6] ;
 wire \i_seal.sealed_value[7] ;
 wire \i_seal.sealed_value[8] ;
 wire \i_seal.sealed_value[9] ;
 wire \i_seal.sensor_id_reg[0] ;
 wire \i_seal.sensor_id_reg[1] ;
 wire \i_seal.sensor_id_reg[2] ;
 wire \i_seal.sensor_id_reg[3] ;
 wire \i_seal.sensor_id_reg[4] ;
 wire \i_seal.sensor_id_reg[5] ;
 wire \i_seal.sensor_id_reg[6] ;
 wire \i_seal.sensor_id_reg[7] ;
 wire \i_seal.session_ctr_in[0] ;
 wire \i_seal.session_ctr_in[1] ;
 wire \i_seal.session_ctr_in[2] ;
 wire \i_seal.session_ctr_in[3] ;
 wire \i_seal.session_ctr_in[4] ;
 wire \i_seal.session_ctr_in[5] ;
 wire \i_seal.session_ctr_in[6] ;
 wire \i_seal.session_ctr_in[7] ;
 wire \i_seal.session_locked ;
 wire \i_seal.state[0] ;
 wire \i_seal.state[1] ;
 wire \i_seal.value_reg[0] ;
 wire \i_seal.value_reg[10] ;
 wire \i_seal.value_reg[11] ;
 wire \i_seal.value_reg[12] ;
 wire \i_seal.value_reg[13] ;
 wire \i_seal.value_reg[14] ;
 wire \i_seal.value_reg[15] ;
 wire \i_seal.value_reg[16] ;
 wire \i_seal.value_reg[17] ;
 wire \i_seal.value_reg[18] ;
 wire \i_seal.value_reg[19] ;
 wire \i_seal.value_reg[1] ;
 wire \i_seal.value_reg[20] ;
 wire \i_seal.value_reg[21] ;
 wire \i_seal.value_reg[22] ;
 wire \i_seal.value_reg[23] ;
 wire \i_seal.value_reg[24] ;
 wire \i_seal.value_reg[25] ;
 wire \i_seal.value_reg[26] ;
 wire \i_seal.value_reg[27] ;
 wire \i_seal.value_reg[28] ;
 wire \i_seal.value_reg[29] ;
 wire \i_seal.value_reg[2] ;
 wire \i_seal.value_reg[30] ;
 wire \i_seal.value_reg[31] ;
 wire \i_seal.value_reg[3] ;
 wire \i_seal.value_reg[4] ;
 wire \i_seal.value_reg[5] ;
 wire \i_seal.value_reg[6] ;
 wire \i_seal.value_reg[7] ;
 wire \i_seal.value_reg[8] ;
 wire \i_seal.value_reg[9] ;
 wire \i_spi.bits_remaining[0] ;
 wire \i_spi.bits_remaining[1] ;
 wire \i_spi.bits_remaining[2] ;
 wire \i_spi.bits_remaining[3] ;
 wire \i_spi.busy ;
 wire \i_spi.clock_count[0] ;
 wire \i_spi.clock_count[1] ;
 wire \i_spi.clock_count[2] ;
 wire \i_spi.clock_count[3] ;
 wire \i_spi.clock_divider[0] ;
 wire \i_spi.clock_divider[1] ;
 wire \i_spi.clock_divider[2] ;
 wire \i_spi.clock_divider[3] ;
 wire \i_spi.data[0] ;
 wire \i_spi.data[1] ;
 wire \i_spi.data[2] ;
 wire \i_spi.data[3] ;
 wire \i_spi.data[4] ;
 wire \i_spi.data[5] ;
 wire \i_spi.data[6] ;
 wire \i_spi.data[7] ;
 wire \i_spi.end_txn_reg ;
 wire \i_spi.read_latency ;
 wire \i_spi.spi_clk_out ;
 wire \i_spi.spi_select ;
 wire \i_tinyqv.cpu.additional_mem_ops[0] ;
 wire \i_tinyqv.cpu.additional_mem_ops[1] ;
 wire \i_tinyqv.cpu.additional_mem_ops[2] ;
 wire \i_tinyqv.cpu.alu_op[0] ;
 wire \i_tinyqv.cpu.alu_op[1] ;
 wire \i_tinyqv.cpu.alu_op[2] ;
 wire \i_tinyqv.cpu.alu_op[3] ;
 wire \i_tinyqv.cpu.counter[2] ;
 wire \i_tinyqv.cpu.counter[3] ;
 wire \i_tinyqv.cpu.counter[4] ;
 wire \i_tinyqv.cpu.data_read_n[0] ;
 wire \i_tinyqv.cpu.data_read_n[1] ;
 wire \i_tinyqv.cpu.data_ready_latch ;
 wire \i_tinyqv.cpu.data_ready_sync ;
 wire \i_tinyqv.cpu.data_write_n[0] ;
 wire \i_tinyqv.cpu.data_write_n[1] ;
 wire \i_tinyqv.cpu.i_core.cmp ;
 wire \i_tinyqv.cpu.i_core.cmp_out ;
 wire \i_tinyqv.cpu.i_core.cy ;
 wire \i_tinyqv.cpu.i_core.cy_out ;
 wire \i_tinyqv.cpu.i_core.cycle[0] ;
 wire \i_tinyqv.cpu.i_core.cycle[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[0] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[2] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[3] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[4] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[5] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[6] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.cy ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.rstn ;
 wire \i_tinyqv.cpu.i_core.i_instrret.add ;
 wire \i_tinyqv.cpu.i_core.i_instrret.cy ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[0] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[1] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[2] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[3] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[10] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[11] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[12] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[13] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[14] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[15] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[16] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[17] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[18] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[19] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[20] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[21] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[22] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[23] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[24] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[25] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[26] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[27] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[28] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[29] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[30] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[31] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[4] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[5] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[6] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[7] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[8] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[9] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[0] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[10] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[11] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[1] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[2] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[3] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[5] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[6] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[7] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[8] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[9] ;
 wire \i_tinyqv.cpu.i_core.is_double_fault_r ;
 wire \i_tinyqv.cpu.i_core.is_interrupt ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.load_done ;
 wire \i_tinyqv.cpu.i_core.load_top_bit ;
 wire \i_tinyqv.cpu.i_core.mcause[0] ;
 wire \i_tinyqv.cpu.i_core.mcause[1] ;
 wire \i_tinyqv.cpu.i_core.mcause[3] ;
 wire \i_tinyqv.cpu.i_core.mcause[4] ;
 wire \i_tinyqv.cpu.i_core.mem_op[0] ;
 wire \i_tinyqv.cpu.i_core.mem_op[1] ;
 wire \i_tinyqv.cpu.i_core.mem_op[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[0] ;
 wire \i_tinyqv.cpu.i_core.mepc[10] ;
 wire \i_tinyqv.cpu.i_core.mepc[11] ;
 wire \i_tinyqv.cpu.i_core.mepc[12] ;
 wire \i_tinyqv.cpu.i_core.mepc[13] ;
 wire \i_tinyqv.cpu.i_core.mepc[14] ;
 wire \i_tinyqv.cpu.i_core.mepc[15] ;
 wire \i_tinyqv.cpu.i_core.mepc[16] ;
 wire \i_tinyqv.cpu.i_core.mepc[17] ;
 wire \i_tinyqv.cpu.i_core.mepc[18] ;
 wire \i_tinyqv.cpu.i_core.mepc[19] ;
 wire \i_tinyqv.cpu.i_core.mepc[1] ;
 wire \i_tinyqv.cpu.i_core.mepc[20] ;
 wire \i_tinyqv.cpu.i_core.mepc[21] ;
 wire \i_tinyqv.cpu.i_core.mepc[22] ;
 wire \i_tinyqv.cpu.i_core.mepc[23] ;
 wire \i_tinyqv.cpu.i_core.mepc[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[3] ;
 wire \i_tinyqv.cpu.i_core.mepc[4] ;
 wire \i_tinyqv.cpu.i_core.mepc[5] ;
 wire \i_tinyqv.cpu.i_core.mepc[6] ;
 wire \i_tinyqv.cpu.i_core.mepc[7] ;
 wire \i_tinyqv.cpu.i_core.mepc[8] ;
 wire \i_tinyqv.cpu.i_core.mepc[9] ;
 wire \i_tinyqv.cpu.i_core.mie[0] ;
 wire \i_tinyqv.cpu.i_core.mie[1] ;
 wire \i_tinyqv.cpu.i_core.mie[2] ;
 wire \i_tinyqv.cpu.i_core.mie[3] ;
 wire \i_tinyqv.cpu.i_core.mie[4] ;
 wire \i_tinyqv.cpu.i_core.mip[0] ;
 wire \i_tinyqv.cpu.i_core.mip[1] ;
 wire \i_tinyqv.cpu.i_core.mstatus_mie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mpie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mte ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[0] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[10] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[11] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[12] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[13] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[14] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[15] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[1] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[2] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[3] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[4] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[5] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[6] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[7] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[8] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[9] ;
 wire \i_tinyqv.cpu.i_core.time_hi[0] ;
 wire \i_tinyqv.cpu.i_core.time_hi[1] ;
 wire \i_tinyqv.cpu.i_core.time_hi[2] ;
 wire \i_tinyqv.cpu.imm[12] ;
 wire \i_tinyqv.cpu.imm[13] ;
 wire \i_tinyqv.cpu.imm[14] ;
 wire \i_tinyqv.cpu.imm[15] ;
 wire \i_tinyqv.cpu.imm[16] ;
 wire \i_tinyqv.cpu.imm[17] ;
 wire \i_tinyqv.cpu.imm[18] ;
 wire \i_tinyqv.cpu.imm[19] ;
 wire \i_tinyqv.cpu.imm[20] ;
 wire \i_tinyqv.cpu.imm[21] ;
 wire \i_tinyqv.cpu.imm[22] ;
 wire \i_tinyqv.cpu.imm[23] ;
 wire \i_tinyqv.cpu.imm[24] ;
 wire \i_tinyqv.cpu.imm[25] ;
 wire \i_tinyqv.cpu.imm[26] ;
 wire \i_tinyqv.cpu.imm[27] ;
 wire \i_tinyqv.cpu.imm[28] ;
 wire \i_tinyqv.cpu.imm[29] ;
 wire \i_tinyqv.cpu.imm[30] ;
 wire \i_tinyqv.cpu.imm[31] ;
 wire \i_tinyqv.cpu.instr_data[0][0] ;
 wire \i_tinyqv.cpu.instr_data[0][10] ;
 wire \i_tinyqv.cpu.instr_data[0][11] ;
 wire \i_tinyqv.cpu.instr_data[0][12] ;
 wire \i_tinyqv.cpu.instr_data[0][13] ;
 wire \i_tinyqv.cpu.instr_data[0][14] ;
 wire \i_tinyqv.cpu.instr_data[0][15] ;
 wire \i_tinyqv.cpu.instr_data[0][1] ;
 wire \i_tinyqv.cpu.instr_data[0][2] ;
 wire \i_tinyqv.cpu.instr_data[0][3] ;
 wire \i_tinyqv.cpu.instr_data[0][4] ;
 wire \i_tinyqv.cpu.instr_data[0][5] ;
 wire \i_tinyqv.cpu.instr_data[0][6] ;
 wire \i_tinyqv.cpu.instr_data[0][7] ;
 wire \i_tinyqv.cpu.instr_data[0][8] ;
 wire \i_tinyqv.cpu.instr_data[0][9] ;
 wire \i_tinyqv.cpu.instr_data[1][0] ;
 wire \i_tinyqv.cpu.instr_data[1][10] ;
 wire \i_tinyqv.cpu.instr_data[1][11] ;
 wire \i_tinyqv.cpu.instr_data[1][12] ;
 wire \i_tinyqv.cpu.instr_data[1][13] ;
 wire \i_tinyqv.cpu.instr_data[1][14] ;
 wire \i_tinyqv.cpu.instr_data[1][15] ;
 wire \i_tinyqv.cpu.instr_data[1][1] ;
 wire \i_tinyqv.cpu.instr_data[1][2] ;
 wire \i_tinyqv.cpu.instr_data[1][3] ;
 wire \i_tinyqv.cpu.instr_data[1][4] ;
 wire \i_tinyqv.cpu.instr_data[1][5] ;
 wire \i_tinyqv.cpu.instr_data[1][6] ;
 wire \i_tinyqv.cpu.instr_data[1][7] ;
 wire \i_tinyqv.cpu.instr_data[1][8] ;
 wire \i_tinyqv.cpu.instr_data[1][9] ;
 wire \i_tinyqv.cpu.instr_data[2][0] ;
 wire \i_tinyqv.cpu.instr_data[2][10] ;
 wire \i_tinyqv.cpu.instr_data[2][11] ;
 wire \i_tinyqv.cpu.instr_data[2][12] ;
 wire \i_tinyqv.cpu.instr_data[2][13] ;
 wire \i_tinyqv.cpu.instr_data[2][14] ;
 wire \i_tinyqv.cpu.instr_data[2][15] ;
 wire \i_tinyqv.cpu.instr_data[2][1] ;
 wire \i_tinyqv.cpu.instr_data[2][2] ;
 wire \i_tinyqv.cpu.instr_data[2][3] ;
 wire \i_tinyqv.cpu.instr_data[2][4] ;
 wire \i_tinyqv.cpu.instr_data[2][5] ;
 wire \i_tinyqv.cpu.instr_data[2][6] ;
 wire \i_tinyqv.cpu.instr_data[2][7] ;
 wire \i_tinyqv.cpu.instr_data[2][8] ;
 wire \i_tinyqv.cpu.instr_data[2][9] ;
 wire \i_tinyqv.cpu.instr_data[3][0] ;
 wire \i_tinyqv.cpu.instr_data[3][10] ;
 wire \i_tinyqv.cpu.instr_data[3][11] ;
 wire \i_tinyqv.cpu.instr_data[3][12] ;
 wire \i_tinyqv.cpu.instr_data[3][13] ;
 wire \i_tinyqv.cpu.instr_data[3][14] ;
 wire \i_tinyqv.cpu.instr_data[3][15] ;
 wire \i_tinyqv.cpu.instr_data[3][1] ;
 wire \i_tinyqv.cpu.instr_data[3][2] ;
 wire \i_tinyqv.cpu.instr_data[3][3] ;
 wire \i_tinyqv.cpu.instr_data[3][4] ;
 wire \i_tinyqv.cpu.instr_data[3][5] ;
 wire \i_tinyqv.cpu.instr_data[3][6] ;
 wire \i_tinyqv.cpu.instr_data[3][7] ;
 wire \i_tinyqv.cpu.instr_data[3][8] ;
 wire \i_tinyqv.cpu.instr_data[3][9] ;
 wire \i_tinyqv.cpu.instr_data_in[0] ;
 wire \i_tinyqv.cpu.instr_data_in[10] ;
 wire \i_tinyqv.cpu.instr_data_in[11] ;
 wire \i_tinyqv.cpu.instr_data_in[12] ;
 wire \i_tinyqv.cpu.instr_data_in[13] ;
 wire \i_tinyqv.cpu.instr_data_in[14] ;
 wire \i_tinyqv.cpu.instr_data_in[15] ;
 wire \i_tinyqv.cpu.instr_data_in[1] ;
 wire \i_tinyqv.cpu.instr_data_in[2] ;
 wire \i_tinyqv.cpu.instr_data_in[3] ;
 wire \i_tinyqv.cpu.instr_data_in[4] ;
 wire \i_tinyqv.cpu.instr_data_in[5] ;
 wire \i_tinyqv.cpu.instr_data_in[6] ;
 wire \i_tinyqv.cpu.instr_data_in[7] ;
 wire \i_tinyqv.cpu.instr_data_in[8] ;
 wire \i_tinyqv.cpu.instr_data_in[9] ;
 wire \i_tinyqv.cpu.instr_data_start[10] ;
 wire \i_tinyqv.cpu.instr_data_start[11] ;
 wire \i_tinyqv.cpu.instr_data_start[12] ;
 wire \i_tinyqv.cpu.instr_data_start[13] ;
 wire \i_tinyqv.cpu.instr_data_start[14] ;
 wire \i_tinyqv.cpu.instr_data_start[15] ;
 wire \i_tinyqv.cpu.instr_data_start[16] ;
 wire \i_tinyqv.cpu.instr_data_start[17] ;
 wire \i_tinyqv.cpu.instr_data_start[18] ;
 wire \i_tinyqv.cpu.instr_data_start[19] ;
 wire \i_tinyqv.cpu.instr_data_start[20] ;
 wire \i_tinyqv.cpu.instr_data_start[21] ;
 wire \i_tinyqv.cpu.instr_data_start[22] ;
 wire \i_tinyqv.cpu.instr_data_start[23] ;
 wire \i_tinyqv.cpu.instr_data_start[3] ;
 wire \i_tinyqv.cpu.instr_data_start[4] ;
 wire \i_tinyqv.cpu.instr_data_start[5] ;
 wire \i_tinyqv.cpu.instr_data_start[6] ;
 wire \i_tinyqv.cpu.instr_data_start[7] ;
 wire \i_tinyqv.cpu.instr_data_start[8] ;
 wire \i_tinyqv.cpu.instr_data_start[9] ;
 wire \i_tinyqv.cpu.instr_fetch_running ;
 wire \i_tinyqv.cpu.instr_fetch_started ;
 wire \i_tinyqv.cpu.instr_fetch_stopped ;
 wire \i_tinyqv.cpu.instr_len[1] ;
 wire \i_tinyqv.cpu.instr_len[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[1] ;
 wire \i_tinyqv.cpu.instr_write_offset[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[3] ;
 wire \i_tinyqv.cpu.is_alu_imm ;
 wire \i_tinyqv.cpu.is_alu_reg ;
 wire \i_tinyqv.cpu.is_auipc ;
 wire \i_tinyqv.cpu.is_branch ;
 wire \i_tinyqv.cpu.is_jal ;
 wire \i_tinyqv.cpu.is_jalr ;
 wire \i_tinyqv.cpu.is_load ;
 wire \i_tinyqv.cpu.is_lui ;
 wire \i_tinyqv.cpu.is_store ;
 wire \i_tinyqv.cpu.is_system ;
 wire \i_tinyqv.cpu.load_started ;
 wire \i_tinyqv.cpu.mem_op_increment_reg ;
 wire \i_tinyqv.cpu.no_write_in_progress ;
 wire \i_tinyqv.cpu.pc[1] ;
 wire \i_tinyqv.cpu.pc[2] ;
 wire \i_tinyqv.cpu.was_early_branch ;
 wire \i_tinyqv.mem.data_from_read[16] ;
 wire \i_tinyqv.mem.data_from_read[17] ;
 wire \i_tinyqv.mem.data_from_read[18] ;
 wire \i_tinyqv.mem.data_from_read[19] ;
 wire \i_tinyqv.mem.data_from_read[20] ;
 wire \i_tinyqv.mem.data_from_read[21] ;
 wire \i_tinyqv.mem.data_from_read[22] ;
 wire \i_tinyqv.mem.data_from_read[23] ;
 wire \i_tinyqv.mem.data_stall ;
 wire \i_tinyqv.mem.instr_active ;
 wire \i_tinyqv.mem.q_ctrl.addr[0] ;
 wire \i_tinyqv.mem.q_ctrl.addr[10] ;
 wire \i_tinyqv.mem.q_ctrl.addr[11] ;
 wire \i_tinyqv.mem.q_ctrl.addr[12] ;
 wire \i_tinyqv.mem.q_ctrl.addr[13] ;
 wire \i_tinyqv.mem.q_ctrl.addr[14] ;
 wire \i_tinyqv.mem.q_ctrl.addr[15] ;
 wire \i_tinyqv.mem.q_ctrl.addr[16] ;
 wire \i_tinyqv.mem.q_ctrl.addr[17] ;
 wire \i_tinyqv.mem.q_ctrl.addr[18] ;
 wire \i_tinyqv.mem.q_ctrl.addr[19] ;
 wire \i_tinyqv.mem.q_ctrl.addr[1] ;
 wire \i_tinyqv.mem.q_ctrl.addr[20] ;
 wire \i_tinyqv.mem.q_ctrl.addr[21] ;
 wire \i_tinyqv.mem.q_ctrl.addr[22] ;
 wire \i_tinyqv.mem.q_ctrl.addr[23] ;
 wire \i_tinyqv.mem.q_ctrl.addr[2] ;
 wire \i_tinyqv.mem.q_ctrl.addr[3] ;
 wire \i_tinyqv.mem.q_ctrl.addr[4] ;
 wire \i_tinyqv.mem.q_ctrl.addr[5] ;
 wire \i_tinyqv.mem.q_ctrl.addr[6] ;
 wire \i_tinyqv.mem.q_ctrl.addr[7] ;
 wire \i_tinyqv.mem.q_ctrl.addr[8] ;
 wire \i_tinyqv.mem.q_ctrl.addr[9] ;
 wire \i_tinyqv.mem.q_ctrl.data_ready ;
 wire \i_tinyqv.mem.q_ctrl.data_req ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[0] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[2] ;
 wire \i_tinyqv.mem.q_ctrl.is_writing ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_a_sel ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_b_sel ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[0] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_neg ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_out ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_pos ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_use_neg ;
 wire \i_tinyqv.mem.q_ctrl.spi_data_oe[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_flash_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_a_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_b_select ;
 wire \i_tinyqv.mem.q_ctrl.stop_txn_reg ;
 wire \i_tinyqv.mem.qspi_data_buf[10] ;
 wire \i_tinyqv.mem.qspi_data_buf[11] ;
 wire \i_tinyqv.mem.qspi_data_buf[12] ;
 wire \i_tinyqv.mem.qspi_data_buf[13] ;
 wire \i_tinyqv.mem.qspi_data_buf[14] ;
 wire \i_tinyqv.mem.qspi_data_buf[15] ;
 wire \i_tinyqv.mem.qspi_data_buf[24] ;
 wire \i_tinyqv.mem.qspi_data_buf[25] ;
 wire \i_tinyqv.mem.qspi_data_buf[26] ;
 wire \i_tinyqv.mem.qspi_data_buf[27] ;
 wire \i_tinyqv.mem.qspi_data_buf[28] ;
 wire \i_tinyqv.mem.qspi_data_buf[29] ;
 wire \i_tinyqv.mem.qspi_data_buf[30] ;
 wire \i_tinyqv.mem.qspi_data_buf[31] ;
 wire \i_tinyqv.mem.qspi_data_buf[8] ;
 wire \i_tinyqv.mem.qspi_data_buf[9] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[0] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[1] ;
 wire \i_tinyqv.mem.qspi_write_done ;
 wire \i_uart_rx.bit_sample ;
 wire \i_uart_rx.cycle_counter[0] ;
 wire \i_uart_rx.cycle_counter[1] ;
 wire \i_uart_rx.cycle_counter[2] ;
 wire \i_uart_rx.cycle_counter[3] ;
 wire \i_uart_rx.cycle_counter[4] ;
 wire \i_uart_rx.cycle_counter[5] ;
 wire \i_uart_rx.cycle_counter[6] ;
 wire \i_uart_rx.cycle_counter[7] ;
 wire \i_uart_rx.cycle_counter[8] ;
 wire \i_uart_rx.fsm_state[0] ;
 wire \i_uart_rx.fsm_state[1] ;
 wire \i_uart_rx.fsm_state[2] ;
 wire \i_uart_rx.fsm_state[3] ;
 wire \i_uart_rx.recieved_data[0] ;
 wire \i_uart_rx.recieved_data[1] ;
 wire \i_uart_rx.recieved_data[2] ;
 wire \i_uart_rx.recieved_data[3] ;
 wire \i_uart_rx.recieved_data[4] ;
 wire \i_uart_rx.recieved_data[5] ;
 wire \i_uart_rx.recieved_data[6] ;
 wire \i_uart_rx.recieved_data[7] ;
 wire \i_uart_rx.rxd_reg[0] ;
 wire \i_uart_rx.rxd_reg[1] ;
 wire \i_uart_tx.cycle_counter[0] ;
 wire \i_uart_tx.cycle_counter[1] ;
 wire \i_uart_tx.cycle_counter[2] ;
 wire \i_uart_tx.cycle_counter[3] ;
 wire \i_uart_tx.cycle_counter[4] ;
 wire \i_uart_tx.cycle_counter[5] ;
 wire \i_uart_tx.cycle_counter[6] ;
 wire \i_uart_tx.cycle_counter[7] ;
 wire \i_uart_tx.cycle_counter[8] ;
 wire \i_uart_tx.data_to_send[0] ;
 wire \i_uart_tx.data_to_send[1] ;
 wire \i_uart_tx.data_to_send[2] ;
 wire \i_uart_tx.data_to_send[3] ;
 wire \i_uart_tx.data_to_send[4] ;
 wire \i_uart_tx.data_to_send[5] ;
 wire \i_uart_tx.data_to_send[6] ;
 wire \i_uart_tx.data_to_send[7] ;
 wire \i_uart_tx.fsm_state[0] ;
 wire \i_uart_tx.fsm_state[1] ;
 wire \i_uart_tx.fsm_state[2] ;
 wire \i_uart_tx.fsm_state[3] ;
 wire \i_uart_tx.txd_reg ;
 wire \i_wdt.counter[0] ;
 wire \i_wdt.counter[10] ;
 wire \i_wdt.counter[11] ;
 wire \i_wdt.counter[12] ;
 wire \i_wdt.counter[13] ;
 wire \i_wdt.counter[14] ;
 wire \i_wdt.counter[15] ;
 wire \i_wdt.counter[16] ;
 wire \i_wdt.counter[17] ;
 wire \i_wdt.counter[18] ;
 wire \i_wdt.counter[19] ;
 wire \i_wdt.counter[1] ;
 wire \i_wdt.counter[20] ;
 wire \i_wdt.counter[21] ;
 wire \i_wdt.counter[22] ;
 wire \i_wdt.counter[23] ;
 wire \i_wdt.counter[24] ;
 wire \i_wdt.counter[25] ;
 wire \i_wdt.counter[26] ;
 wire \i_wdt.counter[27] ;
 wire \i_wdt.counter[28] ;
 wire \i_wdt.counter[29] ;
 wire \i_wdt.counter[2] ;
 wire \i_wdt.counter[30] ;
 wire \i_wdt.counter[31] ;
 wire \i_wdt.counter[3] ;
 wire \i_wdt.counter[4] ;
 wire \i_wdt.counter[5] ;
 wire \i_wdt.counter[6] ;
 wire \i_wdt.counter[7] ;
 wire \i_wdt.counter[8] ;
 wire \i_wdt.counter[9] ;
 wire \i_wdt.enabled ;
 wire \i_wdt.wdt_reset ;
 wire \pps_count[0] ;
 wire \pps_count[10] ;
 wire \pps_count[11] ;
 wire \pps_count[12] ;
 wire \pps_count[13] ;
 wire \pps_count[14] ;
 wire \pps_count[15] ;
 wire \pps_count[1] ;
 wire \pps_count[2] ;
 wire \pps_count[3] ;
 wire \pps_count[4] ;
 wire \pps_count[5] ;
 wire \pps_count[6] ;
 wire \pps_count[7] ;
 wire \pps_count[8] ;
 wire \pps_count[9] ;
 wire pps_prev;
 wire \pps_sync[0] ;
 wire \pps_sync[1] ;
 wire \reset_hold_counter[0] ;
 wire \reset_hold_counter[1] ;
 wire \reset_hold_counter[2] ;
 wire \reset_hold_counter[3] ;
 wire \reset_hold_counter[4] ;
 wire \reset_hold_counter[5] ;
 wire \session_ms_div[0] ;
 wire \session_ms_div[1] ;
 wire \session_ms_div[2] ;
 wire \session_ms_div[3] ;
 wire \session_ms_div[4] ;
 wire \session_ms_div[5] ;
 wire \session_ms_div[6] ;
 wire \session_ms_div[7] ;
 wire \session_ms_div[8] ;
 wire \session_ms_div[9] ;
 wire \timer_count[0] ;
 wire \timer_count[10] ;
 wire \timer_count[11] ;
 wire \timer_count[12] ;
 wire \timer_count[13] ;
 wire \timer_count[14] ;
 wire \timer_count[15] ;
 wire \timer_count[16] ;
 wire \timer_count[17] ;
 wire \timer_count[18] ;
 wire \timer_count[19] ;
 wire \timer_count[1] ;
 wire \timer_count[20] ;
 wire \timer_count[21] ;
 wire \timer_count[22] ;
 wire \timer_count[23] ;
 wire \timer_count[24] ;
 wire \timer_count[25] ;
 wire \timer_count[26] ;
 wire \timer_count[27] ;
 wire \timer_count[28] ;
 wire \timer_count[29] ;
 wire \timer_count[2] ;
 wire \timer_count[30] ;
 wire \timer_count[31] ;
 wire \timer_count[3] ;
 wire \timer_count[4] ;
 wire \timer_count[5] ;
 wire \timer_count[6] ;
 wire \timer_count[7] ;
 wire \timer_count[8] ;
 wire \timer_count[9] ;
 wire timer_irq;
 wire \us_divider[0] ;
 wire \us_divider[1] ;
 wire \us_divider[2] ;
 wire \us_divider[3] ;
 wire \us_divider[4] ;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_88_clk_regs;
 wire clknet_leaf_89_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_106_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_leaf_112_clk_regs;
 wire clknet_leaf_113_clk_regs;
 wire clknet_leaf_114_clk_regs;
 wire clknet_leaf_115_clk_regs;
 wire clknet_leaf_116_clk_regs;
 wire clknet_leaf_117_clk_regs;
 wire clknet_leaf_118_clk_regs;
 wire clknet_leaf_119_clk_regs;
 wire clknet_leaf_120_clk_regs;
 wire clknet_leaf_121_clk_regs;
 wire clknet_leaf_122_clk_regs;
 wire clknet_leaf_123_clk_regs;
 wire clknet_leaf_124_clk_regs;
 wire clknet_leaf_125_clk_regs;
 wire clknet_leaf_126_clk_regs;
 wire clknet_leaf_127_clk_regs;
 wire clknet_leaf_128_clk_regs;
 wire clknet_leaf_129_clk_regs;
 wire clknet_leaf_130_clk_regs;
 wire clknet_leaf_131_clk_regs;
 wire clknet_leaf_132_clk_regs;
 wire clknet_leaf_133_clk_regs;
 wire clknet_leaf_134_clk_regs;
 wire clknet_leaf_135_clk_regs;
 wire clknet_leaf_136_clk_regs;
 wire clknet_leaf_137_clk_regs;
 wire clknet_leaf_138_clk_regs;
 wire clknet_leaf_139_clk_regs;
 wire clknet_leaf_140_clk_regs;
 wire clknet_leaf_141_clk_regs;
 wire clknet_leaf_142_clk_regs;
 wire clknet_leaf_143_clk_regs;
 wire clknet_leaf_144_clk_regs;
 wire clknet_leaf_145_clk_regs;
 wire clknet_leaf_146_clk_regs;
 wire clknet_leaf_147_clk_regs;
 wire clknet_leaf_148_clk_regs;
 wire clknet_leaf_149_clk_regs;
 wire clknet_leaf_150_clk_regs;
 wire clknet_leaf_151_clk_regs;
 wire clknet_leaf_152_clk_regs;
 wire clknet_leaf_153_clk_regs;
 wire clknet_leaf_154_clk_regs;
 wire clknet_leaf_155_clk_regs;
 wire clknet_leaf_156_clk_regs;
 wire clknet_leaf_157_clk_regs;
 wire clknet_leaf_158_clk_regs;
 wire clknet_leaf_159_clk_regs;
 wire clknet_leaf_160_clk_regs;
 wire clknet_leaf_161_clk_regs;
 wire clknet_leaf_162_clk_regs;
 wire clknet_leaf_163_clk_regs;
 wire clknet_leaf_164_clk_regs;
 wire clknet_leaf_165_clk_regs;
 wire clknet_leaf_166_clk_regs;
 wire clknet_leaf_167_clk_regs;
 wire clknet_leaf_168_clk_regs;
 wire clknet_leaf_169_clk_regs;
 wire clknet_leaf_170_clk_regs;
 wire clknet_leaf_171_clk_regs;
 wire clknet_leaf_172_clk_regs;
 wire clknet_leaf_173_clk_regs;
 wire clknet_leaf_174_clk_regs;
 wire clknet_leaf_175_clk_regs;
 wire clknet_leaf_176_clk_regs;
 wire clknet_leaf_177_clk_regs;
 wire clknet_leaf_178_clk_regs;
 wire clknet_leaf_179_clk_regs;
 wire clknet_leaf_180_clk_regs;
 wire clknet_leaf_181_clk_regs;
 wire clknet_leaf_182_clk_regs;
 wire clknet_leaf_183_clk_regs;
 wire clknet_leaf_184_clk_regs;
 wire clknet_leaf_185_clk_regs;
 wire clknet_leaf_186_clk_regs;
 wire clknet_leaf_187_clk_regs;
 wire clknet_leaf_188_clk_regs;
 wire clknet_leaf_189_clk_regs;
 wire clknet_leaf_190_clk_regs;
 wire clknet_leaf_191_clk_regs;
 wire clknet_leaf_192_clk_regs;
 wire clknet_leaf_193_clk_regs;
 wire clknet_leaf_194_clk_regs;
 wire clknet_leaf_195_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_3_0_0_clk_regs;
 wire clknet_3_1_0_clk_regs;
 wire clknet_3_2_0_clk_regs;
 wire clknet_3_3_0_clk_regs;
 wire clknet_3_4_0_clk_regs;
 wire clknet_3_5_0_clk_regs;
 wire clknet_3_6_0_clk_regs;
 wire clknet_3_7_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4181;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4189;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4195;
 wire net4196;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4202;
 wire net4203;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4207;
 wire net4208;
 wire net4209;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4213;
 wire net4214;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4228;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4236;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4241;
 wire net4242;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4246;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4255;
 wire net4256;
 wire net4257;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4276;
 wire net4277;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4285;
 wire net4286;
 wire net4287;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4291;
 wire net4292;
 wire net4293;
 wire net4294;
 wire net4295;
 wire net4296;
 wire net4297;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4301;
 wire net4302;
 wire net4303;
 wire net4304;
 wire net4305;
 wire net4306;
 wire net4307;
 wire net4308;
 wire net4309;
 wire net4310;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4329;
 wire net4330;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4341;
 wire net4342;
 wire net4343;
 wire net4344;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4348;
 wire net4349;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4353;
 wire net4354;
 wire net4355;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4362;
 wire net4363;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4369;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4388;
 wire net4389;
 wire net4390;
 wire net4391;
 wire net4392;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4397;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4401;
 wire net4402;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4409;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4421;
 wire net4422;
 wire net4423;
 wire net4424;
 wire net4425;
 wire net4426;
 wire net4427;
 wire net4428;
 wire net4429;
 wire net4430;
 wire net4431;
 wire net4432;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4442;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4446;
 wire net4447;
 wire net4448;
 wire net4449;
 wire net4450;
 wire net4451;
 wire net4452;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4456;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4460;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4464;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4480;
 wire net4481;
 wire net4482;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4498;
 wire net4499;
 wire net4500;
 wire net4501;
 wire net4502;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4506;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4523;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4528;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4539;
 wire net4540;
 wire net4541;
 wire net4542;
 wire net4543;
 wire net4544;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4557;
 wire net4558;
 wire net4559;
 wire net4560;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4570;
 wire net4571;
 wire net4572;
 wire net4573;
 wire net4574;
 wire net4575;
 wire net4576;
 wire net4577;
 wire net4578;
 wire net4579;
 wire net4580;
 wire net4581;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4585;
 wire net4586;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4592;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4596;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4604;
 wire net4605;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4609;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4623;
 wire net4624;
 wire net4625;
 wire net4626;
 wire net4627;
 wire net4628;
 wire net4629;
 wire net4630;
 wire net4631;
 wire net4632;
 wire net4633;
 wire net4634;
 wire net4635;
 wire net4636;
 wire net4637;
 wire net4638;
 wire net4639;
 wire net4640;
 wire net4641;
 wire net4642;
 wire net4643;
 wire net4644;
 wire net4645;
 wire net4646;
 wire net4647;
 wire net4648;
 wire net4649;
 wire net4650;
 wire net4651;
 wire net4652;
 wire net4653;
 wire net4654;
 wire net4655;
 wire net4656;
 wire net4657;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4662;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4674;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4683;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4689;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net4693;
 wire net4694;
 wire net4695;
 wire net4696;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4708;
 wire net4709;
 wire net4710;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4714;
 wire net4715;
 wire net4716;
 wire net4717;
 wire net4718;
 wire net4719;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4724;
 wire net4725;
 wire net4726;
 wire net4727;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4735;
 wire net4736;
 wire net4737;
 wire net4738;
 wire net4739;
 wire net4740;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4747;
 wire net4748;
 wire net4749;
 wire net4750;
 wire net4751;
 wire net4752;
 wire net4753;
 wire net4754;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4758;
 wire net4759;
 wire net4760;
 wire net4761;
 wire net4762;
 wire net4763;
 wire net4764;
 wire net4765;
 wire net4766;
 wire net4767;
 wire net4768;
 wire net4769;
 wire net4770;
 wire net4771;
 wire net4772;
 wire net4773;
 wire net4774;
 wire net4775;
 wire net4776;
 wire net4777;
 wire net4778;
 wire net4779;
 wire net4780;
 wire net4781;
 wire net4782;
 wire net4783;
 wire net4784;
 wire net4785;
 wire net4786;
 wire net4787;
 wire net4788;
 wire net4789;
 wire net4790;
 wire net4791;
 wire net4792;
 wire net4793;
 wire net4794;
 wire net4795;
 wire net4796;
 wire net4797;
 wire net4798;
 wire net4799;
 wire net4800;
 wire net4801;
 wire net4802;
 wire net4803;
 wire net4804;
 wire net4805;
 wire net4806;
 wire net4807;
 wire net4808;
 wire net4809;
 wire net4810;
 wire net4811;
 wire net4812;
 wire net4813;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4825;
 wire net4826;
 wire net4827;
 wire net4828;
 wire net4829;
 wire net4830;
 wire net4831;
 wire net4832;
 wire net4833;
 wire net4834;
 wire net4835;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4839;
 wire net4840;
 wire net4841;
 wire net4842;
 wire net4843;
 wire net4844;
 wire net4845;
 wire net4846;
 wire net4847;
 wire net4848;
 wire net4849;
 wire net4850;
 wire net4851;
 wire net4852;
 wire net4853;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4858;
 wire net4859;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4879;
 wire net4880;
 wire net4881;
 wire net4882;
 wire net4883;
 wire net4884;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4915;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4935;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4997;
 wire net4998;
 wire net4999;
 wire net5000;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5011;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5023;
 wire net5024;
 wire net5025;
 wire net5026;
 wire net5027;
 wire net5028;
 wire net5029;
 wire net5030;
 wire net5031;
 wire net5032;
 wire net5033;
 wire net5034;
 wire net5035;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5162;
 wire net5163;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5190;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5200;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5211;
 wire net5212;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5227;
 wire net5228;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5235;
 wire net5236;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5241;
 wire net5242;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5251;
 wire net5252;
 wire net5253;
 wire net5254;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5260;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5282;
 wire net5283;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5287;
 wire net5288;
 wire net5289;
 wire net5290;
 wire net5291;
 wire net5292;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5298;
 wire net5299;
 wire net5300;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5327;
 wire net5328;
 wire net5329;
 wire net5330;
 wire net5331;
 wire net5332;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5346;
 wire net5347;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire net5359;
 wire net5360;
 wire net5361;
 wire net5362;
 wire net5363;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;

 sg13g2_inv_1 _09066_ (.Y(_01741_),
    .A(net4637));
 sg13g2_inv_1 _09067_ (.Y(_01742_),
    .A(net3577));
 sg13g2_inv_1 _09068_ (.Y(_01743_),
    .A(\i_latch_mem.genblk1[0].l_ram.data_out[6] ));
 sg13g2_inv_1 _09069_ (.Y(_01744_),
    .A(\i_latch_mem.genblk1[0].l_ram.data_out[5] ));
 sg13g2_inv_1 _09070_ (.Y(_01745_),
    .A(\i_latch_mem.genblk1[0].l_ram.data_out[4] ));
 sg13g2_inv_1 _09071_ (.Y(_01746_),
    .A(\i_spi.clock_count[3] ));
 sg13g2_inv_2 _09072_ (.Y(_01747_),
    .A(net2454));
 sg13g2_inv_1 _09073_ (.Y(_01748_),
    .A(\i_spi.clock_count[1] ));
 sg13g2_inv_1 _09074_ (.Y(_01749_),
    .A(net4740));
 sg13g2_inv_1 _09075_ (.Y(_01750_),
    .A(net4787));
 sg13g2_inv_1 _09076_ (.Y(_01751_),
    .A(\i_uart_rx.rxd_reg[0] ));
 sg13g2_inv_1 _09077_ (.Y(_01752_),
    .A(net4715));
 sg13g2_inv_1 _09078_ (.Y(_01753_),
    .A(net4762));
 sg13g2_inv_2 _09079_ (.Y(_01754_),
    .A(net5040));
 sg13g2_inv_1 _09080_ (.Y(_01755_),
    .A(net4646));
 sg13g2_inv_1 _09081_ (.Y(_01756_),
    .A(net4990));
 sg13g2_inv_1 _09082_ (.Y(_01757_),
    .A(\crc16_read[6] ));
 sg13g2_inv_1 _09083_ (.Y(_01758_),
    .A(\crc16_read[5] ));
 sg13g2_inv_1 _09084_ (.Y(_01759_),
    .A(net4719));
 sg13g2_inv_1 _09085_ (.Y(_01760_),
    .A(net4964));
 sg13g2_inv_1 _09086_ (.Y(_01761_),
    .A(net4874));
 sg13g2_inv_1 _09087_ (.Y(_01762_),
    .A(\crc16_read[1] ));
 sg13g2_inv_1 _09088_ (.Y(_01763_),
    .A(\crc16_read[0] ));
 sg13g2_inv_1 _09089_ (.Y(_01764_),
    .A(net4203));
 sg13g2_inv_1 _09090_ (.Y(_01765_),
    .A(net4313));
 sg13g2_inv_1 _09091_ (.Y(_01766_),
    .A(net3974));
 sg13g2_inv_1 _09092_ (.Y(_01767_),
    .A(net4112));
 sg13g2_inv_1 _09093_ (.Y(_01768_),
    .A(net4064));
 sg13g2_inv_1 _09094_ (.Y(_01769_),
    .A(net4423));
 sg13g2_inv_1 _09095_ (.Y(_01770_),
    .A(net4026));
 sg13g2_inv_1 _09096_ (.Y(_01771_),
    .A(net4486));
 sg13g2_inv_8 _09097_ (.Y(_01772_),
    .A(net2551));
 sg13g2_inv_8 _09098_ (.Y(_01773_),
    .A(net2552));
 sg13g2_inv_8 _09099_ (.Y(_01774_),
    .A(net2553));
 sg13g2_inv_8 _09100_ (.Y(_01775_),
    .A(net2554));
 sg13g2_inv_1 _09101_ (.Y(_01776_),
    .A(net2555));
 sg13g2_inv_8 _09102_ (.Y(_01777_),
    .A(net5012));
 sg13g2_inv_1 _09103_ (.Y(_01778_),
    .A(net2558));
 sg13g2_inv_8 _09104_ (.Y(_01779_),
    .A(net4681));
 sg13g2_inv_8 _09105_ (.Y(_01780_),
    .A(net2547));
 sg13g2_inv_1 _09106_ (.Y(_01781_),
    .A(net4055));
 sg13g2_inv_2 _09107_ (.Y(_01782_),
    .A(net3800));
 sg13g2_inv_1 _09108_ (.Y(_01783_),
    .A(net4258));
 sg13g2_inv_1 _09109_ (.Y(_01784_),
    .A(net4068));
 sg13g2_inv_1 _09110_ (.Y(_01785_),
    .A(net4331));
 sg13g2_inv_1 _09111_ (.Y(_01786_),
    .A(net4359));
 sg13g2_inv_1 _09112_ (.Y(_01787_),
    .A(net4223));
 sg13g2_inv_2 _09113_ (.Y(_01788_),
    .A(net3751));
 sg13g2_inv_1 _09114_ (.Y(_01789_),
    .A(net3988));
 sg13g2_inv_4 _09115_ (.A(net4979),
    .Y(_01790_));
 sg13g2_inv_1 _09116_ (.Y(_01791_),
    .A(\i2c_config_out[14] ));
 sg13g2_inv_4 _09117_ (.A(net4962),
    .Y(_01792_));
 sg13g2_inv_4 _09118_ (.A(net5053),
    .Y(_01793_));
 sg13g2_inv_2 _09119_ (.Y(_01794_),
    .A(net5104));
 sg13g2_inv_4 _09120_ (.A(net4958),
    .Y(_01795_));
 sg13g2_inv_4 _09121_ (.A(net2548),
    .Y(_01796_));
 sg13g2_inv_4 _09122_ (.A(net2550),
    .Y(_01797_));
 sg13g2_inv_1 _09123_ (.Y(_01798_),
    .A(net4897));
 sg13g2_inv_1 _09124_ (.Y(_01799_),
    .A(net4862));
 sg13g2_inv_1 _09125_ (.Y(_01800_),
    .A(\i2c_config_out[3] ));
 sg13g2_inv_1 _09126_ (.Y(_01801_),
    .A(\i2c_config_out[2] ));
 sg13g2_inv_2 _09127_ (.Y(_01802_),
    .A(net4369));
 sg13g2_inv_1 _09128_ (.Y(_01803_),
    .A(net4651));
 sg13g2_inv_2 _09129_ (.Y(_01804_),
    .A(\i_i2c_peri.i_i2c.phy_state_reg[0] ));
 sg13g2_inv_1 _09130_ (.Y(_01805_),
    .A(net4073));
 sg13g2_inv_1 _09131_ (.Y(_01806_),
    .A(net3409));
 sg13g2_inv_2 _09132_ (.Y(_01807_),
    .A(net2471));
 sg13g2_inv_2 _09133_ (.Y(_01808_),
    .A(net4684));
 sg13g2_inv_1 _09134_ (.Y(_01809_),
    .A(net2492));
 sg13g2_inv_2 _09135_ (.Y(_01810_),
    .A(net5345));
 sg13g2_inv_1 _09136_ (.Y(_01811_),
    .A(net4227));
 sg13g2_inv_2 _09137_ (.Y(_01812_),
    .A(net5020));
 sg13g2_inv_1 _09138_ (.Y(_01813_),
    .A(net4077));
 sg13g2_inv_1 _09139_ (.Y(_01814_),
    .A(net5005));
 sg13g2_inv_1 _09140_ (.Y(_01815_),
    .A(net4382));
 sg13g2_inv_2 _09141_ (.Y(_01816_),
    .A(net5055));
 sg13g2_inv_1 _09142_ (.Y(_01817_),
    .A(net4071));
 sg13g2_inv_1 _09143_ (.Y(_01818_),
    .A(net4927));
 sg13g2_inv_1 _09144_ (.Y(_01819_),
    .A(net4327));
 sg13g2_inv_1 _09145_ (.Y(_01820_),
    .A(net5079));
 sg13g2_inv_1 _09146_ (.Y(_01821_),
    .A(net4324));
 sg13g2_inv_1 _09147_ (.Y(_01822_),
    .A(net5054));
 sg13g2_inv_1 _09148_ (.Y(_01823_),
    .A(net4393));
 sg13g2_inv_1 _09149_ (.Y(_01824_),
    .A(net5071));
 sg13g2_inv_1 _09150_ (.Y(_01825_),
    .A(net4189));
 sg13g2_inv_1 _09151_ (.Y(_01826_),
    .A(net4986));
 sg13g2_inv_1 _09152_ (.Y(_01827_),
    .A(net4134));
 sg13g2_inv_1 _09153_ (.Y(_01828_),
    .A(net4928));
 sg13g2_inv_1 _09154_ (.Y(_01829_),
    .A(net4098));
 sg13g2_inv_2 _09155_ (.Y(_01830_),
    .A(net4905));
 sg13g2_inv_1 _09156_ (.Y(_01831_),
    .A(net4155));
 sg13g2_inv_1 _09157_ (.Y(_01832_),
    .A(net4933));
 sg13g2_inv_1 _09158_ (.Y(_01833_),
    .A(net4007));
 sg13g2_inv_1 _09159_ (.Y(_01834_),
    .A(net4994));
 sg13g2_inv_1 _09160_ (.Y(_01835_),
    .A(net4317));
 sg13g2_inv_4 _09161_ (.A(net4912),
    .Y(_01836_));
 sg13g2_inv_1 _09162_ (.Y(_01837_),
    .A(net4016));
 sg13g2_inv_4 _09163_ (.A(net4877),
    .Y(_01838_));
 sg13g2_inv_1 _09164_ (.Y(_01839_),
    .A(net3962));
 sg13g2_inv_4 _09165_ (.A(net4914),
    .Y(_01840_));
 sg13g2_inv_1 _09166_ (.Y(_01841_),
    .A(net4005));
 sg13g2_inv_4 _09167_ (.A(net4892),
    .Y(_01842_));
 sg13g2_inv_1 _09168_ (.Y(_01843_),
    .A(net4118));
 sg13g2_inv_1 _09169_ (.Y(_01844_),
    .A(net4029));
 sg13g2_inv_1 _09170_ (.Y(_01845_),
    .A(net4221));
 sg13g2_inv_1 _09171_ (.Y(_01846_),
    .A(\i_seal.value_reg[12] ));
 sg13g2_inv_1 _09172_ (.Y(_01847_),
    .A(net4430));
 sg13g2_inv_1 _09173_ (.Y(_01848_),
    .A(net4267));
 sg13g2_inv_1 _09174_ (.Y(_01849_),
    .A(net4197));
 sg13g2_inv_1 _09175_ (.Y(_01850_),
    .A(net3785));
 sg13g2_inv_1 _09176_ (.Y(_01851_),
    .A(net3926));
 sg13g2_inv_1 _09177_ (.Y(_01852_),
    .A(net3950));
 sg13g2_inv_1 _09178_ (.Y(_01853_),
    .A(\i_seal.value_reg[5] ));
 sg13g2_inv_1 _09179_ (.Y(_01854_),
    .A(net3956));
 sg13g2_inv_1 _09180_ (.Y(_01855_),
    .A(net4479));
 sg13g2_inv_1 _09181_ (.Y(_01856_),
    .A(net4420));
 sg13g2_inv_1 _09182_ (.Y(_01857_),
    .A(net4572));
 sg13g2_inv_1 _09183_ (.Y(_01858_),
    .A(\i_seal.value_reg[0] ));
 sg13g2_inv_1 _09184_ (.Y(_01859_),
    .A(net4037));
 sg13g2_inv_1 _09185_ (.Y(_01860_),
    .A(net3912));
 sg13g2_inv_1 _09186_ (.Y(_01861_),
    .A(net4047));
 sg13g2_inv_1 _09187_ (.Y(_01862_),
    .A(net3937));
 sg13g2_inv_1 _09188_ (.Y(_01863_),
    .A(net3846));
 sg13g2_inv_1 _09189_ (.Y(_01864_),
    .A(net3685));
 sg13g2_inv_1 _09190_ (.Y(_01865_),
    .A(net4094));
 sg13g2_inv_1 _09191_ (.Y(_01866_),
    .A(net3539));
 sg13g2_inv_1 _09192_ (.Y(_01867_),
    .A(net3844));
 sg13g2_inv_1 _09193_ (.Y(_01868_),
    .A(net3919));
 sg13g2_inv_1 _09194_ (.Y(_01869_),
    .A(net4142));
 sg13g2_inv_1 _09195_ (.Y(_01870_),
    .A(net3917));
 sg13g2_inv_1 _09196_ (.Y(_01871_),
    .A(net3982));
 sg13g2_inv_1 _09197_ (.Y(_01872_),
    .A(net3550));
 sg13g2_inv_1 _09198_ (.Y(_01873_),
    .A(net3825));
 sg13g2_inv_1 _09199_ (.Y(_01874_),
    .A(net3979));
 sg13g2_inv_1 _09200_ (.Y(_01875_),
    .A(net4173));
 sg13g2_inv_1 _09201_ (.Y(_01876_),
    .A(net3673));
 sg13g2_inv_1 _09202_ (.Y(_01877_),
    .A(net4365));
 sg13g2_inv_1 _09203_ (.Y(_01878_),
    .A(net3999));
 sg13g2_inv_1 _09204_ (.Y(_01879_),
    .A(net4559));
 sg13g2_inv_1 _09205_ (.Y(_01880_),
    .A(net4031));
 sg13g2_inv_1 _09206_ (.Y(_01881_),
    .A(net4336));
 sg13g2_inv_1 _09207_ (.Y(_01882_),
    .A(net3835));
 sg13g2_inv_1 _09208_ (.Y(_01883_),
    .A(net4543));
 sg13g2_inv_1 _09209_ (.Y(_01884_),
    .A(net3665));
 sg13g2_inv_1 _09210_ (.Y(_01885_),
    .A(net4059));
 sg13g2_inv_1 _09211_ (.Y(_01886_),
    .A(net3758));
 sg13g2_inv_1 _09212_ (.Y(_01887_),
    .A(net4015));
 sg13g2_inv_1 _09213_ (.Y(_01888_),
    .A(net3971));
 sg13g2_inv_1 _09214_ (.Y(_01889_),
    .A(net4147));
 sg13g2_inv_1 _09215_ (.Y(_01890_),
    .A(net4039));
 sg13g2_inv_1 _09216_ (.Y(_01891_),
    .A(\i_seal.cur_mono[16] ));
 sg13g2_inv_1 _09217_ (.Y(_01892_),
    .A(net3892));
 sg13g2_inv_1 _09218_ (.Y(_01893_),
    .A(net3870));
 sg13g2_inv_1 _09219_ (.Y(_01894_),
    .A(net4777));
 sg13g2_inv_1 _09220_ (.Y(_01895_),
    .A(net3864));
 sg13g2_inv_2 _09221_ (.Y(_01896_),
    .A(net4181));
 sg13g2_inv_1 _09222_ (.Y(_01897_),
    .A(net3901));
 sg13g2_inv_1 _09223_ (.Y(_01898_),
    .A(net3895));
 sg13g2_inv_1 _09224_ (.Y(_01899_),
    .A(net4273));
 sg13g2_inv_1 _09225_ (.Y(_01900_),
    .A(net4555));
 sg13g2_inv_1 _09226_ (.Y(_01901_),
    .A(net3727));
 sg13g2_inv_1 _09227_ (.Y(_01902_),
    .A(\i_seal.cur_mono[9] ));
 sg13g2_inv_1 _09228_ (.Y(_01903_),
    .A(net3654));
 sg13g2_inv_1 _09229_ (.Y(_01904_),
    .A(net3986));
 sg13g2_inv_1 _09230_ (.Y(_01905_),
    .A(net3931));
 sg13g2_inv_2 _09231_ (.Y(_01906_),
    .A(net4253));
 sg13g2_inv_1 _09232_ (.Y(_01907_),
    .A(net4308));
 sg13g2_inv_1 _09233_ (.Y(_01908_),
    .A(net4576));
 sg13g2_inv_1 _09234_ (.Y(_01909_),
    .A(net3713));
 sg13g2_inv_1 _09235_ (.Y(_01910_),
    .A(net4067));
 sg13g2_inv_1 _09236_ (.Y(_01911_),
    .A(net3889));
 sg13g2_inv_1 _09237_ (.Y(_01912_),
    .A(net4114));
 sg13g2_inv_1 _09238_ (.Y(_01913_),
    .A(net4319));
 sg13g2_inv_1 _09239_ (.Y(_01914_),
    .A(net4626));
 sg13g2_inv_2 _09240_ (.Y(_01915_),
    .A(net3954));
 sg13g2_inv_1 _09241_ (.Y(_01916_),
    .A(net4079));
 sg13g2_inv_1 _09242_ (.Y(_01917_),
    .A(net4052));
 sg13g2_inv_1 _09243_ (.Y(_01918_),
    .A(net4110));
 sg13g2_inv_1 _09244_ (.Y(_01919_),
    .A(net4120));
 sg13g2_inv_1 _09245_ (.Y(_01920_),
    .A(net4187));
 sg13g2_inv_2 _09246_ (.Y(_01921_),
    .A(net4202));
 sg13g2_inv_1 _09247_ (.Y(_01922_),
    .A(net3990));
 sg13g2_inv_1 _09248_ (.Y(_01923_),
    .A(net3928));
 sg13g2_inv_2 _09249_ (.Y(_01924_),
    .A(net3885));
 sg13g2_inv_1 _09250_ (.Y(_01925_),
    .A(net3779));
 sg13g2_inv_1 _09251_ (.Y(_01926_),
    .A(net4138));
 sg13g2_inv_1 _09252_ (.Y(_01927_),
    .A(net4311));
 sg13g2_inv_1 _09253_ (.Y(_01928_),
    .A(net3789));
 sg13g2_inv_1 _09254_ (.Y(_01929_),
    .A(net3899));
 sg13g2_inv_1 _09255_ (.Y(_01930_),
    .A(\i_seal.sealed_mono[27] ));
 sg13g2_inv_1 _09256_ (.Y(_01931_),
    .A(\i_seal.sealed_mono[16] ));
 sg13g2_inv_2 _09257_ (.Y(_01932_),
    .A(net3946));
 sg13g2_inv_2 _09258_ (.Y(_01933_),
    .A(\i_seal.sealed_mono[14] ));
 sg13g2_inv_2 _09259_ (.Y(_01934_),
    .A(\i_seal.sealed_mono[13] ));
 sg13g2_inv_2 _09260_ (.Y(_01935_),
    .A(net3765));
 sg13g2_inv_2 _09261_ (.Y(_01936_),
    .A(net3922));
 sg13g2_inv_1 _09262_ (.Y(_01937_),
    .A(\i_seal.sealed_mono[10] ));
 sg13g2_inv_1 _09263_ (.Y(_01938_),
    .A(\i_seal.sealed_mono[9] ));
 sg13g2_inv_1 _09264_ (.Y(_01939_),
    .A(net3568));
 sg13g2_inv_1 _09265_ (.Y(_01940_),
    .A(net3588));
 sg13g2_inv_1 _09266_ (.Y(_01941_),
    .A(net4751));
 sg13g2_inv_1 _09267_ (.Y(_01942_),
    .A(net3668));
 sg13g2_inv_1 _09268_ (.Y(_01943_),
    .A(net3544));
 sg13g2_inv_1 _09269_ (.Y(_01944_),
    .A(net3564));
 sg13g2_inv_1 _09270_ (.Y(_01945_),
    .A(net3677));
 sg13g2_inv_1 _09271_ (.Y(_01946_),
    .A(net3554));
 sg13g2_inv_2 _09272_ (.Y(_01947_),
    .A(net5120));
 sg13g2_inv_1 _09273_ (.Y(_01948_),
    .A(net4363));
 sg13g2_inv_1 _09274_ (.Y(_01949_),
    .A(net5222));
 sg13g2_inv_1 _09275_ (.Y(_01950_),
    .A(net5087));
 sg13g2_inv_1 _09276_ (.Y(_01951_),
    .A(net5176));
 sg13g2_inv_1 _09277_ (.Y(_01952_),
    .A(net5056));
 sg13g2_inv_1 _09278_ (.Y(_01953_),
    .A(net5239));
 sg13g2_inv_1 _09279_ (.Y(_01954_),
    .A(net5332));
 sg13g2_inv_1 _09280_ (.Y(_01955_),
    .A(net5309));
 sg13g2_inv_1 _09281_ (.Y(_01956_),
    .A(net4432));
 sg13g2_inv_1 _09282_ (.Y(_01957_),
    .A(net5125));
 sg13g2_inv_1 _09283_ (.Y(_01958_),
    .A(net3481));
 sg13g2_inv_1 _09284_ (.Y(_01959_),
    .A(net4825));
 sg13g2_inv_2 _09285_ (.Y(_01960_),
    .A(net2498));
 sg13g2_inv_1 _09286_ (.Y(_01961_),
    .A(net3960));
 sg13g2_inv_4 _09287_ (.A(net5061),
    .Y(_01962_));
 sg13g2_inv_1 _09288_ (.Y(_01963_),
    .A(net2510));
 sg13g2_inv_2 _09289_ (.Y(_01964_),
    .A(net4742));
 sg13g2_inv_1 _09290_ (.Y(_01965_),
    .A(\i_tinyqv.cpu.is_jalr ));
 sg13g2_inv_4 _09291_ (.A(net4710),
    .Y(_01966_));
 sg13g2_inv_2 _09292_ (.Y(_01967_),
    .A(net2564));
 sg13g2_inv_1 _09293_ (.Y(_01968_),
    .A(\i_tinyqv.cpu.instr_data_start[22] ));
 sg13g2_inv_2 _09294_ (.Y(_01969_),
    .A(net5145));
 sg13g2_inv_1 _09295_ (.Y(_01970_),
    .A(net2565));
 sg13g2_inv_4 _09296_ (.A(net5256),
    .Y(_01971_));
 sg13g2_inv_1 _09297_ (.Y(_01972_),
    .A(\i_tinyqv.cpu.instr_data_start[15] ));
 sg13g2_inv_1 _09298_ (.Y(_01973_),
    .A(net2568));
 sg13g2_inv_1 _09299_ (.Y(_01974_),
    .A(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_inv_2 _09300_ (.Y(_01975_),
    .A(net5167));
 sg13g2_inv_1 _09301_ (.Y(_01976_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ));
 sg13g2_inv_2 _09302_ (.Y(_01977_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ));
 sg13g2_inv_1 _09303_ (.Y(_01978_),
    .A(\i_spi.clock_divider[3] ));
 sg13g2_inv_1 _09304_ (.Y(_01979_),
    .A(\i_spi.read_latency ));
 sg13g2_inv_1 _09305_ (.Y(_01980_),
    .A(net2608));
 sg13g2_inv_2 _09306_ (.Y(_01981_),
    .A(net2610));
 sg13g2_inv_4 _09307_ (.A(net4625),
    .Y(_01982_));
 sg13g2_inv_1 _09308_ (.Y(_01983_),
    .A(net2612));
 sg13g2_inv_1 _09309_ (.Y(_01984_),
    .A(net5280));
 sg13g2_inv_1 _09310_ (.Y(_01985_),
    .A(net5342));
 sg13g2_inv_1 _09311_ (.Y(_01986_),
    .A(net3935));
 sg13g2_inv_1 _09312_ (.Y(_01987_),
    .A(net4829));
 sg13g2_inv_1 _09313_ (.Y(_01988_),
    .A(net3408));
 sg13g2_inv_2 _09314_ (.Y(_01989_),
    .A(net2539));
 sg13g2_inv_1 _09315_ (.Y(_01990_),
    .A(net2536));
 sg13g2_inv_1 _09316_ (.Y(_01991_),
    .A(\i_tinyqv.cpu.alu_op[3] ));
 sg13g2_inv_1 _09317_ (.Y(_01992_),
    .A(net2524));
 sg13g2_inv_1 _09318_ (.Y(_01993_),
    .A(net5209));
 sg13g2_inv_2 _09319_ (.Y(_01994_),
    .A(net2514));
 sg13g2_inv_2 _09320_ (.Y(_01995_),
    .A(net2515));
 sg13g2_inv_2 _09321_ (.Y(_01996_),
    .A(net2516));
 sg13g2_inv_1 _09322_ (.Y(_01997_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_inv_1 _09323_ (.Y(_01998_),
    .A(\i_tinyqv.cpu.imm[18] ));
 sg13g2_inv_1 _09324_ (.Y(_01999_),
    .A(net4686));
 sg13g2_inv_1 _09325_ (.Y(_02000_),
    .A(net4283));
 sg13g2_inv_2 _09326_ (.Y(_02001_),
    .A(net2529));
 sg13g2_inv_2 _09327_ (.Y(_02002_),
    .A(\i_tinyqv.cpu.instr_write_offset[1] ));
 sg13g2_inv_2 _09328_ (.Y(_02003_),
    .A(\i_tinyqv.mem.q_ctrl.data_ready ));
 sg13g2_inv_1 _09329_ (.Y(_02004_),
    .A(net3772));
 sg13g2_inv_1 _09330_ (.Y(_02005_),
    .A(net3679));
 sg13g2_inv_1 _09331_ (.Y(_02006_),
    .A(net3976));
 sg13g2_inv_1 _09332_ (.Y(_02007_),
    .A(net3841));
 sg13g2_inv_1 _09333_ (.Y(_02008_),
    .A(net3742));
 sg13g2_inv_1 _09334_ (.Y(_02009_),
    .A(net3807));
 sg13g2_inv_1 _09335_ (.Y(_02010_),
    .A(net4049));
 sg13g2_inv_1 _09336_ (.Y(_02011_),
    .A(net3910));
 sg13g2_inv_1 _09337_ (.Y(_02012_),
    .A(net2673));
 sg13g2_inv_8 _09338_ (.Y(_02013_),
    .A(\addr[2] ));
 sg13g2_inv_4 _09339_ (.A(\addr[4] ),
    .Y(_02014_));
 sg13g2_inv_2 _09340_ (.Y(_02015_),
    .A(\addr[6] ));
 sg13g2_inv_1 _09341_ (.Y(_02016_),
    .A(net4566));
 sg13g2_inv_1 _09342_ (.Y(_02017_),
    .A(\i_i2c_peri.i_i2c.addr_reg[3] ));
 sg13g2_inv_1 _09343_ (.Y(_02018_),
    .A(net3652));
 sg13g2_inv_1 _09344_ (.Y(_02019_),
    .A(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ));
 sg13g2_inv_1 _09345_ (.Y(_02020_),
    .A(\i_latch_mem.data_ready ));
 sg13g2_inv_1 _09346_ (.Y(_02021_),
    .A(\i_tinyqv.cpu.instr_fetch_stopped ));
 sg13g2_inv_2 _09347_ (.Y(_02022_),
    .A(net3397));
 sg13g2_inv_2 _09348_ (.Y(_02023_),
    .A(net4865));
 sg13g2_inv_1 _09349_ (.Y(_02024_),
    .A(net4271));
 sg13g2_inv_1 _09350_ (.Y(_02025_),
    .A(\i_seal.crc_feed ));
 sg13g2_inv_1 _09351_ (.Y(_02026_),
    .A(net1));
 sg13g2_inv_1 _09352_ (.Y(_02027_),
    .A(net4339));
 sg13g2_inv_1 _09353_ (.Y(_02028_),
    .A(net4640));
 sg13g2_inv_1 _09354_ (.Y(_02029_),
    .A(net4535));
 sg13g2_inv_1 _09355_ (.Y(_02030_),
    .A(net4374));
 sg13g2_inv_1 _09356_ (.Y(_02031_),
    .A(net4367));
 sg13g2_inv_1 _09357_ (.Y(_02032_),
    .A(net4477));
 sg13g2_inv_1 _09358_ (.Y(_02033_),
    .A(net4441));
 sg13g2_inv_1 _09359_ (.Y(_02034_),
    .A(net4867));
 sg13g2_inv_2 _09360_ (.Y(_02035_),
    .A(net4878));
 sg13g2_inv_2 _09361_ (.Y(_02036_),
    .A(net4564));
 sg13g2_inv_4 _09362_ (.A(net4649),
    .Y(_02037_));
 sg13g2_inv_1 _09363_ (.Y(_02038_),
    .A(net5266));
 sg13g2_inv_1 _09364_ (.Y(_02039_),
    .A(net4341));
 sg13g2_inv_1 _09365_ (.Y(_02040_),
    .A(net3627));
 sg13g2_inv_1 _09366_ (.Y(_02041_),
    .A(net3749));
 sg13g2_inv_2 _09367_ (.Y(_02042_),
    .A(net10));
 sg13g2_inv_1 _09368_ (.Y(_02043_),
    .A(net4003));
 sg13g2_inv_1 _09369_ (.Y(_02044_),
    .A(net3952));
 sg13g2_inv_1 _09370_ (.Y(_02045_),
    .A(net4350));
 sg13g2_inv_1 _09371_ (.Y(_02046_),
    .A(net3380));
 sg13g2_inv_1 _09372_ (.Y(_02047_),
    .A(net2588));
 sg13g2_inv_1 _09373_ (.Y(_02048_),
    .A(net2589));
 sg13g2_inv_1 _09374_ (.Y(_02049_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ));
 sg13g2_inv_1 _09375_ (.Y(_02050_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ));
 sg13g2_inv_1 _09376_ (.Y(_02051_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[6] ));
 sg13g2_inv_1 _09377_ (.Y(_02052_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[7] ));
 sg13g2_inv_1 _09378_ (.Y(_02053_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[8] ));
 sg13g2_inv_1 _09379_ (.Y(_02054_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[9] ));
 sg13g2_inv_1 _09380_ (.Y(_02055_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[10] ));
 sg13g2_inv_1 _09381_ (.Y(_02056_),
    .A(net5380));
 sg13g2_inv_1 _09382_ (.Y(_02057_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[12] ));
 sg13g2_inv_1 _09383_ (.Y(_02058_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[13] ));
 sg13g2_inv_1 _09384_ (.Y(_02059_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[14] ));
 sg13g2_inv_1 _09385_ (.Y(_02060_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[15] ));
 sg13g2_inv_1 _09386_ (.Y(_02061_),
    .A(\i_tinyqv.cpu.i_core.mepc[0] ));
 sg13g2_inv_1 _09387_ (.Y(_02062_),
    .A(net4294));
 sg13g2_inv_1 _09388_ (.Y(_02063_),
    .A(net3724));
 sg13g2_inv_1 _09389_ (.Y(_02064_),
    .A(net3848));
 sg13g2_inv_1 _09390_ (.Y(_02065_),
    .A(\i_latch_mem.data_out[12] ));
 sg13g2_inv_1 _09391_ (.Y(_02066_),
    .A(\i_latch_mem.data_out[20] ));
 sg13g2_inv_1 _09392_ (.Y(_02067_),
    .A(net3641));
 sg13g2_inv_1 _09393_ (.Y(_02068_),
    .A(net2476));
 sg13g2_inv_1 _09394_ (.Y(_02069_),
    .A(\i_latch_mem.data_out[1] ));
 sg13g2_inv_1 _09395_ (.Y(_02070_),
    .A(net3978));
 sg13g2_inv_1 _09396_ (.Y(_02071_),
    .A(net4103));
 sg13g2_inv_1 _09397_ (.Y(_02072_),
    .A(net3878));
 sg13g2_inv_1 _09398_ (.Y(_02073_),
    .A(\i_latch_mem.data_out[25] ));
 sg13g2_inv_1 _09399_ (.Y(_02074_),
    .A(net3623));
 sg13g2_inv_1 _09400_ (.Y(_02075_),
    .A(net4124));
 sg13g2_inv_1 _09401_ (.Y(_02076_),
    .A(net4277));
 sg13g2_inv_1 _09402_ (.Y(_02077_),
    .A(net3740));
 sg13g2_inv_1 _09403_ (.Y(_02078_),
    .A(net3980));
 sg13g2_inv_1 _09404_ (.Y(_02079_),
    .A(\i_latch_mem.data_out[26] ));
 sg13g2_inv_1 _09405_ (.Y(_02080_),
    .A(net3662));
 sg13g2_inv_1 _09406_ (.Y(_02081_),
    .A(net4623));
 sg13g2_inv_1 _09407_ (.Y(_02082_),
    .A(net3823));
 sg13g2_inv_1 _09408_ (.Y(_02083_),
    .A(net3880));
 sg13g2_inv_1 _09409_ (.Y(_02084_),
    .A(\i_latch_mem.data_out[27] ));
 sg13g2_inv_1 _09410_ (.Y(_02085_),
    .A(net3634));
 sg13g2_inv_1 _09411_ (.Y(_02086_),
    .A(\i_latch_mem.data_out[31] ));
 sg13g2_inv_1 _09412_ (.Y(_02087_),
    .A(net4151));
 sg13g2_inv_1 _09413_ (.Y(_02088_),
    .A(net3609));
 sg13g2_inv_1 _16063__2 (.Y(net2722),
    .A(clknet_leaf_65_clk));
 sg13g2_nand2_2 _09415_ (.Y(_02089_),
    .A(\i_tinyqv.cpu.data_write_n[1] ),
    .B(\i_tinyqv.cpu.data_write_n[0] ));
 sg13g2_and2_1 _09416_ (.A(net2471),
    .B(_02089_),
    .X(_02090_));
 sg13g2_nand2_1 _09417_ (.Y(_02091_),
    .A(\addr[0] ),
    .B(\i_latch_mem.cycle[0] ));
 sg13g2_xor2_1 _09418_ (.B(\addr[1] ),
    .A(\i_latch_mem.cycle[1] ),
    .X(_02092_));
 sg13g2_nor2b_1 _09419_ (.A(_02091_),
    .B_N(_02092_),
    .Y(_02093_));
 sg13g2_a21o_2 _09420_ (.A2(\addr[1] ),
    .A1(\i_latch_mem.cycle[1] ),
    .B1(_02093_),
    .X(_02094_));
 sg13g2_nand2_2 _09421_ (.Y(_02095_),
    .A(\addr[2] ),
    .B(\addr[3] ));
 sg13g2_nand2b_2 _09422_ (.Y(_02096_),
    .B(_02094_),
    .A_N(_02095_));
 sg13g2_a21o_1 _09423_ (.A2(_02094_),
    .A1(\addr[2] ),
    .B1(net2466),
    .X(_02097_));
 sg13g2_and2_1 _09424_ (.A(_02096_),
    .B(_02097_),
    .X(_02098_));
 sg13g2_xnor2_1 _09425_ (.Y(_02099_),
    .A(_02013_),
    .B(_02094_));
 sg13g2_nor2_2 _09426_ (.A(_02098_),
    .B(_02099_),
    .Y(_02100_));
 sg13g2_xor2_1 _09427_ (.B(\i_latch_mem.cycle[0] ),
    .A(\addr[0] ),
    .X(_02101_));
 sg13g2_xnor2_1 _09428_ (.Y(_02102_),
    .A(\addr[0] ),
    .B(net2465));
 sg13g2_nand2_2 _09429_ (.Y(_02103_),
    .A(_02092_),
    .B(_02101_));
 sg13g2_nand3_1 _09430_ (.B(_02100_),
    .C(_02101_),
    .A(_02092_),
    .Y(_02104_));
 sg13g2_xnor2_1 _09431_ (.Y(_02105_),
    .A(_02014_),
    .B(_02096_));
 sg13g2_xnor2_1 _09432_ (.Y(_02106_),
    .A(\addr[4] ),
    .B(_02096_));
 sg13g2_nor2_2 _09433_ (.A(_02104_),
    .B(net2140),
    .Y(_02107_));
 sg13g2_nand2_1 _09434_ (.Y(_02108_),
    .A(net2329),
    .B(net1993));
 sg13g2_nor2b_1 _09435_ (.A(\i_latch_mem.cycle[1] ),
    .B_N(net2465),
    .Y(_02109_));
 sg13g2_and2_1 _09436_ (.A(\i_latch_mem.cycle[1] ),
    .B(net2465),
    .X(_02110_));
 sg13g2_nand2_2 _09437_ (.Y(_02111_),
    .A(net5024),
    .B(net2465));
 sg13g2_nor2b_2 _09438_ (.A(net2465),
    .B_N(\i_latch_mem.cycle[1] ),
    .Y(_02112_));
 sg13g2_nor2_1 _09439_ (.A(\i_latch_mem.cycle[1] ),
    .B(net2465),
    .Y(_02113_));
 sg13g2_a22oi_1 _09440_ (.Y(_02114_),
    .B1(net2397),
    .B2(\data_to_write[23] ),
    .A2(net2403),
    .A1(\data_to_write[15] ));
 sg13g2_o21ai_1 _09441_ (.B1(_02114_),
    .Y(_02115_),
    .A1(_01812_),
    .A2(net2399));
 sg13g2_a21oi_2 _09442_ (.B1(_02115_),
    .Y(_02116_),
    .A2(net2393),
    .A1(net2551));
 sg13g2_nand2_1 _09443_ (.Y(_02117_),
    .A(net3526),
    .B(net1919));
 sg13g2_o21ai_1 _09444_ (.B1(_02117_),
    .Y(_01639_),
    .A1(net1919),
    .A2(net2182));
 sg13g2_a22oi_1 _09445_ (.Y(_02118_),
    .B1(net2398),
    .B2(\data_to_write[22] ),
    .A2(net2401),
    .A1(\data_to_write[30] ));
 sg13g2_a22oi_1 _09446_ (.Y(_02119_),
    .B1(net2394),
    .B2(net2552),
    .A2(net2403),
    .A1(\data_to_write[14] ));
 sg13g2_and2_1 _09447_ (.A(_02118_),
    .B(_02119_),
    .X(_02120_));
 sg13g2_nand2_1 _09448_ (.Y(_02121_),
    .A(net3498),
    .B(net1920));
 sg13g2_o21ai_1 _09449_ (.B1(_02121_),
    .Y(_01638_),
    .A1(net1920),
    .A2(net2276));
 sg13g2_a22oi_1 _09450_ (.Y(_02122_),
    .B1(net2398),
    .B2(\data_to_write[21] ),
    .A2(net2401),
    .A1(\data_to_write[29] ));
 sg13g2_a22oi_1 _09451_ (.Y(_02123_),
    .B1(net2393),
    .B2(net2553),
    .A2(net2403),
    .A1(\data_to_write[13] ));
 sg13g2_and2_1 _09452_ (.A(_02122_),
    .B(_02123_),
    .X(_02124_));
 sg13g2_nand2_1 _09453_ (.Y(_02125_),
    .A(net3455),
    .B(net1919));
 sg13g2_o21ai_1 _09454_ (.B1(_02125_),
    .Y(_01637_),
    .A1(net1920),
    .A2(net2270));
 sg13g2_a22oi_1 _09455_ (.Y(_02126_),
    .B1(net2393),
    .B2(net2554),
    .A2(net2401),
    .A1(\data_to_write[28] ));
 sg13g2_a22oi_1 _09456_ (.Y(_02127_),
    .B1(net2398),
    .B2(\data_to_write[20] ),
    .A2(net2403),
    .A1(\data_to_write[12] ));
 sg13g2_and2_1 _09457_ (.A(_02126_),
    .B(_02127_),
    .X(_02128_));
 sg13g2_nand2_1 _09458_ (.Y(_02129_),
    .A(net3531),
    .B(net1920));
 sg13g2_o21ai_1 _09459_ (.B1(_02129_),
    .Y(_01636_),
    .A1(net1920),
    .A2(net2266));
 sg13g2_a22oi_1 _09460_ (.Y(_02130_),
    .B1(net2401),
    .B2(\data_to_write[27] ),
    .A2(net2403),
    .A1(\data_to_write[11] ));
 sg13g2_a22oi_1 _09461_ (.Y(_02131_),
    .B1(net2393),
    .B2(net2555),
    .A2(net2398),
    .A1(\data_to_write[19] ));
 sg13g2_and2_1 _09462_ (.A(_02130_),
    .B(_02131_),
    .X(_02132_));
 sg13g2_nand2_1 _09463_ (.Y(_02133_),
    .A(net3580),
    .B(net1919));
 sg13g2_o21ai_1 _09464_ (.B1(_02133_),
    .Y(_01635_),
    .A1(net1919),
    .A2(net2261));
 sg13g2_a22oi_1 _09465_ (.Y(_02134_),
    .B1(net2394),
    .B2(net2556),
    .A2(net2401),
    .A1(\data_to_write[26] ));
 sg13g2_a22oi_1 _09466_ (.Y(_02135_),
    .B1(net2398),
    .B2(\data_to_write[18] ),
    .A2(net2403),
    .A1(\data_to_write[10] ));
 sg13g2_and2_1 _09467_ (.A(_02134_),
    .B(_02135_),
    .X(_02136_));
 sg13g2_nand2_1 _09468_ (.Y(_02137_),
    .A(net3432),
    .B(net1919));
 sg13g2_o21ai_1 _09469_ (.B1(_02137_),
    .Y(_01634_),
    .A1(_02108_),
    .A2(net2255));
 sg13g2_a22oi_1 _09470_ (.Y(_02138_),
    .B1(net2394),
    .B2(net2557),
    .A2(net2401),
    .A1(\data_to_write[25] ));
 sg13g2_a22oi_1 _09471_ (.Y(_02139_),
    .B1(net2398),
    .B2(\data_to_write[17] ),
    .A2(net2404),
    .A1(\data_to_write[9] ));
 sg13g2_and2_1 _09472_ (.A(_02138_),
    .B(_02139_),
    .X(_02140_));
 sg13g2_nand2_1 _09473_ (.Y(_02141_),
    .A(net3456),
    .B(net1919));
 sg13g2_o21ai_1 _09474_ (.B1(_02141_),
    .Y(_01633_),
    .A1(net1919),
    .A2(net2250));
 sg13g2_a22oi_1 _09475_ (.Y(_02142_),
    .B1(net2401),
    .B2(\data_to_write[24] ),
    .A2(net2404),
    .A1(net2549));
 sg13g2_a22oi_1 _09476_ (.Y(_02143_),
    .B1(net2394),
    .B2(net2559),
    .A2(net2398),
    .A1(\data_to_write[16] ));
 sg13g2_and2_1 _09477_ (.A(_02142_),
    .B(_02143_),
    .X(_02144_));
 sg13g2_nand2_1 _09478_ (.Y(_02145_),
    .A(net3548),
    .B(net1920));
 sg13g2_o21ai_1 _09479_ (.B1(_02145_),
    .Y(_01632_),
    .A1(net1920),
    .A2(net2246));
 sg13g2_nand2_2 _09480_ (.Y(_02146_),
    .A(net2466),
    .B(_02099_));
 sg13g2_nand2b_2 _09481_ (.Y(_02147_),
    .B(_02101_),
    .A_N(_02092_));
 sg13g2_nor3_1 _09482_ (.A(net2141),
    .B(_02146_),
    .C(_02147_),
    .Y(_02148_));
 sg13g2_and2_1 _09483_ (.A(net2327),
    .B(net2101),
    .X(_02149_));
 sg13g2_nor2_1 _09484_ (.A(net4070),
    .B(net2044),
    .Y(_02150_));
 sg13g2_a21oi_1 _09485_ (.A1(net2180),
    .A2(net2044),
    .Y(_01631_),
    .B1(_02150_));
 sg13g2_nor2_1 _09486_ (.A(net4157),
    .B(net2045),
    .Y(_02151_));
 sg13g2_a21oi_1 _09487_ (.A1(net2275),
    .A2(net2045),
    .Y(_01630_),
    .B1(_02151_));
 sg13g2_nor2_1 _09488_ (.A(net3872),
    .B(net2044),
    .Y(_02152_));
 sg13g2_a21oi_1 _09489_ (.A1(net2272),
    .A2(net2044),
    .Y(_01629_),
    .B1(_02152_));
 sg13g2_nor2_1 _09490_ (.A(net3822),
    .B(net2044),
    .Y(_02153_));
 sg13g2_a21oi_1 _09491_ (.A1(net2263),
    .A2(net2044),
    .Y(_01628_),
    .B1(_02153_));
 sg13g2_nor2_1 _09492_ (.A(net4256),
    .B(net2046),
    .Y(_02154_));
 sg13g2_a21oi_1 _09493_ (.A1(net2260),
    .A2(net2046),
    .Y(_01627_),
    .B1(_02154_));
 sg13g2_nor2_1 _09494_ (.A(net3856),
    .B(net2044),
    .Y(_02155_));
 sg13g2_a21oi_1 _09495_ (.A1(net2253),
    .A2(net2044),
    .Y(_01626_),
    .B1(_02155_));
 sg13g2_nor2_1 _09496_ (.A(net4149),
    .B(net2046),
    .Y(_02156_));
 sg13g2_a21oi_1 _09497_ (.A1(net2251),
    .A2(net2046),
    .Y(_01625_),
    .B1(_02156_));
 sg13g2_nor2_1 _09498_ (.A(net4362),
    .B(net2045),
    .Y(_02157_));
 sg13g2_a21oi_1 _09499_ (.A1(net2243),
    .A2(net2045),
    .Y(_01624_),
    .B1(_02157_));
 sg13g2_nor3_2 _09500_ (.A(_02103_),
    .B(net2141),
    .C(_02146_),
    .Y(_02158_));
 sg13g2_and2_1 _09501_ (.A(net2327),
    .B(net2100),
    .X(_02159_));
 sg13g2_nor2_1 _09502_ (.A(net3921),
    .B(net2043),
    .Y(_02160_));
 sg13g2_a21oi_1 _09503_ (.A1(net2179),
    .A2(net2043),
    .Y(_01623_),
    .B1(_02160_));
 sg13g2_nor2_1 _09504_ (.A(net3784),
    .B(net2043),
    .Y(_02161_));
 sg13g2_a21oi_1 _09505_ (.A1(net2275),
    .A2(net2043),
    .Y(_01622_),
    .B1(_02161_));
 sg13g2_nor2_1 _09506_ (.A(net3718),
    .B(net2042),
    .Y(_02162_));
 sg13g2_a21oi_1 _09507_ (.A1(net2269),
    .A2(net2042),
    .Y(_01621_),
    .B1(_02162_));
 sg13g2_nor2_1 _09508_ (.A(net4001),
    .B(net2042),
    .Y(_02163_));
 sg13g2_a21oi_1 _09509_ (.A1(net2264),
    .A2(net2042),
    .Y(_01620_),
    .B1(_02163_));
 sg13g2_nor2_1 _09510_ (.A(net3827),
    .B(net2042),
    .Y(_02164_));
 sg13g2_a21oi_1 _09511_ (.A1(net2258),
    .A2(net2042),
    .Y(_01619_),
    .B1(_02164_));
 sg13g2_nor2_1 _09512_ (.A(net4054),
    .B(net2043),
    .Y(_02165_));
 sg13g2_a21oi_1 _09513_ (.A1(net2253),
    .A2(net2043),
    .Y(_01618_),
    .B1(_02165_));
 sg13g2_nor2_1 _09514_ (.A(net3883),
    .B(net2042),
    .Y(_02166_));
 sg13g2_a21oi_1 _09515_ (.A1(net2248),
    .A2(net2042),
    .Y(_01617_),
    .B1(_02166_));
 sg13g2_nor2_1 _09516_ (.A(net3797),
    .B(net2043),
    .Y(_02167_));
 sg13g2_a21oi_1 _09517_ (.A1(net2243),
    .A2(net2043),
    .Y(_01616_),
    .B1(_02167_));
 sg13g2_nor2_1 _09518_ (.A(_02104_),
    .B(net2139),
    .Y(_02168_));
 sg13g2_nand2_2 _09519_ (.Y(_02169_),
    .A(net2329),
    .B(net1992));
 sg13g2_nand2_1 _09520_ (.Y(_02170_),
    .A(net3672),
    .B(net1917));
 sg13g2_o21ai_1 _09521_ (.B1(_02170_),
    .Y(_01615_),
    .A1(net2183),
    .A2(net1917));
 sg13g2_nand2_1 _09522_ (.Y(_02171_),
    .A(net3657),
    .B(net1917));
 sg13g2_o21ai_1 _09523_ (.B1(_02171_),
    .Y(_01614_),
    .A1(net2277),
    .A2(net1917));
 sg13g2_nand2_1 _09524_ (.Y(_02172_),
    .A(net3457),
    .B(net1917));
 sg13g2_o21ai_1 _09525_ (.B1(_02172_),
    .Y(_01613_),
    .A1(net2271),
    .A2(net1917));
 sg13g2_nand2_1 _09526_ (.Y(_02173_),
    .A(net3537),
    .B(net1917));
 sg13g2_o21ai_1 _09527_ (.B1(_02173_),
    .Y(_01612_),
    .A1(net2266),
    .A2(net1917));
 sg13g2_nand2_1 _09528_ (.Y(_02174_),
    .A(net3538),
    .B(net1918));
 sg13g2_o21ai_1 _09529_ (.B1(_02174_),
    .Y(_01611_),
    .A1(net2261),
    .A2(net1918));
 sg13g2_nand2_1 _09530_ (.Y(_02175_),
    .A(net3611),
    .B(net1918));
 sg13g2_o21ai_1 _09531_ (.B1(_02175_),
    .Y(_01610_),
    .A1(net2255),
    .A2(net1918));
 sg13g2_nand2_1 _09532_ (.Y(_02176_),
    .A(net3563),
    .B(net1918));
 sg13g2_o21ai_1 _09533_ (.B1(_02176_),
    .Y(_01609_),
    .A1(net2250),
    .A2(net1918));
 sg13g2_nand2_1 _09534_ (.Y(_02177_),
    .A(net3586),
    .B(net1918));
 sg13g2_o21ai_1 _09535_ (.B1(_02177_),
    .Y(_01608_),
    .A1(net2246),
    .A2(net1918));
 sg13g2_nand2b_2 _09536_ (.Y(_02178_),
    .B(_02099_),
    .A_N(net2466));
 sg13g2_xnor2_1 _09537_ (.Y(_02179_),
    .A(_02091_),
    .B(_02092_));
 sg13g2_or2_1 _09538_ (.X(_02180_),
    .B(_02179_),
    .A(_02101_));
 sg13g2_inv_2 _09539_ (.Y(_02181_),
    .A(_02180_));
 sg13g2_nor3_1 _09540_ (.A(net2138),
    .B(_02178_),
    .C(_02180_),
    .Y(_02182_));
 sg13g2_nand2_2 _09541_ (.Y(_02183_),
    .A(net2328),
    .B(net2099));
 sg13g2_nand2_1 _09542_ (.Y(_02184_),
    .A(net3533),
    .B(net2041));
 sg13g2_o21ai_1 _09543_ (.B1(_02184_),
    .Y(_01607_),
    .A1(net2181),
    .A2(net2041));
 sg13g2_nand2_1 _09544_ (.Y(_02185_),
    .A(net3638),
    .B(net2040));
 sg13g2_o21ai_1 _09545_ (.B1(_02185_),
    .Y(_01606_),
    .A1(net2274),
    .A2(net2040));
 sg13g2_nand2_1 _09546_ (.Y(_02186_),
    .A(net3421),
    .B(net2041));
 sg13g2_o21ai_1 _09547_ (.B1(_02186_),
    .Y(_01605_),
    .A1(net2268),
    .A2(net2041));
 sg13g2_nand2_1 _09548_ (.Y(_02187_),
    .A(net3508),
    .B(net2041));
 sg13g2_o21ai_1 _09549_ (.B1(_02187_),
    .Y(_01604_),
    .A1(net2264),
    .A2(net2041));
 sg13g2_nand2_1 _09550_ (.Y(_02188_),
    .A(net3903),
    .B(net2041));
 sg13g2_o21ai_1 _09551_ (.B1(_02188_),
    .Y(_01603_),
    .A1(net2258),
    .A2(net2041));
 sg13g2_nand2_1 _09552_ (.Y(_02189_),
    .A(net3463),
    .B(net2040));
 sg13g2_o21ai_1 _09553_ (.B1(_02189_),
    .Y(_01602_),
    .A1(net2254),
    .A2(net2040));
 sg13g2_nand2_1 _09554_ (.Y(_02190_),
    .A(net3596),
    .B(net2040));
 sg13g2_o21ai_1 _09555_ (.B1(_02190_),
    .Y(_01601_),
    .A1(net2248),
    .A2(net2040));
 sg13g2_nand2_1 _09556_ (.Y(_02191_),
    .A(net3520),
    .B(net2040));
 sg13g2_o21ai_1 _09557_ (.B1(_02191_),
    .Y(_01600_),
    .A1(net2245),
    .A2(net2040));
 sg13g2_nor3_2 _09558_ (.A(net2138),
    .B(_02147_),
    .C(_02178_),
    .Y(_02192_));
 sg13g2_nand2_1 _09559_ (.Y(_02193_),
    .A(net2328),
    .B(net2098));
 sg13g2_nand2_1 _09560_ (.Y(_02194_),
    .A(net3934),
    .B(net2038));
 sg13g2_o21ai_1 _09561_ (.B1(_02194_),
    .Y(_01599_),
    .A1(net2181),
    .A2(net2038));
 sg13g2_nand2_1 _09562_ (.Y(_02195_),
    .A(net3753),
    .B(net2039));
 sg13g2_o21ai_1 _09563_ (.B1(_02195_),
    .Y(_01598_),
    .A1(net2274),
    .A2(net2039));
 sg13g2_nand2_1 _09564_ (.Y(_02196_),
    .A(net3512),
    .B(net2038));
 sg13g2_o21ai_1 _09565_ (.B1(_02196_),
    .Y(_01597_),
    .A1(net2268),
    .A2(net2038));
 sg13g2_nand2_1 _09566_ (.Y(_02197_),
    .A(net3601),
    .B(net2039));
 sg13g2_o21ai_1 _09567_ (.B1(_02197_),
    .Y(_01596_),
    .A1(net2264),
    .A2(net2039));
 sg13g2_nand2_1 _09568_ (.Y(_02198_),
    .A(net3582),
    .B(net2039));
 sg13g2_o21ai_1 _09569_ (.B1(_02198_),
    .Y(_01595_),
    .A1(net2258),
    .A2(net2039));
 sg13g2_nand2_1 _09570_ (.Y(_02199_),
    .A(net3574),
    .B(net2039));
 sg13g2_o21ai_1 _09571_ (.B1(_02199_),
    .Y(_01594_),
    .A1(net2254),
    .A2(_02193_));
 sg13g2_nand2_1 _09572_ (.Y(_02200_),
    .A(net3639),
    .B(net2038));
 sg13g2_o21ai_1 _09573_ (.B1(_02200_),
    .Y(_01593_),
    .A1(net2248),
    .A2(net2038));
 sg13g2_nand2_1 _09574_ (.Y(_02201_),
    .A(net3585),
    .B(net2038));
 sg13g2_o21ai_1 _09575_ (.B1(_02201_),
    .Y(_01592_),
    .A1(net2245),
    .A2(net2038));
 sg13g2_nand2_2 _09576_ (.Y(_02202_),
    .A(_02102_),
    .B(_02179_));
 sg13g2_nor3_1 _09577_ (.A(net2138),
    .B(_02178_),
    .C(_02202_),
    .Y(_02203_));
 sg13g2_nand2_1 _09578_ (.Y(_02204_),
    .A(net2328),
    .B(net2097));
 sg13g2_nand2_1 _09579_ (.Y(_02205_),
    .A(net3705),
    .B(net2036));
 sg13g2_o21ai_1 _09580_ (.B1(_02205_),
    .Y(_01591_),
    .A1(net2181),
    .A2(net2036));
 sg13g2_nand2_1 _09581_ (.Y(_02206_),
    .A(net3576),
    .B(net2036));
 sg13g2_o21ai_1 _09582_ (.B1(_02206_),
    .Y(_01590_),
    .A1(net2274),
    .A2(net2036));
 sg13g2_nand2_1 _09583_ (.Y(_02207_),
    .A(net3792),
    .B(net2037));
 sg13g2_o21ai_1 _09584_ (.B1(_02207_),
    .Y(_01589_),
    .A1(net2268),
    .A2(net2037));
 sg13g2_nand2_1 _09585_ (.Y(_02208_),
    .A(net3447),
    .B(net2037));
 sg13g2_o21ai_1 _09586_ (.B1(_02208_),
    .Y(_01588_),
    .A1(net2264),
    .A2(net2037));
 sg13g2_nand2_1 _09587_ (.Y(_02209_),
    .A(net3737),
    .B(net2037));
 sg13g2_o21ai_1 _09588_ (.B1(_02209_),
    .Y(_01587_),
    .A1(net2258),
    .A2(_02204_));
 sg13g2_nand2_1 _09589_ (.Y(_02210_),
    .A(net3494),
    .B(net2036));
 sg13g2_o21ai_1 _09590_ (.B1(_02210_),
    .Y(_01586_),
    .A1(net2254),
    .A2(net2036));
 sg13g2_nand2_1 _09591_ (.Y(_02211_),
    .A(net3469),
    .B(net2037));
 sg13g2_o21ai_1 _09592_ (.B1(_02211_),
    .Y(_01585_),
    .A1(net2248),
    .A2(net2037));
 sg13g2_nand2_1 _09593_ (.Y(_02212_),
    .A(net3428),
    .B(net2036));
 sg13g2_o21ai_1 _09594_ (.B1(_02212_),
    .Y(_01584_),
    .A1(net2245),
    .A2(net2036));
 sg13g2_nor3_1 _09595_ (.A(_02103_),
    .B(net2138),
    .C(_02178_),
    .Y(_02213_));
 sg13g2_nand2_1 _09596_ (.Y(_02214_),
    .A(net2327),
    .B(net2096));
 sg13g2_nand2_1 _09597_ (.Y(_02215_),
    .A(net3488),
    .B(net2033));
 sg13g2_o21ai_1 _09598_ (.B1(_02215_),
    .Y(_01583_),
    .A1(net2179),
    .A2(net2033));
 sg13g2_nand2_1 _09599_ (.Y(_02216_),
    .A(net3424),
    .B(net2033));
 sg13g2_o21ai_1 _09600_ (.B1(_02216_),
    .Y(_01582_),
    .A1(net2275),
    .A2(net2033));
 sg13g2_nand2_1 _09601_ (.Y(_02217_),
    .A(net3461),
    .B(net2035));
 sg13g2_o21ai_1 _09602_ (.B1(_02217_),
    .Y(_01581_),
    .A1(net2268),
    .A2(net2035));
 sg13g2_nand2_1 _09603_ (.Y(_02218_),
    .A(net3462),
    .B(net2034));
 sg13g2_o21ai_1 _09604_ (.B1(_02218_),
    .Y(_01580_),
    .A1(net2263),
    .A2(net2034));
 sg13g2_nand2_1 _09605_ (.Y(_02219_),
    .A(net3485),
    .B(net2033));
 sg13g2_o21ai_1 _09606_ (.B1(_02219_),
    .Y(_01579_),
    .A1(net2260),
    .A2(net2033));
 sg13g2_nand2_1 _09607_ (.Y(_02220_),
    .A(net3495),
    .B(net2035));
 sg13g2_o21ai_1 _09608_ (.B1(_02220_),
    .Y(_01578_),
    .A1(net2254),
    .A2(net2035));
 sg13g2_nand2_1 _09609_ (.Y(_02221_),
    .A(net3510),
    .B(net2033));
 sg13g2_o21ai_1 _09610_ (.B1(_02221_),
    .Y(_01577_),
    .A1(net2251),
    .A2(net2033));
 sg13g2_nand2_1 _09611_ (.Y(_02222_),
    .A(net3595),
    .B(net2034));
 sg13g2_o21ai_1 _09612_ (.B1(_02222_),
    .Y(_01576_),
    .A1(net2244),
    .A2(net2034));
 sg13g2_nand2b_2 _09613_ (.Y(_02223_),
    .B(_02098_),
    .A_N(_02099_));
 sg13g2_nor3_2 _09614_ (.A(net2139),
    .B(_02180_),
    .C(_02223_),
    .Y(_02224_));
 sg13g2_nand2_2 _09615_ (.Y(_02225_),
    .A(net2329),
    .B(net2032));
 sg13g2_nand2_1 _09616_ (.Y(_02226_),
    .A(net3509),
    .B(net1990));
 sg13g2_o21ai_1 _09617_ (.B1(_02226_),
    .Y(_01575_),
    .A1(net2182),
    .A2(net1991));
 sg13g2_nand2_1 _09618_ (.Y(_02227_),
    .A(net3525),
    .B(net1990));
 sg13g2_o21ai_1 _09619_ (.B1(_02227_),
    .Y(_01574_),
    .A1(net2276),
    .A2(net1990));
 sg13g2_nand2_1 _09620_ (.Y(_02228_),
    .A(net3584),
    .B(net1991));
 sg13g2_o21ai_1 _09621_ (.B1(_02228_),
    .Y(_01573_),
    .A1(net2270),
    .A2(net1990));
 sg13g2_nand2_1 _09622_ (.Y(_02229_),
    .A(net3483),
    .B(net1990));
 sg13g2_o21ai_1 _09623_ (.B1(_02229_),
    .Y(_01572_),
    .A1(net2265),
    .A2(net1990));
 sg13g2_nand2_1 _09624_ (.Y(_02230_),
    .A(net3497),
    .B(net1991));
 sg13g2_o21ai_1 _09625_ (.B1(_02230_),
    .Y(_01571_),
    .A1(net2259),
    .A2(net1991));
 sg13g2_nand2_1 _09626_ (.Y(_02231_),
    .A(net3560),
    .B(net1991));
 sg13g2_o21ai_1 _09627_ (.B1(_02231_),
    .Y(_01570_),
    .A1(net2256),
    .A2(net1991));
 sg13g2_nand2_1 _09628_ (.Y(_02232_),
    .A(net3458),
    .B(net1991));
 sg13g2_o21ai_1 _09629_ (.B1(_02232_),
    .Y(_01569_),
    .A1(net2249),
    .A2(net1991));
 sg13g2_nand2_1 _09630_ (.Y(_02233_),
    .A(net3434),
    .B(net1990));
 sg13g2_o21ai_1 _09631_ (.B1(_02233_),
    .Y(_01568_),
    .A1(net2244),
    .A2(net1990));
 sg13g2_nand2_2 _09632_ (.Y(_02234_),
    .A(_02100_),
    .B(_02181_));
 sg13g2_nor2_2 _09633_ (.A(net2139),
    .B(_02234_),
    .Y(_02235_));
 sg13g2_nand3_1 _09634_ (.B(net2140),
    .C(_02181_),
    .A(_02100_),
    .Y(_02236_));
 sg13g2_nand2_2 _09635_ (.Y(_02237_),
    .A(net2328),
    .B(net1989));
 sg13g2_nand2_1 _09636_ (.Y(_02238_),
    .A(net3435),
    .B(net1915));
 sg13g2_o21ai_1 _09637_ (.B1(_02238_),
    .Y(_01567_),
    .A1(net2181),
    .A2(net1915));
 sg13g2_nand2_1 _09638_ (.Y(_02239_),
    .A(net3418),
    .B(net1916));
 sg13g2_o21ai_1 _09639_ (.B1(_02239_),
    .Y(_01566_),
    .A1(net2274),
    .A2(net1916));
 sg13g2_nand2_1 _09640_ (.Y(_02240_),
    .A(net3536),
    .B(net1916));
 sg13g2_o21ai_1 _09641_ (.B1(_02240_),
    .Y(_01565_),
    .A1(net2268),
    .A2(net1916));
 sg13g2_nand2_1 _09642_ (.Y(_02241_),
    .A(net3474),
    .B(net1915));
 sg13g2_o21ai_1 _09643_ (.B1(_02241_),
    .Y(_01564_),
    .A1(net2264),
    .A2(net1915));
 sg13g2_nand2_1 _09644_ (.Y(_02242_),
    .A(net3518),
    .B(net1915));
 sg13g2_o21ai_1 _09645_ (.B1(_02242_),
    .Y(_01563_),
    .A1(net2259),
    .A2(net1915));
 sg13g2_nand2_1 _09646_ (.Y(_02243_),
    .A(net3492),
    .B(net1916));
 sg13g2_o21ai_1 _09647_ (.B1(_02243_),
    .Y(_01562_),
    .A1(net2254),
    .A2(net1916));
 sg13g2_nand2_1 _09648_ (.Y(_02244_),
    .A(net3496),
    .B(net1916));
 sg13g2_o21ai_1 _09649_ (.B1(_02244_),
    .Y(_01561_),
    .A1(net2249),
    .A2(net1916));
 sg13g2_nand2_1 _09650_ (.Y(_02245_),
    .A(net3493),
    .B(net1915));
 sg13g2_o21ai_1 _09651_ (.B1(_02245_),
    .Y(_01560_),
    .A1(net2245),
    .A2(net1915));
 sg13g2_nor3_1 _09652_ (.A(net2139),
    .B(_02202_),
    .C(_02223_),
    .Y(_02246_));
 sg13g2_nand2_1 _09653_ (.Y(_02247_),
    .A(net2329),
    .B(net2031));
 sg13g2_nand2_1 _09654_ (.Y(_02248_),
    .A(net3579),
    .B(net1988));
 sg13g2_o21ai_1 _09655_ (.B1(_02248_),
    .Y(_01559_),
    .A1(net2182),
    .A2(net1988));
 sg13g2_nand2_1 _09656_ (.Y(_02249_),
    .A(net3506),
    .B(net1988));
 sg13g2_o21ai_1 _09657_ (.B1(_02249_),
    .Y(_01558_),
    .A1(net2276),
    .A2(net1988));
 sg13g2_nand2_1 _09658_ (.Y(_02250_),
    .A(net3517),
    .B(net1987));
 sg13g2_o21ai_1 _09659_ (.B1(_02250_),
    .Y(_01557_),
    .A1(net2270),
    .A2(_02247_));
 sg13g2_nand2_1 _09660_ (.Y(_02251_),
    .A(net3640),
    .B(net1987));
 sg13g2_o21ai_1 _09661_ (.B1(_02251_),
    .Y(_01556_),
    .A1(net2265),
    .A2(net1988));
 sg13g2_nand2_1 _09662_ (.Y(_02252_),
    .A(net3738),
    .B(net1987));
 sg13g2_o21ai_1 _09663_ (.B1(_02252_),
    .Y(_01555_),
    .A1(net2262),
    .A2(net1987));
 sg13g2_nand2_1 _09664_ (.Y(_02253_),
    .A(net3464),
    .B(net1988));
 sg13g2_o21ai_1 _09665_ (.B1(_02253_),
    .Y(_01554_),
    .A1(net2255),
    .A2(net1988));
 sg13g2_nand2_1 _09666_ (.Y(_02254_),
    .A(net3739),
    .B(net1987));
 sg13g2_o21ai_1 _09667_ (.B1(_02254_),
    .Y(_01553_),
    .A1(net2250),
    .A2(net1987));
 sg13g2_nand2_1 _09668_ (.Y(_02255_),
    .A(net3597),
    .B(net1987));
 sg13g2_o21ai_1 _09669_ (.B1(_02255_),
    .Y(_01552_),
    .A1(net2244),
    .A2(net1987));
 sg13g2_nor3_2 _09670_ (.A(_02103_),
    .B(net2139),
    .C(_02223_),
    .Y(_02256_));
 sg13g2_nand2_2 _09671_ (.Y(_02257_),
    .A(net2329),
    .B(net2030));
 sg13g2_nand2_1 _09672_ (.Y(_02258_),
    .A(net3821),
    .B(net1986));
 sg13g2_o21ai_1 _09673_ (.B1(_02258_),
    .Y(_01551_),
    .A1(net2180),
    .A2(net1986));
 sg13g2_nand2_1 _09674_ (.Y(_02259_),
    .A(net3453),
    .B(net1985));
 sg13g2_o21ai_1 _09675_ (.B1(_02259_),
    .Y(_01550_),
    .A1(net2278),
    .A2(net1985));
 sg13g2_nand2_1 _09676_ (.Y(_02260_),
    .A(net3532),
    .B(net1986));
 sg13g2_o21ai_1 _09677_ (.B1(_02260_),
    .Y(_01549_),
    .A1(net2270),
    .A2(net1986));
 sg13g2_nand2_1 _09678_ (.Y(_02261_),
    .A(net3593),
    .B(net1985));
 sg13g2_o21ai_1 _09679_ (.B1(_02261_),
    .Y(_01548_),
    .A1(net2265),
    .A2(net1985));
 sg13g2_nand2_1 _09680_ (.Y(_02262_),
    .A(net3587),
    .B(net1986));
 sg13g2_o21ai_1 _09681_ (.B1(_02262_),
    .Y(_01547_),
    .A1(net2261),
    .A2(net1986));
 sg13g2_nand2_1 _09682_ (.Y(_02263_),
    .A(net3468),
    .B(net1986));
 sg13g2_o21ai_1 _09683_ (.B1(_02263_),
    .Y(_01546_),
    .A1(net2255),
    .A2(net1986));
 sg13g2_nand2_1 _09684_ (.Y(_02264_),
    .A(net3572),
    .B(net1985));
 sg13g2_o21ai_1 _09685_ (.B1(_02264_),
    .Y(_01545_),
    .A1(net2249),
    .A2(net1985));
 sg13g2_nand2_1 _09686_ (.Y(_02265_),
    .A(net3422),
    .B(net1985));
 sg13g2_o21ai_1 _09687_ (.B1(_02265_),
    .Y(_01544_),
    .A1(net2244),
    .A2(net1985));
 sg13g2_nand2b_2 _09688_ (.Y(_02266_),
    .B(_02181_),
    .A_N(_02146_));
 sg13g2_nor2_2 _09689_ (.A(net2138),
    .B(_02266_),
    .Y(_02267_));
 sg13g2_and2_1 _09690_ (.A(net2328),
    .B(net2029),
    .X(_02268_));
 sg13g2_nor2_1 _09691_ (.A(net3681),
    .B(net1984),
    .Y(_02269_));
 sg13g2_a21oi_1 _09692_ (.A1(net2181),
    .A2(net1984),
    .Y(_01543_),
    .B1(_02269_));
 sg13g2_nor2_1 _09693_ (.A(net3760),
    .B(net1983),
    .Y(_02270_));
 sg13g2_a21oi_1 _09694_ (.A1(net2274),
    .A2(net1983),
    .Y(_01542_),
    .B1(_02270_));
 sg13g2_nor2_1 _09695_ (.A(net3940),
    .B(net1984),
    .Y(_02271_));
 sg13g2_a21oi_1 _09696_ (.A1(net2268),
    .A2(net1984),
    .Y(_01541_),
    .B1(_02271_));
 sg13g2_nor2_1 _09697_ (.A(net3788),
    .B(net1984),
    .Y(_02272_));
 sg13g2_a21oi_1 _09698_ (.A1(net2264),
    .A2(_02268_),
    .Y(_01540_),
    .B1(_02272_));
 sg13g2_nor2_1 _09699_ (.A(net3696),
    .B(net1983),
    .Y(_02273_));
 sg13g2_a21oi_1 _09700_ (.A1(net2258),
    .A2(net1983),
    .Y(_01539_),
    .B1(_02273_));
 sg13g2_nor2_1 _09701_ (.A(net4002),
    .B(net1983),
    .Y(_02274_));
 sg13g2_a21oi_1 _09702_ (.A1(net2254),
    .A2(net1983),
    .Y(_01538_),
    .B1(_02274_));
 sg13g2_nor2_1 _09703_ (.A(net3869),
    .B(net1984),
    .Y(_02275_));
 sg13g2_a21oi_1 _09704_ (.A1(net2248),
    .A2(net1984),
    .Y(_01537_),
    .B1(_02275_));
 sg13g2_nor2_1 _09705_ (.A(net3863),
    .B(net1983),
    .Y(_02276_));
 sg13g2_a21oi_1 _09706_ (.A1(net2245),
    .A2(net1983),
    .Y(_01536_),
    .B1(_02276_));
 sg13g2_nor3_1 _09707_ (.A(net2138),
    .B(_02146_),
    .C(_02147_),
    .Y(_02277_));
 sg13g2_and2_1 _09708_ (.A(net2328),
    .B(net2095),
    .X(_02278_));
 sg13g2_nor2_1 _09709_ (.A(net3698),
    .B(net2027),
    .Y(_02279_));
 sg13g2_a21oi_1 _09710_ (.A1(net2179),
    .A2(net2027),
    .Y(_01535_),
    .B1(_02279_));
 sg13g2_nor2_1 _09711_ (.A(net4075),
    .B(net2027),
    .Y(_02280_));
 sg13g2_a21oi_1 _09712_ (.A1(net2274),
    .A2(_02278_),
    .Y(_01534_),
    .B1(_02280_));
 sg13g2_nor2_1 _09713_ (.A(net3702),
    .B(net2027),
    .Y(_02281_));
 sg13g2_a21oi_1 _09714_ (.A1(net2269),
    .A2(net2027),
    .Y(_01533_),
    .B1(_02281_));
 sg13g2_nor2_1 _09715_ (.A(net3691),
    .B(net2028),
    .Y(_02282_));
 sg13g2_a21oi_1 _09716_ (.A1(net2264),
    .A2(net2028),
    .Y(_01532_),
    .B1(_02282_));
 sg13g2_nor2_1 _09717_ (.A(net3700),
    .B(net2027),
    .Y(_02283_));
 sg13g2_a21oi_1 _09718_ (.A1(net2258),
    .A2(net2028),
    .Y(_01531_),
    .B1(_02283_));
 sg13g2_nor2_1 _09719_ (.A(net3658),
    .B(net2027),
    .Y(_02284_));
 sg13g2_a21oi_1 _09720_ (.A1(net2253),
    .A2(net2027),
    .Y(_01530_),
    .B1(_02284_));
 sg13g2_nor2_1 _09721_ (.A(net3873),
    .B(net2028),
    .Y(_02285_));
 sg13g2_a21oi_1 _09722_ (.A1(net2248),
    .A2(net2028),
    .Y(_01529_),
    .B1(_02285_));
 sg13g2_nor2_1 _09723_ (.A(net3699),
    .B(net2028),
    .Y(_02286_));
 sg13g2_a21oi_1 _09724_ (.A1(net2245),
    .A2(net2028),
    .Y(_01528_),
    .B1(_02286_));
 sg13g2_or2_1 _09725_ (.X(_02287_),
    .B(_02202_),
    .A(_02146_));
 sg13g2_nor2_2 _09726_ (.A(net2138),
    .B(_02287_),
    .Y(_02288_));
 sg13g2_and2_1 _09727_ (.A(net2331),
    .B(net2026),
    .X(_02289_));
 sg13g2_nor2_1 _09728_ (.A(net4150),
    .B(net1982),
    .Y(_02290_));
 sg13g2_a21oi_1 _09729_ (.A1(net2179),
    .A2(net1982),
    .Y(_01527_),
    .B1(_02290_));
 sg13g2_nor2_1 _09730_ (.A(net4220),
    .B(net1981),
    .Y(_02291_));
 sg13g2_a21oi_1 _09731_ (.A1(net2275),
    .A2(net1982),
    .Y(_01526_),
    .B1(_02291_));
 sg13g2_nor2_1 _09732_ (.A(net3701),
    .B(net1981),
    .Y(_02292_));
 sg13g2_a21oi_1 _09733_ (.A1(net2269),
    .A2(net1981),
    .Y(_01525_),
    .B1(_02292_));
 sg13g2_nor2_1 _09734_ (.A(net4087),
    .B(net1981),
    .Y(_02293_));
 sg13g2_a21oi_1 _09735_ (.A1(net2267),
    .A2(net1981),
    .Y(_01524_),
    .B1(_02293_));
 sg13g2_nor2_1 _09736_ (.A(net4028),
    .B(net1982),
    .Y(_02294_));
 sg13g2_a21oi_1 _09737_ (.A1(net2260),
    .A2(net1982),
    .Y(_01523_),
    .B1(_02294_));
 sg13g2_nor2_1 _09738_ (.A(net3731),
    .B(_02289_),
    .Y(_02295_));
 sg13g2_a21oi_1 _09739_ (.A1(net2253),
    .A2(net1981),
    .Y(_01522_),
    .B1(_02295_));
 sg13g2_nor2_1 _09740_ (.A(net3783),
    .B(net1981),
    .Y(_02296_));
 sg13g2_a21oi_1 _09741_ (.A1(net2251),
    .A2(net1981),
    .Y(_01521_),
    .B1(_02296_));
 sg13g2_nor2_1 _09742_ (.A(net4219),
    .B(net1982),
    .Y(_02297_));
 sg13g2_a21oi_1 _09743_ (.A1(net2244),
    .A2(net1982),
    .Y(_01520_),
    .B1(_02297_));
 sg13g2_nor3_1 _09744_ (.A(_02103_),
    .B(net2138),
    .C(_02146_),
    .Y(_02298_));
 sg13g2_and2_1 _09745_ (.A(net2328),
    .B(net2094),
    .X(_02299_));
 sg13g2_nor2_1 _09746_ (.A(net3868),
    .B(net2024),
    .Y(_02300_));
 sg13g2_a21oi_1 _09747_ (.A1(net2181),
    .A2(net2024),
    .Y(_01519_),
    .B1(_02300_));
 sg13g2_nor2_1 _09748_ (.A(net3987),
    .B(_02299_),
    .Y(_02301_));
 sg13g2_a21oi_1 _09749_ (.A1(net2274),
    .A2(net2024),
    .Y(_01518_),
    .B1(_02301_));
 sg13g2_nor2_1 _09750_ (.A(net3833),
    .B(net2025),
    .Y(_02302_));
 sg13g2_a21oi_1 _09751_ (.A1(net2269),
    .A2(net2025),
    .Y(_01517_),
    .B1(_02302_));
 sg13g2_nor2_1 _09752_ (.A(net3664),
    .B(net2024),
    .Y(_02303_));
 sg13g2_a21oi_1 _09753_ (.A1(net2264),
    .A2(net2024),
    .Y(_01516_),
    .B1(_02303_));
 sg13g2_nor2_1 _09754_ (.A(net3799),
    .B(net2025),
    .Y(_02304_));
 sg13g2_a21oi_1 _09755_ (.A1(net2260),
    .A2(net2025),
    .Y(_01515_),
    .B1(_02304_));
 sg13g2_nor2_1 _09756_ (.A(net3771),
    .B(net2024),
    .Y(_02305_));
 sg13g2_a21oi_1 _09757_ (.A1(net2254),
    .A2(net2024),
    .Y(_01514_),
    .B1(_02305_));
 sg13g2_nor2_1 _09758_ (.A(net3695),
    .B(net2024),
    .Y(_02306_));
 sg13g2_a21oi_1 _09759_ (.A1(net2248),
    .A2(net2025),
    .Y(_01513_),
    .B1(_02306_));
 sg13g2_nor2_1 _09760_ (.A(net3900),
    .B(net2025),
    .Y(_02307_));
 sg13g2_a21oi_1 _09761_ (.A1(net2243),
    .A2(net2025),
    .Y(_01512_),
    .B1(_02307_));
 sg13g2_nor2_2 _09762_ (.A(net2140),
    .B(_02234_),
    .Y(_02308_));
 sg13g2_nand2_1 _09763_ (.Y(_02309_),
    .A(net2329),
    .B(_02308_));
 sg13g2_nand2_1 _09764_ (.Y(_02310_),
    .A(net3459),
    .B(net1913));
 sg13g2_o21ai_1 _09765_ (.B1(_02310_),
    .Y(_01511_),
    .A1(net2182),
    .A2(net1913));
 sg13g2_nand2_1 _09766_ (.Y(_02311_),
    .A(net3489),
    .B(net1914));
 sg13g2_o21ai_1 _09767_ (.B1(_02311_),
    .Y(_01510_),
    .A1(net2277),
    .A2(net1914));
 sg13g2_nand2_1 _09768_ (.Y(_02312_),
    .A(net3513),
    .B(net1913));
 sg13g2_o21ai_1 _09769_ (.B1(_02312_),
    .Y(_01509_),
    .A1(net2271),
    .A2(net1914));
 sg13g2_nand2_1 _09770_ (.Y(_02313_),
    .A(net3529),
    .B(net1913));
 sg13g2_o21ai_1 _09771_ (.B1(_02313_),
    .Y(_01508_),
    .A1(net2265),
    .A2(net1913));
 sg13g2_nand2_1 _09772_ (.Y(_02314_),
    .A(net3599),
    .B(net1914));
 sg13g2_o21ai_1 _09773_ (.B1(_02314_),
    .Y(_01507_),
    .A1(net2261),
    .A2(net1914));
 sg13g2_nand2_1 _09774_ (.Y(_02315_),
    .A(net3437),
    .B(_02309_));
 sg13g2_o21ai_1 _09775_ (.B1(_02315_),
    .Y(_01506_),
    .A1(net2255),
    .A2(net1913));
 sg13g2_nand2_1 _09776_ (.Y(_02316_),
    .A(net3530),
    .B(net1914));
 sg13g2_o21ai_1 _09777_ (.B1(_02316_),
    .Y(_01505_),
    .A1(net2250),
    .A2(net1914));
 sg13g2_nand2_1 _09778_ (.Y(_02317_),
    .A(net3590),
    .B(net1913));
 sg13g2_o21ai_1 _09779_ (.B1(_02317_),
    .Y(_01504_),
    .A1(net2247),
    .A2(net1913));
 sg13g2_or3_1 _09780_ (.A(_02098_),
    .B(_02099_),
    .C(_02147_),
    .X(_02318_));
 sg13g2_nor2_1 _09781_ (.A(net2140),
    .B(_02318_),
    .Y(_02319_));
 sg13g2_nand2_1 _09782_ (.Y(_02320_),
    .A(net2330),
    .B(net2023));
 sg13g2_nand2_1 _09783_ (.Y(_02321_),
    .A(net3504),
    .B(net1978));
 sg13g2_o21ai_1 _09784_ (.B1(_02321_),
    .Y(_01503_),
    .A1(net2184),
    .A2(net1978));
 sg13g2_nand2_1 _09785_ (.Y(_02322_),
    .A(net3451),
    .B(net1978));
 sg13g2_o21ai_1 _09786_ (.B1(_02322_),
    .Y(_01502_),
    .A1(net2278),
    .A2(net1978));
 sg13g2_nand2_1 _09787_ (.Y(_02323_),
    .A(net3778),
    .B(_02320_));
 sg13g2_o21ai_1 _09788_ (.B1(_02323_),
    .Y(_01501_),
    .A1(net2273),
    .A2(net1979));
 sg13g2_nand2_1 _09789_ (.Y(_02324_),
    .A(net3500),
    .B(net1978));
 sg13g2_o21ai_1 _09790_ (.B1(_02324_),
    .Y(_01500_),
    .A1(net2267),
    .A2(net1978));
 sg13g2_nand2_1 _09791_ (.Y(_02325_),
    .A(net3546),
    .B(net1979));
 sg13g2_o21ai_1 _09792_ (.B1(_02325_),
    .Y(_01499_),
    .A1(net2258),
    .A2(net1979));
 sg13g2_nand2_1 _09793_ (.Y(_02326_),
    .A(net3454),
    .B(net1979));
 sg13g2_o21ai_1 _09794_ (.B1(_02326_),
    .Y(_01498_),
    .A1(net2256),
    .A2(net1979));
 sg13g2_nand2_1 _09795_ (.Y(_02327_),
    .A(net3436),
    .B(net1979));
 sg13g2_o21ai_1 _09796_ (.B1(_02327_),
    .Y(_01497_),
    .A1(net2249),
    .A2(net1979));
 sg13g2_nand2_1 _09797_ (.Y(_02328_),
    .A(net3420),
    .B(net1978));
 sg13g2_o21ai_1 _09798_ (.B1(_02328_),
    .Y(_01496_),
    .A1(net2246),
    .A2(net1978));
 sg13g2_nand3_1 _09799_ (.B(_02102_),
    .C(_02179_),
    .A(_02100_),
    .Y(_02329_));
 sg13g2_nor2_2 _09800_ (.A(_02105_),
    .B(_02329_),
    .Y(_02330_));
 sg13g2_nand2_2 _09801_ (.Y(_02331_),
    .A(net2329),
    .B(net1977));
 sg13g2_nand2_1 _09802_ (.Y(_02332_),
    .A(net3476),
    .B(net1912));
 sg13g2_o21ai_1 _09803_ (.B1(_02332_),
    .Y(_01495_),
    .A1(net2183),
    .A2(net1912));
 sg13g2_nand2_1 _09804_ (.Y(_02333_),
    .A(net3559),
    .B(net1911));
 sg13g2_o21ai_1 _09805_ (.B1(_02333_),
    .Y(_01494_),
    .A1(net2277),
    .A2(net1911));
 sg13g2_nand2_1 _09806_ (.Y(_02334_),
    .A(net3499),
    .B(net1911));
 sg13g2_o21ai_1 _09807_ (.B1(_02334_),
    .Y(_01493_),
    .A1(net2270),
    .A2(net1911));
 sg13g2_nand2_1 _09808_ (.Y(_02335_),
    .A(net3689),
    .B(net1912));
 sg13g2_o21ai_1 _09809_ (.B1(_02335_),
    .Y(_01492_),
    .A1(net2265),
    .A2(net1912));
 sg13g2_nand2_1 _09810_ (.Y(_02336_),
    .A(net3449),
    .B(net1911));
 sg13g2_o21ai_1 _09811_ (.B1(_02336_),
    .Y(_01491_),
    .A1(net2261),
    .A2(net1911));
 sg13g2_nand2_1 _09812_ (.Y(_02337_),
    .A(net3898),
    .B(net1912));
 sg13g2_o21ai_1 _09813_ (.B1(_02337_),
    .Y(_01490_),
    .A1(net2255),
    .A2(net1912));
 sg13g2_nand2_1 _09814_ (.Y(_02338_),
    .A(net3661),
    .B(net1911));
 sg13g2_o21ai_1 _09815_ (.B1(_02338_),
    .Y(_01489_),
    .A1(net2250),
    .A2(net1911));
 sg13g2_nand2_1 _09816_ (.Y(_02339_),
    .A(net3442),
    .B(net1912));
 sg13g2_o21ai_1 _09817_ (.B1(_02339_),
    .Y(_01488_),
    .A1(net2247),
    .A2(net1912));
 sg13g2_nor2_2 _09818_ (.A(net2139),
    .B(_02318_),
    .Y(_02340_));
 sg13g2_nand2_2 _09819_ (.Y(_02341_),
    .A(net2330),
    .B(net2022));
 sg13g2_nand2_1 _09820_ (.Y(_02342_),
    .A(net3618),
    .B(net1975));
 sg13g2_o21ai_1 _09821_ (.B1(_02342_),
    .Y(_01487_),
    .A1(net2183),
    .A2(net1975));
 sg13g2_nand2_1 _09822_ (.Y(_02343_),
    .A(net3541),
    .B(net1976));
 sg13g2_o21ai_1 _09823_ (.B1(_02343_),
    .Y(_01486_),
    .A1(net2276),
    .A2(net1975));
 sg13g2_nand2_1 _09824_ (.Y(_02344_),
    .A(net3439),
    .B(net1975));
 sg13g2_o21ai_1 _09825_ (.B1(_02344_),
    .Y(_01485_),
    .A1(net2271),
    .A2(net1975));
 sg13g2_nand2_1 _09826_ (.Y(_02345_),
    .A(net3472),
    .B(net1975));
 sg13g2_o21ai_1 _09827_ (.B1(_02345_),
    .Y(_01484_),
    .A1(net2266),
    .A2(net1975));
 sg13g2_nand2_1 _09828_ (.Y(_02346_),
    .A(net3419),
    .B(net1976));
 sg13g2_o21ai_1 _09829_ (.B1(_02346_),
    .Y(_01483_),
    .A1(net2258),
    .A2(net1976));
 sg13g2_nand2_1 _09830_ (.Y(_02347_),
    .A(net3600),
    .B(net1976));
 sg13g2_o21ai_1 _09831_ (.B1(_02347_),
    .Y(_01482_),
    .A1(net2256),
    .A2(net1976));
 sg13g2_nand2_1 _09832_ (.Y(_02348_),
    .A(net3438),
    .B(net1976));
 sg13g2_o21ai_1 _09833_ (.B1(_02348_),
    .Y(_01481_),
    .A1(net2249),
    .A2(net1976));
 sg13g2_nand2_1 _09834_ (.Y(_02349_),
    .A(net3467),
    .B(net1976));
 sg13g2_o21ai_1 _09835_ (.B1(_02349_),
    .Y(_01480_),
    .A1(net2246),
    .A2(net1975));
 sg13g2_nor3_1 _09836_ (.A(net2141),
    .B(_02178_),
    .C(_02180_),
    .Y(_02350_));
 sg13g2_and2_1 _09837_ (.A(net2327),
    .B(net2093),
    .X(_02351_));
 sg13g2_nor2_1 _09838_ (.A(net3909),
    .B(net2021),
    .Y(_02352_));
 sg13g2_a21oi_1 _09839_ (.A1(net2180),
    .A2(net2021),
    .Y(_01479_),
    .B1(_02352_));
 sg13g2_nor2_1 _09840_ (.A(net3754),
    .B(net2020),
    .Y(_02353_));
 sg13g2_a21oi_1 _09841_ (.A1(net2275),
    .A2(net2020),
    .Y(_01478_),
    .B1(_02353_));
 sg13g2_nor2_1 _09842_ (.A(net3804),
    .B(net2020),
    .Y(_02354_));
 sg13g2_a21oi_1 _09843_ (.A1(net2269),
    .A2(net2020),
    .Y(_01477_),
    .B1(_02354_));
 sg13g2_nor2_1 _09844_ (.A(net3998),
    .B(net2020),
    .Y(_02355_));
 sg13g2_a21oi_1 _09845_ (.A1(net2267),
    .A2(net2020),
    .Y(_01476_),
    .B1(_02355_));
 sg13g2_nor2_1 _09846_ (.A(net4051),
    .B(net2021),
    .Y(_02356_));
 sg13g2_a21oi_1 _09847_ (.A1(net2260),
    .A2(net2021),
    .Y(_01475_),
    .B1(_02356_));
 sg13g2_nor2_1 _09848_ (.A(net3798),
    .B(net2021),
    .Y(_02357_));
 sg13g2_a21oi_1 _09849_ (.A1(net2253),
    .A2(net2021),
    .Y(_01474_),
    .B1(_02357_));
 sg13g2_nor2_1 _09850_ (.A(net3941),
    .B(net2020),
    .Y(_02358_));
 sg13g2_a21oi_1 _09851_ (.A1(net2251),
    .A2(net2020),
    .Y(_01473_),
    .B1(_02358_));
 sg13g2_nor2_1 _09852_ (.A(net3709),
    .B(net2021),
    .Y(_02359_));
 sg13g2_a21oi_1 _09853_ (.A1(net2244),
    .A2(net2021),
    .Y(_01472_),
    .B1(_02359_));
 sg13g2_nor3_2 _09854_ (.A(net2141),
    .B(_02147_),
    .C(_02178_),
    .Y(_02360_));
 sg13g2_and2_1 _09855_ (.A(net2327),
    .B(net2092),
    .X(_02361_));
 sg13g2_nor2_1 _09856_ (.A(net4288),
    .B(net2018),
    .Y(_02362_));
 sg13g2_a21oi_1 _09857_ (.A1(net2179),
    .A2(net2018),
    .Y(_01471_),
    .B1(_02362_));
 sg13g2_nor2_1 _09858_ (.A(net4066),
    .B(net2019),
    .Y(_02363_));
 sg13g2_a21oi_1 _09859_ (.A1(net2275),
    .A2(net2019),
    .Y(_01470_),
    .B1(_02363_));
 sg13g2_nor2_1 _09860_ (.A(net3925),
    .B(net2018),
    .Y(_02364_));
 sg13g2_a21oi_1 _09861_ (.A1(net2269),
    .A2(net2018),
    .Y(_01469_),
    .B1(_02364_));
 sg13g2_nor2_1 _09862_ (.A(net4274),
    .B(net2018),
    .Y(_02365_));
 sg13g2_a21oi_1 _09863_ (.A1(net2263),
    .A2(net2018),
    .Y(_01468_),
    .B1(_02365_));
 sg13g2_nor2_1 _09864_ (.A(net3884),
    .B(net2019),
    .Y(_02366_));
 sg13g2_a21oi_1 _09865_ (.A1(net2260),
    .A2(net2019),
    .Y(_01467_),
    .B1(_02366_));
 sg13g2_nor2_1 _09866_ (.A(net3852),
    .B(net2019),
    .Y(_02367_));
 sg13g2_a21oi_1 _09867_ (.A1(net2257),
    .A2(_02361_),
    .Y(_01466_),
    .B1(_02367_));
 sg13g2_nor2_1 _09868_ (.A(net3791),
    .B(net2018),
    .Y(_02368_));
 sg13g2_a21oi_1 _09869_ (.A1(net2251),
    .A2(net2018),
    .Y(_01465_),
    .B1(_02368_));
 sg13g2_nor2_1 _09870_ (.A(net4083),
    .B(net2019),
    .Y(_02369_));
 sg13g2_a21oi_1 _09871_ (.A1(net2243),
    .A2(net2019),
    .Y(_01464_),
    .B1(_02369_));
 sg13g2_nor3_1 _09872_ (.A(net2141),
    .B(_02178_),
    .C(_02202_),
    .Y(_02370_));
 sg13g2_and2_1 _09873_ (.A(net2327),
    .B(net2091),
    .X(_02371_));
 sg13g2_nor2_1 _09874_ (.A(net3706),
    .B(net2017),
    .Y(_02372_));
 sg13g2_a21oi_1 _09875_ (.A1(net2179),
    .A2(net2017),
    .Y(_01463_),
    .B1(_02372_));
 sg13g2_nor2_1 _09876_ (.A(net4107),
    .B(_02371_),
    .Y(_02373_));
 sg13g2_a21oi_1 _09877_ (.A1(net2275),
    .A2(net2017),
    .Y(_01462_),
    .B1(_02373_));
 sg13g2_nor2_1 _09878_ (.A(net3735),
    .B(net2017),
    .Y(_02374_));
 sg13g2_a21oi_1 _09879_ (.A1(net2269),
    .A2(net2017),
    .Y(_01461_),
    .B1(_02374_));
 sg13g2_nor2_1 _09880_ (.A(net3776),
    .B(net2016),
    .Y(_02375_));
 sg13g2_a21oi_1 _09881_ (.A1(net2263),
    .A2(net2016),
    .Y(_01460_),
    .B1(_02375_));
 sg13g2_nor2_1 _09882_ (.A(net3707),
    .B(net2017),
    .Y(_02376_));
 sg13g2_a21oi_1 _09883_ (.A1(net2260),
    .A2(net2017),
    .Y(_01459_),
    .B1(_02376_));
 sg13g2_nor2_1 _09884_ (.A(net3967),
    .B(net2016),
    .Y(_02377_));
 sg13g2_a21oi_1 _09885_ (.A1(net2253),
    .A2(net2016),
    .Y(_01458_),
    .B1(_02377_));
 sg13g2_nor2_1 _09886_ (.A(net3970),
    .B(net2016),
    .Y(_02378_));
 sg13g2_a21oi_1 _09887_ (.A1(net2251),
    .A2(net2016),
    .Y(_01457_),
    .B1(_02378_));
 sg13g2_nor2_1 _09888_ (.A(net3667),
    .B(net2016),
    .Y(_02379_));
 sg13g2_a21oi_1 _09889_ (.A1(net2243),
    .A2(net2016),
    .Y(_01456_),
    .B1(_02379_));
 sg13g2_nor3_2 _09890_ (.A(_02103_),
    .B(net2141),
    .C(_02178_),
    .Y(_02380_));
 sg13g2_and2_1 _09891_ (.A(net2331),
    .B(net2090),
    .X(_02381_));
 sg13g2_nor2_1 _09892_ (.A(net3732),
    .B(net2014),
    .Y(_02382_));
 sg13g2_a21oi_1 _09893_ (.A1(net2179),
    .A2(net2014),
    .Y(_01455_),
    .B1(_02382_));
 sg13g2_nor2_1 _09894_ (.A(net3688),
    .B(net2014),
    .Y(_02383_));
 sg13g2_a21oi_1 _09895_ (.A1(net2279),
    .A2(net2014),
    .Y(_01454_),
    .B1(_02383_));
 sg13g2_nor2_1 _09896_ (.A(net3726),
    .B(net2015),
    .Y(_02384_));
 sg13g2_a21oi_1 _09897_ (.A1(net2272),
    .A2(net2015),
    .Y(_01453_),
    .B1(_02384_));
 sg13g2_nor2_1 _09898_ (.A(net3837),
    .B(net2015),
    .Y(_02385_));
 sg13g2_a21oi_1 _09899_ (.A1(net2263),
    .A2(net2015),
    .Y(_01452_),
    .B1(_02385_));
 sg13g2_nor2_1 _09900_ (.A(net4036),
    .B(net2015),
    .Y(_02386_));
 sg13g2_a21oi_1 _09901_ (.A1(net2262),
    .A2(net2015),
    .Y(_01451_),
    .B1(_02386_));
 sg13g2_nor2_1 _09902_ (.A(net3862),
    .B(_02381_),
    .Y(_02387_));
 sg13g2_a21oi_1 _09903_ (.A1(net2257),
    .A2(net2015),
    .Y(_01450_),
    .B1(_02387_));
 sg13g2_nor2_1 _09904_ (.A(net3924),
    .B(net2014),
    .Y(_02388_));
 sg13g2_a21oi_1 _09905_ (.A1(net2251),
    .A2(net2014),
    .Y(_01449_),
    .B1(_02388_));
 sg13g2_nor2_1 _09906_ (.A(net3882),
    .B(net2014),
    .Y(_02389_));
 sg13g2_a21oi_1 _09907_ (.A1(net2243),
    .A2(net2014),
    .Y(_01448_),
    .B1(_02389_));
 sg13g2_nor3_2 _09908_ (.A(net2140),
    .B(_02180_),
    .C(_02223_),
    .Y(_02390_));
 sg13g2_nand2_2 _09909_ (.Y(_02391_),
    .A(net2330),
    .B(_02390_));
 sg13g2_nand2_1 _09910_ (.Y(_02392_),
    .A(net3425),
    .B(net1974));
 sg13g2_o21ai_1 _09911_ (.B1(_02392_),
    .Y(_01447_),
    .A1(net2184),
    .A2(net1974));
 sg13g2_nand2_1 _09912_ (.Y(_02393_),
    .A(net3445),
    .B(net1973));
 sg13g2_o21ai_1 _09913_ (.B1(_02393_),
    .Y(_01446_),
    .A1(net2276),
    .A2(net1973));
 sg13g2_nand2_1 _09914_ (.Y(_02394_),
    .A(net3534),
    .B(net1974));
 sg13g2_o21ai_1 _09915_ (.B1(_02394_),
    .Y(_01445_),
    .A1(net2268),
    .A2(net1974));
 sg13g2_nand2_1 _09916_ (.Y(_02395_),
    .A(net3549),
    .B(net1973));
 sg13g2_o21ai_1 _09917_ (.B1(_02395_),
    .Y(_01444_),
    .A1(net2265),
    .A2(net1973));
 sg13g2_nand2_1 _09918_ (.Y(_02396_),
    .A(net3505),
    .B(net1973));
 sg13g2_o21ai_1 _09919_ (.B1(_02396_),
    .Y(_01443_),
    .A1(net2259),
    .A2(net1973));
 sg13g2_nand2_1 _09920_ (.Y(_02397_),
    .A(net3478),
    .B(net1973));
 sg13g2_o21ai_1 _09921_ (.B1(_02397_),
    .Y(_01442_),
    .A1(net2256),
    .A2(net1973));
 sg13g2_nand2_1 _09922_ (.Y(_02398_),
    .A(net3433),
    .B(net1974));
 sg13g2_o21ai_1 _09923_ (.B1(_02398_),
    .Y(_01441_),
    .A1(net2249),
    .A2(net1974));
 sg13g2_nand2_1 _09924_ (.Y(_02399_),
    .A(net3622),
    .B(net1974));
 sg13g2_o21ai_1 _09925_ (.B1(_02399_),
    .Y(_01440_),
    .A1(net2246),
    .A2(net1974));
 sg13g2_nor3_1 _09926_ (.A(net2140),
    .B(_02147_),
    .C(_02223_),
    .Y(_02400_));
 sg13g2_nand2_2 _09927_ (.Y(_02401_),
    .A(net2330),
    .B(net2012));
 sg13g2_nand2_1 _09928_ (.Y(_02402_),
    .A(net3524),
    .B(net1971));
 sg13g2_o21ai_1 _09929_ (.B1(_02402_),
    .Y(_01439_),
    .A1(net2182),
    .A2(net1971));
 sg13g2_nand2_1 _09930_ (.Y(_02403_),
    .A(net3511),
    .B(net1972));
 sg13g2_o21ai_1 _09931_ (.B1(_02403_),
    .Y(_01438_),
    .A1(net2276),
    .A2(net1972));
 sg13g2_nand2_1 _09932_ (.Y(_02404_),
    .A(net3452),
    .B(net1972));
 sg13g2_o21ai_1 _09933_ (.B1(_02404_),
    .Y(_01437_),
    .A1(net2270),
    .A2(net1972));
 sg13g2_nand2_1 _09934_ (.Y(_02405_),
    .A(net3656),
    .B(net1971));
 sg13g2_o21ai_1 _09935_ (.B1(_02405_),
    .Y(_01436_),
    .A1(net2265),
    .A2(net1971));
 sg13g2_nand2_1 _09936_ (.Y(_02406_),
    .A(net3519),
    .B(net1972));
 sg13g2_o21ai_1 _09937_ (.B1(_02406_),
    .Y(_01435_),
    .A1(net2261),
    .A2(net1972));
 sg13g2_nand2_1 _09938_ (.Y(_02407_),
    .A(net3470),
    .B(net1971));
 sg13g2_o21ai_1 _09939_ (.B1(_02407_),
    .Y(_01434_),
    .A1(net2255),
    .A2(net1971));
 sg13g2_nand2_1 _09940_ (.Y(_02408_),
    .A(net3581),
    .B(net1972));
 sg13g2_o21ai_1 _09941_ (.B1(_02408_),
    .Y(_01433_),
    .A1(net2250),
    .A2(net1972));
 sg13g2_nand2_1 _09942_ (.Y(_02409_),
    .A(net3573),
    .B(net1971));
 sg13g2_o21ai_1 _09943_ (.B1(_02409_),
    .Y(_01432_),
    .A1(net2244),
    .A2(net1971));
 sg13g2_nor3_1 _09944_ (.A(net2140),
    .B(_02202_),
    .C(_02223_),
    .Y(_02410_));
 sg13g2_nand2_1 _09945_ (.Y(_02411_),
    .A(net2330),
    .B(net2011));
 sg13g2_nand2_1 _09946_ (.Y(_02412_),
    .A(net3440),
    .B(net1970));
 sg13g2_o21ai_1 _09947_ (.B1(_02412_),
    .Y(_01431_),
    .A1(net2182),
    .A2(net1970));
 sg13g2_nand2_1 _09948_ (.Y(_02413_),
    .A(net3502),
    .B(net1970));
 sg13g2_o21ai_1 _09949_ (.B1(_02413_),
    .Y(_01430_),
    .A1(net2276),
    .A2(net1970));
 sg13g2_nand2_1 _09950_ (.Y(_02414_),
    .A(net3501),
    .B(net1969));
 sg13g2_o21ai_1 _09951_ (.B1(_02414_),
    .Y(_01429_),
    .A1(net2270),
    .A2(net1969));
 sg13g2_nand2_1 _09952_ (.Y(_02415_),
    .A(net3733),
    .B(net1969));
 sg13g2_o21ai_1 _09953_ (.B1(_02415_),
    .Y(_01428_),
    .A1(net2265),
    .A2(net1969));
 sg13g2_nand2_1 _09954_ (.Y(_02416_),
    .A(net3460),
    .B(_02411_));
 sg13g2_o21ai_1 _09955_ (.B1(_02416_),
    .Y(_01427_),
    .A1(net2261),
    .A2(net1970));
 sg13g2_nand2_1 _09956_ (.Y(_02417_),
    .A(net3535),
    .B(net1969));
 sg13g2_o21ai_1 _09957_ (.B1(_02417_),
    .Y(_01426_),
    .A1(net2255),
    .A2(net1969));
 sg13g2_nand2_1 _09958_ (.Y(_02418_),
    .A(net3473),
    .B(net1970));
 sg13g2_o21ai_1 _09959_ (.B1(_02418_),
    .Y(_01425_),
    .A1(net2250),
    .A2(net1970));
 sg13g2_nand2_1 _09960_ (.Y(_02419_),
    .A(net3523),
    .B(net1969));
 sg13g2_o21ai_1 _09961_ (.B1(_02419_),
    .Y(_01424_),
    .A1(net2246),
    .A2(net1969));
 sg13g2_nor3_2 _09962_ (.A(_02103_),
    .B(net2140),
    .C(_02223_),
    .Y(_02420_));
 sg13g2_nand2_2 _09963_ (.Y(_02421_),
    .A(net2330),
    .B(net2010));
 sg13g2_nand2_1 _09964_ (.Y(_02422_),
    .A(net3547),
    .B(net1968));
 sg13g2_o21ai_1 _09965_ (.B1(_02422_),
    .Y(_01423_),
    .A1(net2183),
    .A2(net1968));
 sg13g2_nand2_1 _09966_ (.Y(_02423_),
    .A(net3503),
    .B(net1968));
 sg13g2_o21ai_1 _09967_ (.B1(_02423_),
    .Y(_01422_),
    .A1(net2278),
    .A2(net1968));
 sg13g2_nand2_1 _09968_ (.Y(_02424_),
    .A(net3441),
    .B(net1968));
 sg13g2_o21ai_1 _09969_ (.B1(_02424_),
    .Y(_01421_),
    .A1(net2273),
    .A2(net1968));
 sg13g2_nand2_1 _09970_ (.Y(_02425_),
    .A(net3466),
    .B(net1968));
 sg13g2_o21ai_1 _09971_ (.B1(_02425_),
    .Y(_01420_),
    .A1(net2266),
    .A2(net1968));
 sg13g2_nand2_1 _09972_ (.Y(_02426_),
    .A(net3446),
    .B(net1967));
 sg13g2_o21ai_1 _09973_ (.B1(_02426_),
    .Y(_01419_),
    .A1(net2259),
    .A2(net1967));
 sg13g2_nand2_1 _09974_ (.Y(_02427_),
    .A(net3426),
    .B(net1967));
 sg13g2_o21ai_1 _09975_ (.B1(_02427_),
    .Y(_01418_),
    .A1(net2256),
    .A2(net1967));
 sg13g2_nand2_1 _09976_ (.Y(_02428_),
    .A(net3507),
    .B(net1967));
 sg13g2_o21ai_1 _09977_ (.B1(_02428_),
    .Y(_01417_),
    .A1(net2250),
    .A2(net1967));
 sg13g2_nand2_1 _09978_ (.Y(_02429_),
    .A(net3484),
    .B(net1967));
 sg13g2_o21ai_1 _09979_ (.B1(_02429_),
    .Y(_01416_),
    .A1(net2246),
    .A2(net1967));
 sg13g2_nor2_2 _09980_ (.A(net2141),
    .B(_02266_),
    .Y(_02430_));
 sg13g2_and2_1 _09981_ (.A(net2327),
    .B(net2009),
    .X(_02431_));
 sg13g2_nor2_1 _09982_ (.A(net3859),
    .B(net1964),
    .Y(_02432_));
 sg13g2_a21oi_1 _09983_ (.A1(net2179),
    .A2(net1964),
    .Y(_01415_),
    .B1(_02432_));
 sg13g2_nor2_1 _09984_ (.A(net3762),
    .B(net1966),
    .Y(_02433_));
 sg13g2_a21oi_1 _09985_ (.A1(net2274),
    .A2(net1966),
    .Y(_01414_),
    .B1(_02433_));
 sg13g2_nor2_1 _09986_ (.A(net3708),
    .B(net1964),
    .Y(_02434_));
 sg13g2_a21oi_1 _09987_ (.A1(net2269),
    .A2(net1964),
    .Y(_01413_),
    .B1(_02434_));
 sg13g2_nor2_1 _09988_ (.A(net3840),
    .B(net1964),
    .Y(_02435_));
 sg13g2_a21oi_1 _09989_ (.A1(net2263),
    .A2(net1964),
    .Y(_01412_),
    .B1(_02435_));
 sg13g2_nor2_1 _09990_ (.A(net3697),
    .B(net1965),
    .Y(_02436_));
 sg13g2_a21oi_1 _09991_ (.A1(net2260),
    .A2(net1965),
    .Y(_01411_),
    .B1(_02436_));
 sg13g2_nor2_1 _09992_ (.A(net3763),
    .B(net1964),
    .Y(_02437_));
 sg13g2_a21oi_1 _09993_ (.A1(net2253),
    .A2(net1964),
    .Y(_01410_),
    .B1(_02437_));
 sg13g2_nor2_1 _09994_ (.A(net3684),
    .B(net1966),
    .Y(_02438_));
 sg13g2_a21oi_1 _09995_ (.A1(net2248),
    .A2(net1966),
    .Y(_01409_),
    .B1(_02438_));
 sg13g2_nor2_1 _09996_ (.A(net3782),
    .B(net1965),
    .Y(_02439_));
 sg13g2_a21oi_1 _09997_ (.A1(net2243),
    .A2(net1965),
    .Y(_01408_),
    .B1(_02439_));
 sg13g2_nor2_2 _09998_ (.A(net2139),
    .B(_02329_),
    .Y(_02440_));
 sg13g2_nand2_1 _09999_ (.Y(_02441_),
    .A(net2329),
    .B(_02440_));
 sg13g2_nand2_1 _10000_ (.Y(_02442_),
    .A(net3443),
    .B(net1910));
 sg13g2_o21ai_1 _10001_ (.B1(_02442_),
    .Y(_01407_),
    .A1(net2182),
    .A2(net1910));
 sg13g2_nand2_1 _10002_ (.Y(_02443_),
    .A(net3583),
    .B(net1909));
 sg13g2_o21ai_1 _10003_ (.B1(_02443_),
    .Y(_01406_),
    .A1(net2277),
    .A2(net1909));
 sg13g2_nand2_1 _10004_ (.Y(_02444_),
    .A(net3598),
    .B(net1910));
 sg13g2_o21ai_1 _10005_ (.B1(_02444_),
    .Y(_01405_),
    .A1(net2270),
    .A2(net1910));
 sg13g2_nand2_1 _10006_ (.Y(_02445_),
    .A(net3471),
    .B(net1909));
 sg13g2_o21ai_1 _10007_ (.B1(_02445_),
    .Y(_01404_),
    .A1(net2266),
    .A2(net1909));
 sg13g2_nand2_1 _10008_ (.Y(_02446_),
    .A(net3475),
    .B(net1910));
 sg13g2_o21ai_1 _10009_ (.B1(_02446_),
    .Y(_01403_),
    .A1(net2261),
    .A2(net1909));
 sg13g2_nand2_1 _10010_ (.Y(_02447_),
    .A(net3558),
    .B(net1909));
 sg13g2_o21ai_1 _10011_ (.B1(_02447_),
    .Y(_01402_),
    .A1(net2256),
    .A2(_02441_));
 sg13g2_nand2_1 _10012_ (.Y(_02448_),
    .A(net3429),
    .B(net1910));
 sg13g2_o21ai_1 _10013_ (.B1(_02448_),
    .Y(_01401_),
    .A1(net2252),
    .A2(net1910));
 sg13g2_nand2_1 _10014_ (.Y(_02449_),
    .A(net3423),
    .B(net1909));
 sg13g2_o21ai_1 _10015_ (.B1(_02449_),
    .Y(_01400_),
    .A1(net2246),
    .A2(net1909));
 sg13g2_nor2_2 _10016_ (.A(net2141),
    .B(_02287_),
    .Y(_02450_));
 sg13g2_and2_1 _10017_ (.A(net2327),
    .B(net2008),
    .X(_02451_));
 sg13g2_nor2_1 _10018_ (.A(net3796),
    .B(net1961),
    .Y(_02452_));
 sg13g2_a21oi_1 _10019_ (.A1(net2180),
    .A2(net1961),
    .Y(_01399_),
    .B1(_02452_));
 sg13g2_nor2_1 _10020_ (.A(net3715),
    .B(net1961),
    .Y(_02453_));
 sg13g2_a21oi_1 _10021_ (.A1(net2279),
    .A2(net1961),
    .Y(_01398_),
    .B1(_02453_));
 sg13g2_nor2_1 _10022_ (.A(net3817),
    .B(net1962),
    .Y(_02454_));
 sg13g2_a21oi_1 _10023_ (.A1(net2272),
    .A2(net1962),
    .Y(_01397_),
    .B1(_02454_));
 sg13g2_nor2_1 _10024_ (.A(net3966),
    .B(net1962),
    .Y(_02455_));
 sg13g2_a21oi_1 _10025_ (.A1(net2263),
    .A2(_02451_),
    .Y(_01396_),
    .B1(_02455_));
 sg13g2_nor2_1 _10026_ (.A(net3777),
    .B(net1961),
    .Y(_02456_));
 sg13g2_a21oi_1 _10027_ (.A1(net2262),
    .A2(net1961),
    .Y(_01395_),
    .B1(_02456_));
 sg13g2_nor2_1 _10028_ (.A(net3692),
    .B(net1962),
    .Y(_02457_));
 sg13g2_a21oi_1 _10029_ (.A1(net2253),
    .A2(net1962),
    .Y(_01394_),
    .B1(_02457_));
 sg13g2_nor2_1 _10030_ (.A(net4102),
    .B(net1961),
    .Y(_02458_));
 sg13g2_a21oi_1 _10031_ (.A1(net2251),
    .A2(net1961),
    .Y(_01393_),
    .B1(_02458_));
 sg13g2_nor2_1 _10032_ (.A(net3855),
    .B(net1962),
    .Y(_02459_));
 sg13g2_a21oi_1 _10033_ (.A1(net2243),
    .A2(net1962),
    .Y(_01392_),
    .B1(_02459_));
 sg13g2_nor3_2 _10034_ (.A(net2139),
    .B(_02147_),
    .C(_02223_),
    .Y(_02460_));
 sg13g2_nand2_2 _10035_ (.Y(_02461_),
    .A(net2330),
    .B(net2007));
 sg13g2_nand2_1 _10036_ (.Y(_02462_),
    .A(net3444),
    .B(net1960));
 sg13g2_o21ai_1 _10037_ (.B1(_02462_),
    .Y(_01106_),
    .A1(net2182),
    .A2(net1960));
 sg13g2_nand2_1 _10038_ (.Y(_02463_),
    .A(net3448),
    .B(net1960));
 sg13g2_o21ai_1 _10039_ (.B1(_02463_),
    .Y(_01105_),
    .A1(net2276),
    .A2(net1960));
 sg13g2_nand2_1 _10040_ (.Y(_02464_),
    .A(net3427),
    .B(net1959));
 sg13g2_o21ai_1 _10041_ (.B1(_02464_),
    .Y(_01104_),
    .A1(net2268),
    .A2(net1959));
 sg13g2_nand2_1 _10042_ (.Y(_02465_),
    .A(net3553),
    .B(net1959));
 sg13g2_o21ai_1 _10043_ (.B1(_02465_),
    .Y(_01103_),
    .A1(net2263),
    .A2(net1959));
 sg13g2_nand2_1 _10044_ (.Y(_02466_),
    .A(net3465),
    .B(net1959));
 sg13g2_o21ai_1 _10045_ (.B1(_02466_),
    .Y(_01102_),
    .A1(net2259),
    .A2(net1959));
 sg13g2_nand2_1 _10046_ (.Y(_02467_),
    .A(net3477),
    .B(net1960));
 sg13g2_o21ai_1 _10047_ (.B1(_02467_),
    .Y(_01101_),
    .A1(net2256),
    .A2(net1960));
 sg13g2_nand2_1 _10048_ (.Y(_02468_),
    .A(net3516),
    .B(net1960));
 sg13g2_o21ai_1 _10049_ (.B1(_02468_),
    .Y(_01100_),
    .A1(net2249),
    .A2(net1960));
 sg13g2_nand2_1 _10050_ (.Y(_02469_),
    .A(net3450),
    .B(net1959));
 sg13g2_o21ai_1 _10051_ (.B1(_02469_),
    .Y(_01099_),
    .A1(net2244),
    .A2(net1959));
 sg13g2_nor3_2 _10052_ (.A(\addr[27] ),
    .B(net2472),
    .C(\addr[25] ),
    .Y(_02470_));
 sg13g2_or3_1 _10053_ (.A(\addr[27] ),
    .B(net2472),
    .C(\addr[25] ),
    .X(_02471_));
 sg13g2_and2_1 _10054_ (.A(_02089_),
    .B(net2388),
    .X(_02472_));
 sg13g2_nand2_2 _10055_ (.Y(_02473_),
    .A(_02089_),
    .B(net2387));
 sg13g2_nor2_1 _10056_ (.A(net2466),
    .B(\addr[6] ),
    .Y(_02474_));
 sg13g2_nand2_2 _10057_ (.Y(_02475_),
    .A(\addr[2] ),
    .B(_02474_));
 sg13g2_nor4_1 _10058_ (.A(\addr[24] ),
    .B(\addr[1] ),
    .C(\addr[8] ),
    .D(\addr[7] ),
    .Y(_02476_));
 sg13g2_nor3_1 _10059_ (.A(\addr[0] ),
    .B(net2472),
    .C(\addr[25] ),
    .Y(_02477_));
 sg13g2_nand3_1 _10060_ (.B(_02476_),
    .C(_02477_),
    .A(\addr[27] ),
    .Y(_02478_));
 sg13g2_nor4_1 _10061_ (.A(\addr[14] ),
    .B(\addr[13] ),
    .C(\addr[16] ),
    .D(\addr[15] ),
    .Y(_02479_));
 sg13g2_nor4_1 _10062_ (.A(\addr[10] ),
    .B(\addr[9] ),
    .C(\addr[12] ),
    .D(\addr[11] ),
    .Y(_02480_));
 sg13g2_nand2_2 _10063_ (.Y(_02481_),
    .A(_02479_),
    .B(_02480_));
 sg13g2_nor3_1 _10064_ (.A(\addr[22] ),
    .B(\addr[21] ),
    .C(\addr[23] ),
    .Y(_02482_));
 sg13g2_nor4_1 _10065_ (.A(\addr[18] ),
    .B(\addr[17] ),
    .C(\addr[20] ),
    .D(\addr[19] ),
    .Y(_02483_));
 sg13g2_nand2_2 _10066_ (.Y(_02484_),
    .A(_02482_),
    .B(_02483_));
 sg13g2_nor3_2 _10067_ (.A(_02478_),
    .B(_02481_),
    .C(_02484_),
    .Y(_02485_));
 sg13g2_and2_1 _10068_ (.A(_02014_),
    .B(_02485_),
    .X(_02486_));
 sg13g2_nand2_2 _10069_ (.Y(_02487_),
    .A(\addr[5] ),
    .B(_02486_));
 sg13g2_nor2_2 _10070_ (.A(_02475_),
    .B(_02487_),
    .Y(_02488_));
 sg13g2_nor3_2 _10071_ (.A(_02478_),
    .B(_02481_),
    .C(_02484_),
    .Y(_02489_));
 sg13g2_a21o_2 _10072_ (.A2(_02488_),
    .A1(net2326),
    .B1(net2414),
    .X(_02490_));
 sg13g2_nor2_1 _10073_ (.A(net4260),
    .B(net2006),
    .Y(_02491_));
 sg13g2_a21oi_1 _10074_ (.A1(net2453),
    .A2(net2006),
    .Y(_00595_),
    .B1(_02491_));
 sg13g2_nor2_1 _10075_ (.A(net3939),
    .B(net2006),
    .Y(_02492_));
 sg13g2_a21oi_1 _10076_ (.A1(_01777_),
    .A2(net2006),
    .Y(_00594_),
    .B1(_02492_));
 sg13g2_nor2_1 _10077_ (.A(net4082),
    .B(net2006),
    .Y(_02493_));
 sg13g2_a21oi_1 _10078_ (.A1(net2452),
    .A2(net2006),
    .Y(_00593_),
    .B1(_02493_));
 sg13g2_nor2_1 _10079_ (.A(net4018),
    .B(net2006),
    .Y(_02494_));
 sg13g2_a21oi_1 _10080_ (.A1(_01779_),
    .A2(net2006),
    .Y(_00592_),
    .B1(_02494_));
 sg13g2_nor2_1 _10081_ (.A(net3916),
    .B(_02490_),
    .Y(_02495_));
 sg13g2_a21oi_1 _10082_ (.A1(_01797_),
    .A2(_02490_),
    .Y(_00591_),
    .B1(_02495_));
 sg13g2_nand2_2 _10083_ (.Y(_02496_),
    .A(net2510),
    .B(\i_tinyqv.cpu.is_auipc ));
 sg13g2_o21ai_1 _10084_ (.B1(_02496_),
    .Y(_02497_),
    .A1(_01963_),
    .A2(_01964_));
 sg13g2_o21ai_1 _10085_ (.B1(net2510),
    .Y(_02498_),
    .A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_auipc ));
 sg13g2_nor2b_2 _10086_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .Y(_02499_));
 sg13g2_nor2_2 _10087_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .Y(_02500_));
 sg13g2_and2_1 _10088_ (.A(_02499_),
    .B(_02500_),
    .X(_02501_));
 sg13g2_and2_1 _10089_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .X(_02502_));
 sg13g2_and2_1 _10090_ (.A(_02500_),
    .B(_02502_),
    .X(_02503_));
 sg13g2_nand2_1 _10091_ (.Y(_02504_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .B(_02503_));
 sg13g2_and2_1 _10092_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .X(_02505_));
 sg13g2_and2_1 _10093_ (.A(_02502_),
    .B(net2386),
    .X(_02506_));
 sg13g2_nor2b_2 _10094_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .Y(_02507_));
 sg13g2_and2_1 _10095_ (.A(_02502_),
    .B(_02507_),
    .X(_02508_));
 sg13g2_a22oi_1 _10096_ (.Y(_02509_),
    .B1(_02508_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .A2(_02506_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ));
 sg13g2_nor2b_2 _10097_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .Y(_02510_));
 sg13g2_and2_1 _10098_ (.A(_02507_),
    .B(net2385),
    .X(_02511_));
 sg13g2_nand3_1 _10099_ (.B(_02507_),
    .C(net2385),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .Y(_02512_));
 sg13g2_nor2b_2 _10100_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .Y(_02513_));
 sg13g2_and2_1 _10101_ (.A(_02499_),
    .B(_02513_),
    .X(_02514_));
 sg13g2_and2_1 _10102_ (.A(_02499_),
    .B(_02507_),
    .X(_02515_));
 sg13g2_nand3_1 _10103_ (.B(_02499_),
    .C(_02507_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .Y(_02516_));
 sg13g2_nor2_2 _10104_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .Y(_02517_));
 sg13g2_and2_1 _10105_ (.A(_02513_),
    .B(_02517_),
    .X(_02518_));
 sg13g2_nand3_1 _10106_ (.B(_02513_),
    .C(_02517_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .Y(_02519_));
 sg13g2_and2_1 _10107_ (.A(_02507_),
    .B(_02517_),
    .X(_02520_));
 sg13g2_nand2_1 _10108_ (.Y(_02521_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .B(_02520_));
 sg13g2_nor2b_1 _10109_ (.A(net2539),
    .B_N(net2538),
    .Y(_02522_));
 sg13g2_nand2b_2 _10110_ (.Y(_02523_),
    .B(net2537),
    .A_N(net2539));
 sg13g2_nand2_2 _10111_ (.Y(_02524_),
    .A(net2536),
    .B(net2384));
 sg13g2_and4_1 _10112_ (.A(net2536),
    .B(_02500_),
    .C(net2385),
    .D(net2384),
    .X(_02525_));
 sg13g2_and2_1 _10113_ (.A(_02502_),
    .B(_02513_),
    .X(_02526_));
 sg13g2_nand2_1 _10114_ (.Y(_02527_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .B(_02526_));
 sg13g2_nand3_1 _10115_ (.B(net2386),
    .C(net2385),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .Y(_02528_));
 sg13g2_and2_1 _10116_ (.A(_02499_),
    .B(net2386),
    .X(_02529_));
 sg13g2_nand3_1 _10117_ (.B(_02499_),
    .C(net2386),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .Y(_02530_));
 sg13g2_and2_1 _10118_ (.A(net2385),
    .B(_02513_),
    .X(_02531_));
 sg13g2_nand2_1 _10119_ (.Y(_02532_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .B(_02531_));
 sg13g2_a221oi_1 _10120_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .C1(_02525_),
    .B1(_02514_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .Y(_02533_),
    .A2(_02501_));
 sg13g2_and4_1 _10121_ (.A(_02504_),
    .B(_02521_),
    .C(_02532_),
    .D(_02533_),
    .X(_02534_));
 sg13g2_and4_1 _10122_ (.A(_02512_),
    .B(_02516_),
    .C(_02519_),
    .D(_02530_),
    .X(_02535_));
 sg13g2_and4_1 _10123_ (.A(_02509_),
    .B(_02527_),
    .C(_02528_),
    .D(_02535_),
    .X(_02536_));
 sg13g2_nand2_2 _10124_ (.Y(_02537_),
    .A(_02534_),
    .B(_02536_));
 sg13g2_nor2_2 _10125_ (.A(net2537),
    .B(net2542),
    .Y(_02538_));
 sg13g2_or2_1 _10126_ (.X(_02539_),
    .B(net2539),
    .A(net2537));
 sg13g2_and2_1 _10127_ (.A(net2537),
    .B(net2541),
    .X(_02540_));
 sg13g2_nand2_1 _10128_ (.Y(_02541_),
    .A(net2537),
    .B(net2541));
 sg13g2_a22oi_1 _10129_ (.Y(_02542_),
    .B1(net2373),
    .B2(\i_tinyqv.cpu.instr_data_start[15] ),
    .A2(net2377),
    .A1(net2574));
 sg13g2_nor2b_1 _10130_ (.A(net2537),
    .B_N(net2541),
    .Y(_02543_));
 sg13g2_nand2b_2 _10131_ (.Y(_02544_),
    .B(net2539),
    .A_N(net2538));
 sg13g2_a22oi_1 _10132_ (.Y(_02545_),
    .B1(net2368),
    .B2(net2572),
    .A2(net2382),
    .A1(\i_tinyqv.cpu.instr_data_start[11] ));
 sg13g2_a21oi_1 _10133_ (.A1(_02542_),
    .A2(_02545_),
    .Y(_02546_),
    .B1(net2532));
 sg13g2_nand2b_2 _10134_ (.Y(_02547_),
    .B(net2534),
    .A_N(net2538));
 sg13g2_nor2_1 _10135_ (.A(net2435),
    .B(_02539_),
    .Y(_02548_));
 sg13g2_nand2_2 _10136_ (.Y(_02549_),
    .A(net2534),
    .B(net2378));
 sg13g2_nor2_2 _10137_ (.A(net2435),
    .B(_02544_),
    .Y(_02550_));
 sg13g2_nand2_2 _10138_ (.Y(_02551_),
    .A(net2534),
    .B(net2369));
 sg13g2_a22oi_1 _10139_ (.Y(_02552_),
    .B1(_02550_),
    .B2(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(net2323),
    .A1(\i_tinyqv.cpu.instr_data_start[19] ));
 sg13g2_nand2b_2 _10140_ (.Y(_02553_),
    .B(_02552_),
    .A_N(_02546_));
 sg13g2_and3_2 _10141_ (.X(_02554_),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .B(net2527),
    .C(net2524));
 sg13g2_nand3_1 _10142_ (.B(net2527),
    .C(net2524),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .Y(_02555_));
 sg13g2_o21ai_1 _10143_ (.B1(_02555_),
    .Y(_02556_),
    .A1(_02498_),
    .A2(_02553_));
 sg13g2_inv_1 _10144_ (.Y(_02557_),
    .A(_02556_));
 sg13g2_o21ai_1 _10145_ (.B1(_02557_),
    .Y(_02558_),
    .A1(_02497_),
    .A2(_02537_));
 sg13g2_o21ai_1 _10146_ (.B1(net2527),
    .Y(_02559_),
    .A1(_01991_),
    .A2(net2434));
 sg13g2_o21ai_1 _10147_ (.B1(net2365),
    .Y(_02560_),
    .A1(\i_tinyqv.cpu.alu_op[3] ),
    .A2(net2527));
 sg13g2_inv_2 _10148_ (.Y(_02561_),
    .A(_02560_));
 sg13g2_and2_1 _10149_ (.A(net2509),
    .B(\i_tinyqv.cpu.is_branch ),
    .X(_02562_));
 sg13g2_nand2_1 _10150_ (.Y(_02563_),
    .A(net2509),
    .B(\i_tinyqv.cpu.is_branch ));
 sg13g2_o21ai_1 _10151_ (.B1(net2509),
    .Y(_02564_),
    .A1(\i_tinyqv.cpu.is_branch ),
    .A2(\i_tinyqv.cpu.is_alu_reg ));
 sg13g2_a21oi_1 _10152_ (.A1(\i_tinyqv.cpu.imm[15] ),
    .A2(net2372),
    .Y(_02565_),
    .B1(net2532));
 sg13g2_a22oi_1 _10153_ (.Y(_02566_),
    .B1(net2367),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .A2(net2376),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[3] ));
 sg13g2_nand2_1 _10154_ (.Y(_02567_),
    .A(_02565_),
    .B(_02566_));
 sg13g2_a21oi_1 _10155_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .A2(net2381),
    .Y(_02568_),
    .B1(_02567_));
 sg13g2_a22oi_1 _10156_ (.Y(_02569_),
    .B1(net2372),
    .B2(\i_tinyqv.cpu.imm[31] ),
    .A2(net2376),
    .A1(\i_tinyqv.cpu.imm[19] ));
 sg13g2_a221oi_1 _10157_ (.B2(\i_tinyqv.cpu.imm[23] ),
    .C1(net2437),
    .B1(net2367),
    .A1(\i_tinyqv.cpu.imm[27] ),
    .Y(_02570_),
    .A2(net2381));
 sg13g2_a21o_2 _10158_ (.A2(_02570_),
    .A1(_02569_),
    .B1(_02568_),
    .X(_02571_));
 sg13g2_nor2b_1 _10159_ (.A(net2514),
    .B_N(net2513),
    .Y(_02572_));
 sg13g2_nand3b_1 _10160_ (.B(net2513),
    .C(net2515),
    .Y(_02573_),
    .A_N(net2514));
 sg13g2_nor2_2 _10161_ (.A(net2516),
    .B(_02573_),
    .Y(_02574_));
 sg13g2_nand2b_1 _10162_ (.Y(_02575_),
    .B(net2515),
    .A_N(net2513));
 sg13g2_nand3b_1 _10163_ (.B(net2515),
    .C(net2514),
    .Y(_02576_),
    .A_N(net2513));
 sg13g2_nor2_2 _10164_ (.A(_01996_),
    .B(_02576_),
    .Y(_02577_));
 sg13g2_nand2_2 _10165_ (.Y(_02578_),
    .A(net2514),
    .B(net2513));
 sg13g2_nor3_2 _10166_ (.A(_01995_),
    .B(_01996_),
    .C(_02578_),
    .Y(_02579_));
 sg13g2_nor2_1 _10167_ (.A(net2514),
    .B(net2513),
    .Y(_02580_));
 sg13g2_nor3_2 _10168_ (.A(net2514),
    .B(net2516),
    .C(_02575_),
    .Y(_02581_));
 sg13g2_nor3_2 _10169_ (.A(_01995_),
    .B(net2516),
    .C(_02578_),
    .Y(_02582_));
 sg13g2_a22oi_1 _10170_ (.Y(_02583_),
    .B1(_02582_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .A2(_02581_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_nor2_2 _10171_ (.A(net2516),
    .B(_02576_),
    .Y(_02584_));
 sg13g2_nor2_2 _10172_ (.A(_01996_),
    .B(_02573_),
    .Y(_02585_));
 sg13g2_nor2_1 _10173_ (.A(net2515),
    .B(net2516),
    .Y(_02586_));
 sg13g2_and2_1 _10174_ (.A(_02572_),
    .B(_02586_),
    .X(_02587_));
 sg13g2_nor2b_1 _10175_ (.A(net2515),
    .B_N(net2516),
    .Y(_02588_));
 sg13g2_nand2b_2 _10176_ (.Y(_02589_),
    .B(net2516),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ));
 sg13g2_and2_1 _10177_ (.A(_02572_),
    .B(_02588_),
    .X(_02590_));
 sg13g2_nand2_1 _10178_ (.Y(_02591_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .B(_02586_));
 sg13g2_nor3_1 _10179_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .B(_02524_),
    .C(_02591_),
    .Y(_02592_));
 sg13g2_and2_1 _10180_ (.A(_02580_),
    .B(_02588_),
    .X(_02593_));
 sg13g2_nor3_2 _10181_ (.A(_01994_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .C(_02589_),
    .Y(_02594_));
 sg13g2_a22oi_1 _10182_ (.Y(_02595_),
    .B1(_02594_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .A2(_02593_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ));
 sg13g2_nor2b_2 _10183_ (.A(_02578_),
    .B_N(_02586_),
    .Y(_02596_));
 sg13g2_nand2_1 _10184_ (.Y(_02597_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .B(_02596_));
 sg13g2_nor2_2 _10185_ (.A(_02578_),
    .B(_02589_),
    .Y(_02598_));
 sg13g2_a22oi_1 _10186_ (.Y(_02599_),
    .B1(_02598_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .A2(_02587_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ));
 sg13g2_a22oi_1 _10187_ (.Y(_02600_),
    .B1(_02590_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A2(_02577_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_a22oi_1 _10188_ (.Y(_02601_),
    .B1(_02584_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .A2(_02574_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ));
 sg13g2_and4_1 _10189_ (.A(_02595_),
    .B(_02599_),
    .C(_02600_),
    .D(_02601_),
    .X(_02602_));
 sg13g2_a221oi_1 _10190_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .C1(_02592_),
    .B1(_02585_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .Y(_02603_),
    .A2(_02579_));
 sg13g2_nand4_1 _10191_ (.B(_02597_),
    .C(_02602_),
    .A(_02583_),
    .Y(_02604_),
    .D(_02603_));
 sg13g2_nor2_1 _10192_ (.A(_02564_),
    .B(_02604_),
    .Y(_02605_));
 sg13g2_a21oi_2 _10193_ (.B1(_02605_),
    .Y(_02606_),
    .A2(_02571_),
    .A1(_02564_));
 sg13g2_xnor2_1 _10194_ (.Y(_02607_),
    .A(_02561_),
    .B(_02606_));
 sg13g2_nor2_1 _10195_ (.A(_02558_),
    .B(_02607_),
    .Y(_02608_));
 sg13g2_a22oi_1 _10196_ (.Y(_02609_),
    .B1(_02515_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A2(_02508_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ));
 sg13g2_nand3_1 _10197_ (.B(_02507_),
    .C(_02517_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .Y(_02610_));
 sg13g2_nand3_1 _10198_ (.B(_02500_),
    .C(_02502_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .Y(_02611_));
 sg13g2_nand3_1 _10199_ (.B(net2386),
    .C(net2385),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .Y(_02612_));
 sg13g2_and2_1 _10200_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .B(_02501_),
    .X(_02613_));
 sg13g2_nand3_1 _10201_ (.B(_02499_),
    .C(_02505_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .Y(_02614_));
 sg13g2_and2_1 _10202_ (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .B(_02511_),
    .X(_02615_));
 sg13g2_nand2_1 _10203_ (.Y(_02616_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .B(_02514_));
 sg13g2_nand3_1 _10204_ (.B(_02513_),
    .C(_02517_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .Y(_02617_));
 sg13g2_a22oi_1 _10205_ (.Y(_02618_),
    .B1(_02526_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .A2(_02506_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ));
 sg13g2_nor2_2 _10206_ (.A(net2535),
    .B(net2379),
    .Y(_02619_));
 sg13g2_nand4_1 _10207_ (.B(net2386),
    .C(_02517_),
    .A(net2436),
    .Y(_02620_),
    .D(net2384));
 sg13g2_nand3_1 _10208_ (.B(_02510_),
    .C(_02513_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .Y(_02621_));
 sg13g2_nand4_1 _10209_ (.B(_02611_),
    .C(_02620_),
    .A(_02610_),
    .Y(_02622_),
    .D(_02621_));
 sg13g2_and4_1 _10210_ (.A(_02609_),
    .B(_02612_),
    .C(_02616_),
    .D(_02618_),
    .X(_02623_));
 sg13g2_nand2_1 _10211_ (.Y(_02624_),
    .A(_02614_),
    .B(_02617_));
 sg13g2_nor4_2 _10212_ (.A(_02613_),
    .B(_02615_),
    .C(_02622_),
    .Y(_02625_),
    .D(_02624_));
 sg13g2_nand2_2 _10213_ (.Y(_02626_),
    .A(_02623_),
    .B(_02625_));
 sg13g2_a22oi_1 _10214_ (.Y(_02627_),
    .B1(net2373),
    .B2(net2568),
    .A2(net2377),
    .A1(\i_tinyqv.cpu.pc[2] ));
 sg13g2_a22oi_1 _10215_ (.Y(_02628_),
    .B1(net2368),
    .B2(\i_tinyqv.cpu.instr_data_start[6] ),
    .A2(net2382),
    .A1(net2571));
 sg13g2_a21oi_1 _10216_ (.A1(_02627_),
    .A2(_02628_),
    .Y(_02629_),
    .B1(net2532));
 sg13g2_a22oi_1 _10217_ (.Y(_02630_),
    .B1(_02550_),
    .B2(\i_tinyqv.cpu.instr_data_start[22] ),
    .A2(net2323),
    .A1(\i_tinyqv.cpu.instr_data_start[18] ));
 sg13g2_nand2b_2 _10218_ (.Y(_02631_),
    .B(_02630_),
    .A_N(_02629_));
 sg13g2_o21ai_1 _10219_ (.B1(_02555_),
    .Y(_02632_),
    .A1(_02498_),
    .A2(_02631_));
 sg13g2_inv_1 _10220_ (.Y(_02633_),
    .A(_02632_));
 sg13g2_o21ai_1 _10221_ (.B1(_02633_),
    .Y(_02634_),
    .A1(_02497_),
    .A2(_02626_));
 sg13g2_a21oi_1 _10222_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .A2(net2367),
    .Y(_02635_),
    .B1(net2532));
 sg13g2_and2_1 _10223_ (.A(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .B(net2376),
    .X(_02636_));
 sg13g2_a221oi_1 _10224_ (.B2(\i_tinyqv.cpu.imm[14] ),
    .C1(_02636_),
    .B1(net2372),
    .A1(net2531),
    .Y(_02637_),
    .A2(net2381));
 sg13g2_a22oi_1 _10225_ (.Y(_02638_),
    .B1(net2372),
    .B2(\i_tinyqv.cpu.imm[30] ),
    .A2(net2376),
    .A1(\i_tinyqv.cpu.imm[18] ));
 sg13g2_a221oi_1 _10226_ (.B2(\i_tinyqv.cpu.imm[22] ),
    .C1(net2437),
    .B1(net2367),
    .A1(\i_tinyqv.cpu.imm[26] ),
    .Y(_02639_),
    .A2(net2381));
 sg13g2_a22oi_1 _10227_ (.Y(_02640_),
    .B1(_02638_),
    .B2(_02639_),
    .A2(_02637_),
    .A1(_02635_));
 sg13g2_inv_1 _10228_ (.Y(_02641_),
    .A(_02640_));
 sg13g2_nand4_1 _10229_ (.B(net2517),
    .C(_02580_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .Y(_02642_),
    .D(_02619_));
 sg13g2_a22oi_1 _10230_ (.Y(_02643_),
    .B1(_02593_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .A2(_02590_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ));
 sg13g2_nand2_1 _10231_ (.Y(_02644_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .B(_02594_));
 sg13g2_a22oi_1 _10232_ (.Y(_02645_),
    .B1(_02598_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .A2(_02582_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ));
 sg13g2_a22oi_1 _10233_ (.Y(_02646_),
    .B1(_02587_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A2(_02581_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ));
 sg13g2_a22oi_1 _10234_ (.Y(_02647_),
    .B1(_02585_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .A2(_02574_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_nand4_1 _10235_ (.B(_02645_),
    .C(_02646_),
    .A(_02643_),
    .Y(_02648_),
    .D(_02647_));
 sg13g2_a22oi_1 _10236_ (.Y(_02649_),
    .B1(_02584_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .A2(_02577_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ));
 sg13g2_a22oi_1 _10237_ (.Y(_02650_),
    .B1(_02596_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .A2(_02579_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ));
 sg13g2_nand4_1 _10238_ (.B(_02644_),
    .C(_02649_),
    .A(_02642_),
    .Y(_02651_),
    .D(_02650_));
 sg13g2_or2_1 _10239_ (.X(_02652_),
    .B(_02651_),
    .A(_02648_));
 sg13g2_mux2_1 _10240_ (.A0(_02652_),
    .A1(_02640_),
    .S(_02564_),
    .X(_02653_));
 sg13g2_xnor2_1 _10241_ (.Y(_02654_),
    .A(_02560_),
    .B(_02653_));
 sg13g2_nand2b_1 _10242_ (.Y(_02655_),
    .B(_02654_),
    .A_N(_02634_));
 sg13g2_inv_1 _10243_ (.Y(_02656_),
    .A(_02655_));
 sg13g2_nand2_1 _10244_ (.Y(_02657_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .B(_02508_));
 sg13g2_a22oi_1 _10245_ (.Y(_02658_),
    .B1(_02520_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .A2(_02518_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_and3_1 _10246_ (.X(_02659_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .B(_02505_),
    .C(net2385));
 sg13g2_nand2_1 _10247_ (.Y(_02660_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .B(_02531_));
 sg13g2_a22oi_1 _10248_ (.Y(_02661_),
    .B1(_02526_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .A2(_02503_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ));
 sg13g2_and3_2 _10249_ (.X(_02662_),
    .A(_02658_),
    .B(_02660_),
    .C(_02661_));
 sg13g2_a221oi_1 _10250_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .C1(_02659_),
    .B1(_02511_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .Y(_02663_),
    .A2(_02506_));
 sg13g2_a22oi_1 _10251_ (.Y(_02664_),
    .B1(_02529_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A2(_02501_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ));
 sg13g2_a22oi_1 _10252_ (.Y(_02665_),
    .B1(_02515_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A2(_02514_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ));
 sg13g2_and4_1 _10253_ (.A(_02657_),
    .B(_02663_),
    .C(_02664_),
    .D(_02665_),
    .X(_02666_));
 sg13g2_nand2_2 _10254_ (.Y(_02667_),
    .A(_02662_),
    .B(_02666_));
 sg13g2_a22oi_1 _10255_ (.Y(_02668_),
    .B1(net2373),
    .B2(net2569),
    .A2(net2381),
    .A1(\i_tinyqv.cpu.instr_data_start[9] ));
 sg13g2_a22oi_1 _10256_ (.Y(_02669_),
    .B1(net2368),
    .B2(\i_tinyqv.cpu.instr_data_start[5] ),
    .A2(net2377),
    .A1(\i_tinyqv.cpu.pc[1] ));
 sg13g2_a21oi_1 _10257_ (.A1(_02668_),
    .A2(_02669_),
    .Y(_02670_),
    .B1(net2532));
 sg13g2_a221oi_1 _10258_ (.B2(\i_tinyqv.cpu.instr_data_start[21] ),
    .C1(_02670_),
    .B1(_02550_),
    .A1(\i_tinyqv.cpu.instr_data_start[17] ),
    .Y(_02671_),
    .A2(net2323));
 sg13g2_a21oi_1 _10259_ (.A1(_02497_),
    .A2(_02671_),
    .Y(_02672_),
    .B1(_02554_));
 sg13g2_o21ai_1 _10260_ (.B1(_02672_),
    .Y(_02673_),
    .A1(_02497_),
    .A2(_02667_));
 sg13g2_inv_1 _10261_ (.Y(_02674_),
    .A(_02673_));
 sg13g2_nand2_1 _10262_ (.Y(_02675_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .B(_02590_));
 sg13g2_a22oi_1 _10263_ (.Y(_02676_),
    .B1(_02582_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A2(_02579_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ));
 sg13g2_a22oi_1 _10264_ (.Y(_02677_),
    .B1(_02584_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .A2(_02577_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ));
 sg13g2_a22oi_1 _10265_ (.Y(_02678_),
    .B1(_02594_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .A2(_02581_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ));
 sg13g2_a22oi_1 _10266_ (.Y(_02679_),
    .B1(_02598_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .A2(_02596_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ));
 sg13g2_a22oi_1 _10267_ (.Y(_02680_),
    .B1(_02585_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A2(_02574_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_a22oi_1 _10268_ (.Y(_02681_),
    .B1(_02593_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .A2(_02587_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ));
 sg13g2_and4_1 _10269_ (.A(_02675_),
    .B(_02677_),
    .C(_02680_),
    .D(_02681_),
    .X(_02682_));
 sg13g2_nand4_1 _10270_ (.B(_02678_),
    .C(_02679_),
    .A(_02676_),
    .Y(_02683_),
    .D(_02682_));
 sg13g2_a22oi_1 _10271_ (.Y(_02684_),
    .B1(net2367),
    .B2(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .A2(net2372),
    .A1(\i_tinyqv.cpu.imm[13] ));
 sg13g2_a221oi_1 _10272_ (.B2(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .C1(net2532),
    .B1(net2376),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .Y(_02685_),
    .A2(net2381));
 sg13g2_and2_1 _10273_ (.A(\i_tinyqv.cpu.imm[21] ),
    .B(net2367),
    .X(_02686_));
 sg13g2_a221oi_1 _10274_ (.B2(\i_tinyqv.cpu.imm[29] ),
    .C1(_02686_),
    .B1(net2372),
    .A1(\i_tinyqv.cpu.imm[25] ),
    .Y(_02687_),
    .A2(net2381));
 sg13g2_a21oi_1 _10275_ (.A1(\i_tinyqv.cpu.imm[17] ),
    .A2(net2376),
    .Y(_02688_),
    .B1(net2437));
 sg13g2_a22oi_1 _10276_ (.Y(_02689_),
    .B1(_02687_),
    .B2(_02688_),
    .A2(_02685_),
    .A1(_02684_));
 sg13g2_mux2_1 _10277_ (.A0(_02683_),
    .A1(_02689_),
    .S(_02564_),
    .X(_02690_));
 sg13g2_xnor2_1 _10278_ (.Y(_02691_),
    .A(_02561_),
    .B(_02690_));
 sg13g2_nand2b_1 _10279_ (.Y(_02692_),
    .B(_02674_),
    .A_N(_02691_));
 sg13g2_nand4_1 _10280_ (.B(net2386),
    .C(_02517_),
    .A(net2536),
    .Y(_02693_),
    .D(net2384));
 sg13g2_nand3_1 _10281_ (.B(net2386),
    .C(net2385),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .Y(_02694_));
 sg13g2_a22oi_1 _10282_ (.Y(_02695_),
    .B1(_02526_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .A2(_02518_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ));
 sg13g2_a22oi_1 _10283_ (.Y(_02696_),
    .B1(_02514_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A2(_02503_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ));
 sg13g2_a22oi_1 _10284_ (.Y(_02697_),
    .B1(_02520_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .A2(_02506_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ));
 sg13g2_a22oi_1 _10285_ (.Y(_02698_),
    .B1(_02531_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A2(_02511_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ));
 sg13g2_a22oi_1 _10286_ (.Y(_02699_),
    .B1(_02529_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .A2(_02515_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_and4_1 _10287_ (.A(_02696_),
    .B(_02697_),
    .C(_02698_),
    .D(_02699_),
    .X(_02700_));
 sg13g2_a22oi_1 _10288_ (.Y(_02701_),
    .B1(_02508_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A2(_02501_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ));
 sg13g2_and4_1 _10289_ (.A(_02693_),
    .B(_02694_),
    .C(_02695_),
    .D(_02701_),
    .X(_02702_));
 sg13g2_nand2_2 _10290_ (.Y(_02703_),
    .A(_02700_),
    .B(_02702_));
 sg13g2_nand3_1 _10291_ (.B(_02700_),
    .C(_02702_),
    .A(_02498_),
    .Y(_02704_));
 sg13g2_nor2_2 _10292_ (.A(net2533),
    .B(net2371),
    .Y(_02705_));
 sg13g2_a22oi_1 _10293_ (.Y(_02706_),
    .B1(_02705_),
    .B2(\i_tinyqv.cpu.instr_data_start[12] ),
    .A2(net2323),
    .A1(net2567));
 sg13g2_nor2_1 _10294_ (.A(net2538),
    .B(net2534),
    .Y(_02707_));
 sg13g2_nor2_2 _10295_ (.A(net2535),
    .B(net2366),
    .Y(_02708_));
 sg13g2_nand2_1 _10296_ (.Y(_02709_),
    .A(\i_tinyqv.cpu.instr_data_start[4] ),
    .B(net2322));
 sg13g2_a22oi_1 _10297_ (.Y(_02710_),
    .B1(_02619_),
    .B2(\i_tinyqv.cpu.instr_data_start[8] ),
    .A2(_02550_),
    .A1(\i_tinyqv.cpu.instr_data_start[20] ));
 sg13g2_nand3_1 _10298_ (.B(_02709_),
    .C(_02710_),
    .A(_02706_),
    .Y(_02711_));
 sg13g2_or2_1 _10299_ (.X(_02712_),
    .B(_02711_),
    .A(_02498_));
 sg13g2_nand3_1 _10300_ (.B(_02704_),
    .C(_02712_),
    .A(net2365),
    .Y(_02713_));
 sg13g2_a21oi_1 _10301_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .A2(net2367),
    .Y(_02714_),
    .B1(net2532));
 sg13g2_and2_1 _10302_ (.A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .B(net2376),
    .X(_02715_));
 sg13g2_a221oi_1 _10303_ (.B2(\i_tinyqv.cpu.imm[12] ),
    .C1(_02715_),
    .B1(net2372),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .Y(_02716_),
    .A2(net2381));
 sg13g2_a22oi_1 _10304_ (.Y(_02717_),
    .B1(net2367),
    .B2(\i_tinyqv.cpu.imm[20] ),
    .A2(net2376),
    .A1(\i_tinyqv.cpu.imm[16] ));
 sg13g2_a221oi_1 _10305_ (.B2(\i_tinyqv.cpu.imm[28] ),
    .C1(net2437),
    .B1(net2372),
    .A1(\i_tinyqv.cpu.imm[24] ),
    .Y(_02718_),
    .A2(net2383));
 sg13g2_a22oi_1 _10306_ (.Y(_02719_),
    .B1(_02717_),
    .B2(_02718_),
    .A2(_02716_),
    .A1(_02714_));
 sg13g2_or4_1 _10307_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .B(_01996_),
    .C(_02524_),
    .D(_02575_),
    .X(_02720_));
 sg13g2_nand2_1 _10308_ (.Y(_02721_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .B(_02582_));
 sg13g2_a22oi_1 _10309_ (.Y(_02722_),
    .B1(_02593_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .A2(_02585_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_a22oi_1 _10310_ (.Y(_02723_),
    .B1(_02584_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .A2(_02577_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_a22oi_1 _10311_ (.Y(_02724_),
    .B1(_02596_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .A2(_02594_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_a22oi_1 _10312_ (.Y(_02725_),
    .B1(_02587_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .A2(_02581_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ));
 sg13g2_and4_1 _10313_ (.A(_02722_),
    .B(_02723_),
    .C(_02724_),
    .D(_02725_),
    .X(_02726_));
 sg13g2_a22oi_1 _10314_ (.Y(_02727_),
    .B1(_02590_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A2(_02574_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ));
 sg13g2_a22oi_1 _10315_ (.Y(_02728_),
    .B1(_02598_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .A2(_02579_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ));
 sg13g2_and4_1 _10316_ (.A(_02720_),
    .B(_02721_),
    .C(_02727_),
    .D(_02728_),
    .X(_02729_));
 sg13g2_nand2_2 _10317_ (.Y(_02730_),
    .A(_02726_),
    .B(_02729_));
 sg13g2_nand3b_1 _10318_ (.B(_02726_),
    .C(_02729_),
    .Y(_02731_),
    .A_N(_02564_));
 sg13g2_nand2b_1 _10319_ (.Y(_02732_),
    .B(_02564_),
    .A_N(_02719_));
 sg13g2_nand2_1 _10320_ (.Y(_02733_),
    .A(_02731_),
    .B(_02732_));
 sg13g2_and3_1 _10321_ (.X(_02734_),
    .A(_02561_),
    .B(_02731_),
    .C(_02732_));
 sg13g2_a21oi_1 _10322_ (.A1(_02731_),
    .A2(_02732_),
    .Y(_02735_),
    .B1(_02561_));
 sg13g2_nor3_1 _10323_ (.A(_02713_),
    .B(_02734_),
    .C(_02735_),
    .Y(_02736_));
 sg13g2_o21ai_1 _10324_ (.B1(_02713_),
    .Y(_02737_),
    .A1(_02734_),
    .A2(_02735_));
 sg13g2_nand2b_1 _10325_ (.Y(_02738_),
    .B(_02737_),
    .A_N(_02736_));
 sg13g2_nor2_1 _10326_ (.A(net2534),
    .B(_02539_),
    .Y(_02739_));
 sg13g2_nand2_1 _10327_ (.Y(_02740_),
    .A(net2435),
    .B(net2378));
 sg13g2_nand2_1 _10328_ (.Y(_02741_),
    .A(\i_tinyqv.cpu.i_core.cy ),
    .B(net2319));
 sg13g2_o21ai_1 _10329_ (.B1(_02741_),
    .Y(_02742_),
    .A1(_02560_),
    .A2(net2319));
 sg13g2_a21oi_1 _10330_ (.A1(_02737_),
    .A2(_02742_),
    .Y(_02743_),
    .B1(_02736_));
 sg13g2_xnor2_1 _10331_ (.Y(_02744_),
    .A(_02673_),
    .B(_02691_));
 sg13g2_o21ai_1 _10332_ (.B1(_02692_),
    .Y(_02745_),
    .A1(_02743_),
    .A2(_02744_));
 sg13g2_nand2b_1 _10333_ (.Y(_02746_),
    .B(_02634_),
    .A_N(_02654_));
 sg13g2_nand2_1 _10334_ (.Y(_02747_),
    .A(_02655_),
    .B(_02746_));
 sg13g2_a21oi_1 _10335_ (.A1(_02745_),
    .A2(_02746_),
    .Y(_02748_),
    .B1(_02656_));
 sg13g2_xnor2_1 _10336_ (.Y(_02749_),
    .A(_02558_),
    .B(_02607_));
 sg13g2_nor2_1 _10337_ (.A(_02748_),
    .B(_02749_),
    .Y(_02750_));
 sg13g2_or2_1 _10338_ (.X(\i_tinyqv.cpu.i_core.cy_out ),
    .B(_02750_),
    .A(_02608_));
 sg13g2_nor2_1 _10339_ (.A(\reset_hold_counter[4] ),
    .B(\reset_hold_counter[3] ),
    .Y(_02751_));
 sg13g2_nor3_1 _10340_ (.A(\reset_hold_counter[2] ),
    .B(\reset_hold_counter[1] ),
    .C(net3430),
    .Y(_02752_));
 sg13g2_nand2_1 _10341_ (.Y(_02753_),
    .A(_02751_),
    .B(_02752_));
 sg13g2_nor2_1 _10342_ (.A(net3405),
    .B(_02753_),
    .Y(_02754_));
 sg13g2_nor3_1 _10343_ (.A(net3405),
    .B(_02026_),
    .C(_02753_),
    .Y(combined_rst_n));
 sg13g2_nand2_2 _10344_ (.Y(_02755_),
    .A(net4920),
    .B(net5142));
 sg13g2_nand2_1 _10345_ (.Y(_02756_),
    .A(net4949),
    .B(net5122));
 sg13g2_and2_1 _10346_ (.A(net2390),
    .B(_02756_),
    .X(_02757_));
 sg13g2_and2_1 _10347_ (.A(_02755_),
    .B(_02757_),
    .X(_02758_));
 sg13g2_nand2_1 _10348_ (.Y(_02759_),
    .A(net2612),
    .B(_02757_));
 sg13g2_o21ai_1 _10349_ (.B1(_02759_),
    .Y(_02760_),
    .A1(net2613),
    .A2(_02758_));
 sg13g2_nand2_1 _10350_ (.Y(_02761_),
    .A(net2613),
    .B(_02758_));
 sg13g2_o21ai_1 _10351_ (.B1(_02761_),
    .Y(_02762_),
    .A1(net2612),
    .A2(_02757_));
 sg13g2_nor2_2 _10352_ (.A(_02760_),
    .B(_02762_),
    .Y(_02763_));
 sg13g2_and2_1 _10353_ (.A(net4873),
    .B(_02763_),
    .X(_00098_));
 sg13g2_nor2_1 _10354_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.is_load ),
    .Y(_02764_));
 sg13g2_and2_1 _10355_ (.A(net2510),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .X(_02765_));
 sg13g2_nand2_1 _10356_ (.Y(_02766_),
    .A(net2510),
    .B(\i_tinyqv.cpu.no_write_in_progress ));
 sg13g2_nand2_1 _10357_ (.Y(_02767_),
    .A(net2511),
    .B(_02764_));
 sg13g2_o21ai_1 _10358_ (.B1(net2511),
    .Y(_02768_),
    .A1(net5124),
    .A2(_02764_));
 sg13g2_nor2_2 _10359_ (.A(net2435),
    .B(net2370),
    .Y(_02769_));
 sg13g2_nand2_2 _10360_ (.Y(_02770_),
    .A(net2535),
    .B(net2374));
 sg13g2_a21oi_1 _10361_ (.A1(_02558_),
    .A2(_02606_),
    .Y(_02771_),
    .B1(_02559_));
 sg13g2_o21ai_1 _10362_ (.B1(_02771_),
    .Y(_02772_),
    .A1(_02748_),
    .A2(_02749_));
 sg13g2_o21ai_1 _10363_ (.B1(_02559_),
    .Y(_02773_),
    .A1(\i_tinyqv.cpu.i_core.cmp ),
    .A2(net2320));
 sg13g2_xor2_1 _10364_ (.B(_02733_),
    .A(_02713_),
    .X(_02774_));
 sg13g2_nand2_1 _10365_ (.Y(_02775_),
    .A(_02674_),
    .B(_02690_));
 sg13g2_xnor2_1 _10366_ (.Y(_02776_),
    .A(_02673_),
    .B(_02690_));
 sg13g2_nor2b_1 _10367_ (.A(_02606_),
    .B_N(_02558_),
    .Y(_02777_));
 sg13g2_nand2b_1 _10368_ (.Y(_02778_),
    .B(_02606_),
    .A_N(_02558_));
 sg13g2_xor2_1 _10369_ (.B(_02606_),
    .A(_02558_),
    .X(_02779_));
 sg13g2_nand2b_1 _10370_ (.Y(_02780_),
    .B(_02653_),
    .A_N(_02634_));
 sg13g2_nor2b_1 _10371_ (.A(_02653_),
    .B_N(_02634_),
    .Y(_02781_));
 sg13g2_xnor2_1 _10372_ (.Y(_02782_),
    .A(_02634_),
    .B(_02653_));
 sg13g2_nand2b_1 _10373_ (.Y(_02783_),
    .B(_02779_),
    .A_N(_02773_));
 sg13g2_nor4_1 _10374_ (.A(_02774_),
    .B(_02776_),
    .C(_02782_),
    .D(_02783_),
    .Y(_02784_));
 sg13g2_inv_1 _10375_ (.Y(_02785_),
    .A(_02784_));
 sg13g2_nor4_1 _10376_ (.A(_02001_),
    .B(_02554_),
    .C(_02608_),
    .D(_02750_),
    .Y(_02786_));
 sg13g2_a22oi_1 _10377_ (.Y(_02787_),
    .B1(_02772_),
    .B2(_02785_),
    .A2(net2365),
    .A1(net2529));
 sg13g2_or2_1 _10378_ (.X(\i_tinyqv.cpu.i_core.cmp_out ),
    .B(_02787_),
    .A(_02786_));
 sg13g2_nor3_1 _10379_ (.A(_02001_),
    .B(_02786_),
    .C(_02787_),
    .Y(_02788_));
 sg13g2_a21oi_1 _10380_ (.A1(_02772_),
    .A2(_02785_),
    .Y(_02789_),
    .B1(net2529));
 sg13g2_or3_1 _10381_ (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .B(net2365),
    .C(_02789_),
    .X(_02790_));
 sg13g2_nand2_2 _10382_ (.Y(_02791_),
    .A(net2511),
    .B(net5029));
 sg13g2_o21ai_1 _10383_ (.B1(net2512),
    .Y(_02792_),
    .A1(\i_tinyqv.cpu.is_alu_reg ),
    .A2(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_nor2_1 _10384_ (.A(net2527),
    .B(_02001_),
    .Y(_02793_));
 sg13g2_nand2b_2 _10385_ (.Y(_02794_),
    .B(net2530),
    .A_N(net2528));
 sg13g2_nor2b_2 _10386_ (.A(net2524),
    .B_N(net2527),
    .Y(_02795_));
 sg13g2_inv_1 _10387_ (.Y(_02796_),
    .A(_02795_));
 sg13g2_nor2_1 _10388_ (.A(_02793_),
    .B(_02795_),
    .Y(_02797_));
 sg13g2_xnor2_1 _10389_ (.Y(_02798_),
    .A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .B(_02797_));
 sg13g2_nand4_1 _10390_ (.B(\i_tinyqv.cpu.i_core.load_done ),
    .C(_02765_),
    .A(\i_tinyqv.cpu.is_load ),
    .Y(_02799_),
    .D(_02792_));
 sg13g2_and2_1 _10391_ (.A(net2365),
    .B(_02799_),
    .X(_02800_));
 sg13g2_o21ai_1 _10392_ (.B1(_02800_),
    .Y(_02801_),
    .A1(_02792_),
    .A2(_02798_));
 sg13g2_o21ai_1 _10393_ (.B1(_02801_),
    .Y(_02802_),
    .A1(_02788_),
    .A2(_02790_));
 sg13g2_a21oi_2 _10394_ (.B1(_01963_),
    .Y(_02803_),
    .A2(_01965_),
    .A1(_01964_));
 sg13g2_nand2_2 _10395_ (.Y(_02804_),
    .A(net2511),
    .B(\i_tinyqv.cpu.is_lui ));
 sg13g2_nand2_1 _10396_ (.Y(_02805_),
    .A(_02496_),
    .B(_02804_));
 sg13g2_or2_1 _10397_ (.X(_02806_),
    .B(_02805_),
    .A(_02803_));
 sg13g2_and2_1 _10398_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .X(_02807_));
 sg13g2_nand2_1 _10399_ (.Y(_02808_),
    .A(net5112),
    .B(net5073));
 sg13g2_and2_1 _10400_ (.A(net2510),
    .B(\i_tinyqv.cpu.is_system ),
    .X(_02809_));
 sg13g2_nand2_2 _10401_ (.Y(_02810_),
    .A(net2510),
    .B(\i_tinyqv.cpu.is_system ));
 sg13g2_or4_1 _10402_ (.A(net4937),
    .B(net2364),
    .C(net2357),
    .D(_02809_),
    .X(_02811_));
 sg13g2_nor3_1 _10403_ (.A(_02768_),
    .B(_02806_),
    .C(_02811_),
    .Y(_02812_));
 sg13g2_a21oi_2 _10404_ (.B1(net2315),
    .Y(_02813_),
    .A2(_02812_),
    .A1(_02802_));
 sg13g2_a221oi_1 _10405_ (.B2(_02812_),
    .C1(net2315),
    .B1(_02802_),
    .A1(_02766_),
    .Y(_02814_),
    .A2(_02767_));
 sg13g2_nand2b_1 _10406_ (.Y(_02815_),
    .B(_02813_),
    .A_N(_02768_));
 sg13g2_a21o_1 _10407_ (.A2(_02813_),
    .A1(net4937),
    .B1(_02814_),
    .X(_00045_));
 sg13g2_and2_1 _10408_ (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .B(net2616),
    .X(uio_oe[5]));
 sg13g2_mux2_1 _10409_ (.A0(\i_uart_tx.txd_reg ),
    .A1(\gpio_out[0] ),
    .S(\gpio_out_sel[0] ),
    .X(uo_out[0]));
 sg13g2_nand2b_2 _10410_ (.Y(uo_out[1]),
    .B(\gpio_out_sel[1] ),
    .A_N(\gpio_out[1] ));
 sg13g2_mux2_1 _10411_ (.A0(\i_i2c_peri.i_i2c.scl_o_reg ),
    .A1(\gpio_out[2] ),
    .S(\gpio_out_sel[2] ),
    .X(uo_out[2]));
 sg13g2_mux2_1 _10412_ (.A0(\i_spi.data[7] ),
    .A1(\gpio_out[3] ),
    .S(\gpio_out_sel[3] ),
    .X(uo_out[3]));
 sg13g2_mux2_1 _10413_ (.A0(\i_spi.spi_select ),
    .A1(\gpio_out[4] ),
    .S(\gpio_out_sel[4] ),
    .X(uo_out[4]));
 sg13g2_mux2_1 _10414_ (.A0(\i_spi.spi_clk_out ),
    .A1(\gpio_out[5] ),
    .S(\gpio_out_sel[5] ),
    .X(uo_out[5]));
 sg13g2_mux2_1 _10415_ (.A0(\i_i2c_peri.i_i2c.sda_o_reg ),
    .A1(\gpio_out[6] ),
    .S(\gpio_out_sel[6] ),
    .X(uo_out[6]));
 sg13g2_nand2_1 _10416_ (.Y(_02816_),
    .A(\i_tinyqv.mem.q_ctrl.spi_clk_neg ),
    .B(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ));
 sg13g2_o21ai_1 _10417_ (.B1(_02816_),
    .Y(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .A1(_01982_),
    .A2(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ));
 sg13g2_nor2_2 _10418_ (.A(net4136),
    .B(\i_tinyqv.cpu.i_core.cycle[0] ),
    .Y(_02817_));
 sg13g2_or2_1 _10419_ (.X(_02818_),
    .B(net5156),
    .A(net4136));
 sg13g2_nand4_1 _10420_ (.B(_02765_),
    .C(net2317),
    .A(net5112),
    .Y(_02819_),
    .D(_02817_));
 sg13g2_nor4_1 _10421_ (.A(_02764_),
    .B(_02766_),
    .C(net2315),
    .D(_02818_),
    .Y(_02820_));
 sg13g2_and2_1 _10422_ (.A(\i_tinyqv.cpu.is_store ),
    .B(net2240),
    .X(_02821_));
 sg13g2_nor2_1 _10423_ (.A(net5050),
    .B(net5352),
    .Y(_02822_));
 sg13g2_nor3_2 _10424_ (.A(net4315),
    .B(net5050),
    .C(net5352),
    .Y(_02823_));
 sg13g2_nand2b_2 _10425_ (.Y(_02824_),
    .B(_02822_),
    .A_N(net4315));
 sg13g2_o21ai_1 _10426_ (.B1(net2501),
    .Y(_02825_),
    .A1(net3652),
    .A2(_02821_));
 sg13g2_a21oi_1 _10427_ (.A1(_02821_),
    .A2(_02823_),
    .Y(_02826_),
    .B1(_02825_));
 sg13g2_nand2_2 _10428_ (.Y(_02827_),
    .A(_02814_),
    .B(_02823_));
 sg13g2_nand2_1 _10429_ (.Y(_02828_),
    .A(\i_tinyqv.cpu.is_load ),
    .B(_02827_));
 sg13g2_nand3_1 _10430_ (.B(net2240),
    .C(_02827_),
    .A(net5326),
    .Y(_02829_));
 sg13g2_mux2_1 _10431_ (.A0(_02824_),
    .A1(_02826_),
    .S(_02829_),
    .X(_00044_));
 sg13g2_a21oi_1 _10432_ (.A1(_02623_),
    .A2(_02625_),
    .Y(_02830_),
    .B1(_01962_));
 sg13g2_a21oi_1 _10433_ (.A1(_02700_),
    .A2(_02702_),
    .Y(_02831_),
    .B1(_01962_));
 sg13g2_a21oi_1 _10434_ (.A1(_02534_),
    .A2(_02536_),
    .Y(_02832_),
    .B1(_01962_));
 sg13g2_a21oi_1 _10435_ (.A1(_02662_),
    .A2(_02666_),
    .Y(_02833_),
    .B1(_01962_));
 sg13g2_nor4_1 _10436_ (.A(net2137),
    .B(net2133),
    .C(net2131),
    .D(net2128),
    .Y(_02834_));
 sg13g2_nand2_1 _10437_ (.Y(_02835_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net2133));
 sg13g2_nand2_1 _10438_ (.Y(_02836_),
    .A(net2588),
    .B(net2137));
 sg13g2_nand2_1 _10439_ (.Y(_02837_),
    .A(net2589),
    .B(net2128));
 sg13g2_nor2_1 _10440_ (.A(_02836_),
    .B(_02837_),
    .Y(_02838_));
 sg13g2_a22oi_1 _10441_ (.Y(_02839_),
    .B1(net2128),
    .B2(net2588),
    .A2(net2137),
    .A1(net2589));
 sg13g2_nor2_1 _10442_ (.A(_02838_),
    .B(_02839_),
    .Y(_02840_));
 sg13g2_nor2b_1 _10443_ (.A(_02835_),
    .B_N(_02840_),
    .Y(_02841_));
 sg13g2_and2_1 _10444_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net2133),
    .X(_02842_));
 sg13g2_nand2_1 _10445_ (.Y(_02843_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net2128));
 sg13g2_and2_1 _10446_ (.A(net2588),
    .B(net2131),
    .X(_02844_));
 sg13g2_and4_1 _10447_ (.A(net2588),
    .B(net2589),
    .C(net2137),
    .D(net2131),
    .X(_02845_));
 sg13g2_a22oi_1 _10448_ (.Y(_02846_),
    .B1(net2131),
    .B2(net2589),
    .A2(net2137),
    .A1(net2588));
 sg13g2_or3_1 _10449_ (.A(_02843_),
    .B(_02845_),
    .C(_02846_),
    .X(_02847_));
 sg13g2_o21ai_1 _10450_ (.B1(_02843_),
    .Y(_02848_),
    .A1(_02845_),
    .A2(_02846_));
 sg13g2_nand3_1 _10451_ (.B(_02847_),
    .C(_02848_),
    .A(_02838_),
    .Y(_02849_));
 sg13g2_a21o_1 _10452_ (.A2(_02848_),
    .A1(_02847_),
    .B1(_02838_),
    .X(_02850_));
 sg13g2_nand3_1 _10453_ (.B(_02849_),
    .C(_02850_),
    .A(_02842_),
    .Y(_02851_));
 sg13g2_a21o_1 _10454_ (.A2(_02850_),
    .A1(_02849_),
    .B1(_02842_),
    .X(_02852_));
 sg13g2_nand3_1 _10455_ (.B(_02851_),
    .C(_02852_),
    .A(_02841_),
    .Y(_02853_));
 sg13g2_a21o_1 _10456_ (.A2(_02852_),
    .A1(_02851_),
    .B1(_02841_),
    .X(_02854_));
 sg13g2_nand3_1 _10457_ (.B(_02853_),
    .C(_02854_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .Y(_02855_));
 sg13g2_a21o_1 _10458_ (.A2(_02854_),
    .A1(_02853_),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .X(_02856_));
 sg13g2_nand4_1 _10459_ (.B(net2589),
    .C(net2133),
    .A(net2588),
    .Y(_02857_),
    .D(net2128));
 sg13g2_inv_1 _10460_ (.Y(_02858_),
    .A(_02857_));
 sg13g2_xnor2_1 _10461_ (.Y(_02859_),
    .A(_02835_),
    .B(_02840_));
 sg13g2_and2_1 _10462_ (.A(_02858_),
    .B(_02859_),
    .X(_02860_));
 sg13g2_xnor2_1 _10463_ (.Y(_02861_),
    .A(_02857_),
    .B(_02859_));
 sg13g2_a21o_1 _10464_ (.A2(_02861_),
    .A1(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .B1(_02860_),
    .X(_02862_));
 sg13g2_and3_1 _10465_ (.X(_02863_),
    .A(_02855_),
    .B(_02856_),
    .C(_02862_));
 sg13g2_nand3_1 _10466_ (.B(_02856_),
    .C(_02862_),
    .A(_02855_),
    .Y(_02864_));
 sg13g2_nand2_1 _10467_ (.Y(_02865_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(net2133));
 sg13g2_a21oi_1 _10468_ (.A1(_02837_),
    .A2(_02865_),
    .Y(_02866_),
    .B1(_02858_));
 sg13g2_nand3_1 _10469_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .C(net2133),
    .A(net2589),
    .Y(_02867_));
 sg13g2_xnor2_1 _10470_ (.Y(_02868_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .B(_02866_));
 sg13g2_nor2_1 _10471_ (.A(_02867_),
    .B(_02868_),
    .Y(_02869_));
 sg13g2_a21oi_1 _10472_ (.A1(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .A2(_02866_),
    .Y(_02870_),
    .B1(_02869_));
 sg13g2_xnor2_1 _10473_ (.Y(_02871_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .B(_02861_));
 sg13g2_or2_1 _10474_ (.X(_02872_),
    .B(_02871_),
    .A(_02870_));
 sg13g2_a21oi_1 _10475_ (.A1(_02855_),
    .A2(_02856_),
    .Y(_02873_),
    .B1(_02862_));
 sg13g2_or2_1 _10476_ (.X(_02874_),
    .B(_02873_),
    .A(_02863_));
 sg13g2_nor2_1 _10477_ (.A(_02872_),
    .B(_02874_),
    .Y(_02875_));
 sg13g2_nor2_1 _10478_ (.A(_02863_),
    .B(_02875_),
    .Y(_02876_));
 sg13g2_o21ai_1 _10479_ (.B1(_02864_),
    .Y(_02877_),
    .A1(_02872_),
    .A2(_02873_));
 sg13g2_nand2_1 _10480_ (.Y(_02878_),
    .A(_02849_),
    .B(_02851_));
 sg13g2_nand2_1 _10481_ (.Y(_02879_),
    .A(net2587),
    .B(net2133));
 sg13g2_nand2b_1 _10482_ (.Y(_02880_),
    .B(_02847_),
    .A_N(_02845_));
 sg13g2_nand2_1 _10483_ (.Y(_02881_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net2128));
 sg13g2_nand2_2 _10484_ (.Y(_02882_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net2131));
 sg13g2_nand2_1 _10485_ (.Y(_02883_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net2137));
 sg13g2_xnor2_1 _10486_ (.Y(_02884_),
    .A(_02844_),
    .B(_02883_));
 sg13g2_nand2b_1 _10487_ (.Y(_02885_),
    .B(_02884_),
    .A_N(_02881_));
 sg13g2_xnor2_1 _10488_ (.Y(_02886_),
    .A(_02881_),
    .B(_02884_));
 sg13g2_nand2_1 _10489_ (.Y(_02887_),
    .A(_02880_),
    .B(_02886_));
 sg13g2_xnor2_1 _10490_ (.Y(_02888_),
    .A(_02880_),
    .B(_02886_));
 sg13g2_xor2_1 _10491_ (.B(_02888_),
    .A(_02879_),
    .X(_02889_));
 sg13g2_nand2_1 _10492_ (.Y(_02890_),
    .A(_02878_),
    .B(_02889_));
 sg13g2_xnor2_1 _10493_ (.Y(_02891_),
    .A(_02878_),
    .B(_02889_));
 sg13g2_xnor2_1 _10494_ (.Y(_02892_),
    .A(_02049_),
    .B(_02891_));
 sg13g2_nand2_1 _10495_ (.Y(_02893_),
    .A(_02853_),
    .B(_02855_));
 sg13g2_nor2b_1 _10496_ (.A(_02892_),
    .B_N(_02893_),
    .Y(_02894_));
 sg13g2_xnor2_1 _10497_ (.Y(_02895_),
    .A(_02892_),
    .B(_02893_));
 sg13g2_inv_1 _10498_ (.Y(_02896_),
    .A(_02895_));
 sg13g2_nand2_1 _10499_ (.Y(_02897_),
    .A(_02877_),
    .B(_02895_));
 sg13g2_a21oi_1 _10500_ (.A1(_02876_),
    .A2(_02896_),
    .Y(_02898_),
    .B1(_02834_));
 sg13g2_a22oi_1 _10501_ (.Y(_02899_),
    .B1(_02897_),
    .B2(_02898_),
    .A2(_02834_),
    .A1(net4776));
 sg13g2_inv_1 _10502_ (.Y(_00000_),
    .A(_02899_));
 sg13g2_a21oi_1 _10503_ (.A1(_02877_),
    .A2(_02895_),
    .Y(_02900_),
    .B1(_02894_));
 sg13g2_o21ai_1 _10504_ (.B1(_02887_),
    .Y(_02901_),
    .A1(_02879_),
    .A2(_02888_));
 sg13g2_nand2_1 _10505_ (.Y(_02902_),
    .A(net2586),
    .B(net2133));
 sg13g2_o21ai_1 _10506_ (.B1(_02885_),
    .Y(_02903_),
    .A1(_02836_),
    .A2(_02882_));
 sg13g2_and2_1 _10507_ (.A(net2587),
    .B(net2128),
    .X(_02904_));
 sg13g2_nand2_1 _10508_ (.Y(_02905_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net2130));
 sg13g2_nand2_1 _10509_ (.Y(_02906_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net2137));
 sg13g2_xor2_1 _10510_ (.B(_02906_),
    .A(_02882_),
    .X(_02907_));
 sg13g2_nand2_1 _10511_ (.Y(_02908_),
    .A(_02904_),
    .B(_02907_));
 sg13g2_xor2_1 _10512_ (.B(_02907_),
    .A(_02904_),
    .X(_02909_));
 sg13g2_nand2_1 _10513_ (.Y(_02910_),
    .A(_02903_),
    .B(_02909_));
 sg13g2_xnor2_1 _10514_ (.Y(_02911_),
    .A(_02903_),
    .B(_02909_));
 sg13g2_xor2_1 _10515_ (.B(_02911_),
    .A(_02902_),
    .X(_02912_));
 sg13g2_nand2_1 _10516_ (.Y(_02913_),
    .A(_02901_),
    .B(_02912_));
 sg13g2_xnor2_1 _10517_ (.Y(_02914_),
    .A(_02901_),
    .B(_02912_));
 sg13g2_xnor2_1 _10518_ (.Y(_02915_),
    .A(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .B(_02914_));
 sg13g2_o21ai_1 _10519_ (.B1(_02890_),
    .Y(_02916_),
    .A1(_02049_),
    .A2(_02891_));
 sg13g2_nor2_1 _10520_ (.A(_02915_),
    .B(_02916_),
    .Y(_02917_));
 sg13g2_xnor2_1 _10521_ (.Y(_02918_),
    .A(_02915_),
    .B(_02916_));
 sg13g2_xor2_1 _10522_ (.B(_02918_),
    .A(_02900_),
    .X(_00003_));
 sg13g2_o21ai_1 _10523_ (.B1(_02910_),
    .Y(_02919_),
    .A1(_02902_),
    .A2(_02911_));
 sg13g2_nand2_1 _10524_ (.Y(_02920_),
    .A(net2585),
    .B(net2134));
 sg13g2_o21ai_1 _10525_ (.B1(_02908_),
    .Y(_02921_),
    .A1(_02882_),
    .A2(_02906_));
 sg13g2_nand2_1 _10526_ (.Y(_02922_),
    .A(net2586),
    .B(net2127));
 sg13g2_nand2_1 _10527_ (.Y(_02923_),
    .A(net2587),
    .B(net2130));
 sg13g2_nand2_1 _10528_ (.Y(_02924_),
    .A(net2587),
    .B(net2136));
 sg13g2_xor2_1 _10529_ (.B(_02924_),
    .A(_02905_),
    .X(_02925_));
 sg13g2_nand2b_1 _10530_ (.Y(_02926_),
    .B(_02925_),
    .A_N(_02922_));
 sg13g2_xnor2_1 _10531_ (.Y(_02927_),
    .A(_02922_),
    .B(_02925_));
 sg13g2_nand2_1 _10532_ (.Y(_02928_),
    .A(_02921_),
    .B(_02927_));
 sg13g2_xnor2_1 _10533_ (.Y(_02929_),
    .A(_02921_),
    .B(_02927_));
 sg13g2_xor2_1 _10534_ (.B(_02929_),
    .A(_02920_),
    .X(_02930_));
 sg13g2_nand2_1 _10535_ (.Y(_02931_),
    .A(_02919_),
    .B(_02930_));
 sg13g2_xnor2_1 _10536_ (.Y(_02932_),
    .A(_02919_),
    .B(_02930_));
 sg13g2_xnor2_1 _10537_ (.Y(_02933_),
    .A(_02051_),
    .B(_02932_));
 sg13g2_o21ai_1 _10538_ (.B1(_02913_),
    .Y(_02934_),
    .A1(_02050_),
    .A2(_02914_));
 sg13g2_nor2b_1 _10539_ (.A(_02933_),
    .B_N(_02934_),
    .Y(_02935_));
 sg13g2_inv_1 _10540_ (.Y(_02936_),
    .A(_02935_));
 sg13g2_xor2_1 _10541_ (.B(_02934_),
    .A(_02933_),
    .X(_02937_));
 sg13g2_a221oi_1 _10542_ (.B2(_02916_),
    .C1(_02894_),
    .B1(_02915_),
    .A1(_02877_),
    .Y(_02938_),
    .A2(_02895_));
 sg13g2_or3_1 _10543_ (.A(_02917_),
    .B(_02937_),
    .C(_02938_),
    .X(_02939_));
 sg13g2_o21ai_1 _10544_ (.B1(_02937_),
    .Y(_02940_),
    .A1(_02917_),
    .A2(_02938_));
 sg13g2_and2_1 _10545_ (.A(_02939_),
    .B(_02940_),
    .X(_00004_));
 sg13g2_and2_1 _10546_ (.A(_02936_),
    .B(_02939_),
    .X(_02941_));
 sg13g2_o21ai_1 _10547_ (.B1(_02928_),
    .Y(_02942_),
    .A1(_02920_),
    .A2(_02929_));
 sg13g2_nand2_1 _10548_ (.Y(_02943_),
    .A(net2584),
    .B(net2134));
 sg13g2_o21ai_1 _10549_ (.B1(_02926_),
    .Y(_02944_),
    .A1(_02905_),
    .A2(_02924_));
 sg13g2_nand2_1 _10550_ (.Y(_02945_),
    .A(net2585),
    .B(net2127));
 sg13g2_nand2_1 _10551_ (.Y(_02946_),
    .A(net2586),
    .B(net2130));
 sg13g2_nand2_1 _10552_ (.Y(_02947_),
    .A(net2586),
    .B(net2136));
 sg13g2_xor2_1 _10553_ (.B(_02947_),
    .A(_02923_),
    .X(_02948_));
 sg13g2_nand2b_1 _10554_ (.Y(_02949_),
    .B(_02948_),
    .A_N(_02945_));
 sg13g2_xnor2_1 _10555_ (.Y(_02950_),
    .A(_02945_),
    .B(_02948_));
 sg13g2_nand2_1 _10556_ (.Y(_02951_),
    .A(_02944_),
    .B(_02950_));
 sg13g2_xnor2_1 _10557_ (.Y(_02952_),
    .A(_02944_),
    .B(_02950_));
 sg13g2_xor2_1 _10558_ (.B(_02952_),
    .A(_02943_),
    .X(_02953_));
 sg13g2_nand2_1 _10559_ (.Y(_02954_),
    .A(_02942_),
    .B(_02953_));
 sg13g2_xnor2_1 _10560_ (.Y(_02955_),
    .A(_02942_),
    .B(_02953_));
 sg13g2_xnor2_1 _10561_ (.Y(_02956_),
    .A(_02052_),
    .B(_02955_));
 sg13g2_o21ai_1 _10562_ (.B1(_02931_),
    .Y(_02957_),
    .A1(_02051_),
    .A2(_02932_));
 sg13g2_nor2b_1 _10563_ (.A(_02956_),
    .B_N(_02957_),
    .Y(_02958_));
 sg13g2_xnor2_1 _10564_ (.Y(_02959_),
    .A(_02956_),
    .B(_02957_));
 sg13g2_inv_1 _10565_ (.Y(_02960_),
    .A(_02959_));
 sg13g2_a21oi_2 _10566_ (.B1(_02960_),
    .Y(_02961_),
    .A2(_02939_),
    .A1(_02936_));
 sg13g2_xnor2_1 _10567_ (.Y(_00005_),
    .A(_02941_),
    .B(_02959_));
 sg13g2_nor2_1 _10568_ (.A(_02958_),
    .B(_02961_),
    .Y(_02962_));
 sg13g2_o21ai_1 _10569_ (.B1(_02951_),
    .Y(_02963_),
    .A1(_02943_),
    .A2(_02952_));
 sg13g2_nand2_1 _10570_ (.Y(_02964_),
    .A(net2583),
    .B(net2132));
 sg13g2_o21ai_1 _10571_ (.B1(_02949_),
    .Y(_02965_),
    .A1(_02923_),
    .A2(_02947_));
 sg13g2_nand2_1 _10572_ (.Y(_02966_),
    .A(net2584),
    .B(net2126));
 sg13g2_nand2_1 _10573_ (.Y(_02967_),
    .A(net2585),
    .B(net2130));
 sg13g2_nand2_1 _10574_ (.Y(_02968_),
    .A(net2585),
    .B(net2136));
 sg13g2_xor2_1 _10575_ (.B(_02968_),
    .A(_02946_),
    .X(_02969_));
 sg13g2_nand2b_1 _10576_ (.Y(_02970_),
    .B(_02969_),
    .A_N(_02966_));
 sg13g2_xnor2_1 _10577_ (.Y(_02971_),
    .A(_02966_),
    .B(_02969_));
 sg13g2_nand2_1 _10578_ (.Y(_02972_),
    .A(_02965_),
    .B(_02971_));
 sg13g2_xnor2_1 _10579_ (.Y(_02973_),
    .A(_02965_),
    .B(_02971_));
 sg13g2_xor2_1 _10580_ (.B(_02973_),
    .A(_02964_),
    .X(_02974_));
 sg13g2_nand2_1 _10581_ (.Y(_02975_),
    .A(_02963_),
    .B(_02974_));
 sg13g2_xnor2_1 _10582_ (.Y(_02976_),
    .A(_02963_),
    .B(_02974_));
 sg13g2_xnor2_1 _10583_ (.Y(_02977_),
    .A(_02053_),
    .B(_02976_));
 sg13g2_o21ai_1 _10584_ (.B1(_02954_),
    .Y(_02978_),
    .A1(_02052_),
    .A2(_02955_));
 sg13g2_nand2b_1 _10585_ (.Y(_02979_),
    .B(_02978_),
    .A_N(_02977_));
 sg13g2_xnor2_1 _10586_ (.Y(_02980_),
    .A(_02977_),
    .B(_02978_));
 sg13g2_inv_1 _10587_ (.Y(_02981_),
    .A(_02980_));
 sg13g2_xnor2_1 _10588_ (.Y(_00006_),
    .A(_02962_),
    .B(_02980_));
 sg13g2_o21ai_1 _10589_ (.B1(_02979_),
    .Y(_02982_),
    .A1(_02962_),
    .A2(_02981_));
 sg13g2_o21ai_1 _10590_ (.B1(_02975_),
    .Y(_02983_),
    .A1(_02053_),
    .A2(_02976_));
 sg13g2_o21ai_1 _10591_ (.B1(_02972_),
    .Y(_02984_),
    .A1(_02964_),
    .A2(_02973_));
 sg13g2_nand2_1 _10592_ (.Y(_02985_),
    .A(net2582),
    .B(net2132));
 sg13g2_o21ai_1 _10593_ (.B1(_02970_),
    .Y(_02986_),
    .A1(_02946_),
    .A2(_02968_));
 sg13g2_nand2_1 _10594_ (.Y(_02987_),
    .A(net2583),
    .B(net2126));
 sg13g2_nand2_1 _10595_ (.Y(_02988_),
    .A(net2584),
    .B(net2130));
 sg13g2_nand2_1 _10596_ (.Y(_02989_),
    .A(net2584),
    .B(net2135));
 sg13g2_xor2_1 _10597_ (.B(_02989_),
    .A(_02967_),
    .X(_02990_));
 sg13g2_nand2b_1 _10598_ (.Y(_02991_),
    .B(_02990_),
    .A_N(_02987_));
 sg13g2_xnor2_1 _10599_ (.Y(_02992_),
    .A(_02987_),
    .B(_02990_));
 sg13g2_nand2_1 _10600_ (.Y(_02993_),
    .A(_02986_),
    .B(_02992_));
 sg13g2_xnor2_1 _10601_ (.Y(_02994_),
    .A(_02986_),
    .B(_02992_));
 sg13g2_xor2_1 _10602_ (.B(_02994_),
    .A(_02985_),
    .X(_02995_));
 sg13g2_nand2_1 _10603_ (.Y(_02996_),
    .A(_02984_),
    .B(_02995_));
 sg13g2_xnor2_1 _10604_ (.Y(_02997_),
    .A(_02984_),
    .B(_02995_));
 sg13g2_xnor2_1 _10605_ (.Y(_02998_),
    .A(_02054_),
    .B(_02997_));
 sg13g2_nor2b_1 _10606_ (.A(_02983_),
    .B_N(_02998_),
    .Y(_02999_));
 sg13g2_nor2b_1 _10607_ (.A(_02998_),
    .B_N(_02983_),
    .Y(_03000_));
 sg13g2_or2_1 _10608_ (.X(_03001_),
    .B(_03000_),
    .A(_02999_));
 sg13g2_xnor2_1 _10609_ (.Y(_00007_),
    .A(_02982_),
    .B(_03001_));
 sg13g2_o21ai_1 _10610_ (.B1(_02993_),
    .Y(_03002_),
    .A1(_02985_),
    .A2(_02994_));
 sg13g2_nand2_1 _10611_ (.Y(_03003_),
    .A(net2581),
    .B(net2132));
 sg13g2_o21ai_1 _10612_ (.B1(_02991_),
    .Y(_03004_),
    .A1(_02967_),
    .A2(_02989_));
 sg13g2_nand2_1 _10613_ (.Y(_03005_),
    .A(net2582),
    .B(net2127));
 sg13g2_nand2_1 _10614_ (.Y(_03006_),
    .A(net2583),
    .B(net2129));
 sg13g2_nand2_1 _10615_ (.Y(_03007_),
    .A(net2583),
    .B(net2136));
 sg13g2_xor2_1 _10616_ (.B(_03007_),
    .A(_02988_),
    .X(_03008_));
 sg13g2_nand2b_1 _10617_ (.Y(_03009_),
    .B(_03008_),
    .A_N(_03005_));
 sg13g2_xnor2_1 _10618_ (.Y(_03010_),
    .A(_03005_),
    .B(_03008_));
 sg13g2_nand2_1 _10619_ (.Y(_03011_),
    .A(_03004_),
    .B(_03010_));
 sg13g2_xnor2_1 _10620_ (.Y(_03012_),
    .A(_03004_),
    .B(_03010_));
 sg13g2_xor2_1 _10621_ (.B(_03012_),
    .A(_03003_),
    .X(_03013_));
 sg13g2_nand2_1 _10622_ (.Y(_03014_),
    .A(_03002_),
    .B(_03013_));
 sg13g2_xnor2_1 _10623_ (.Y(_03015_),
    .A(_03002_),
    .B(_03013_));
 sg13g2_xnor2_1 _10624_ (.Y(_03016_),
    .A(_02055_),
    .B(_03015_));
 sg13g2_o21ai_1 _10625_ (.B1(_02996_),
    .Y(_03017_),
    .A1(_02054_),
    .A2(_02997_));
 sg13g2_nor2b_1 _10626_ (.A(_03016_),
    .B_N(_03017_),
    .Y(_03018_));
 sg13g2_nand2b_1 _10627_ (.Y(_03019_),
    .B(_03017_),
    .A_N(_03016_));
 sg13g2_xnor2_1 _10628_ (.Y(_03020_),
    .A(_03016_),
    .B(_03017_));
 sg13g2_nor2_1 _10629_ (.A(_02981_),
    .B(_03001_),
    .Y(_03021_));
 sg13g2_o21ai_1 _10630_ (.B1(_03021_),
    .Y(_03022_),
    .A1(_02958_),
    .A2(_02961_));
 sg13g2_nor2_1 _10631_ (.A(_02979_),
    .B(_02999_),
    .Y(_03023_));
 sg13g2_nor2_1 _10632_ (.A(_03000_),
    .B(_03023_),
    .Y(_03024_));
 sg13g2_nand2_1 _10633_ (.Y(_03025_),
    .A(_03022_),
    .B(_03024_));
 sg13g2_xor2_1 _10634_ (.B(_03025_),
    .A(_03020_),
    .X(_00008_));
 sg13g2_o21ai_1 _10635_ (.B1(_03014_),
    .Y(_03026_),
    .A1(_02055_),
    .A2(_03015_));
 sg13g2_o21ai_1 _10636_ (.B1(_03011_),
    .Y(_03027_),
    .A1(_03003_),
    .A2(_03012_));
 sg13g2_nand2_1 _10637_ (.Y(_03028_),
    .A(net2580),
    .B(net2132));
 sg13g2_o21ai_1 _10638_ (.B1(_03009_),
    .Y(_03029_),
    .A1(_02988_),
    .A2(_03007_));
 sg13g2_nand2_1 _10639_ (.Y(_03030_),
    .A(net2581),
    .B(net2126));
 sg13g2_nand2_1 _10640_ (.Y(_03031_),
    .A(net2582),
    .B(net2129));
 sg13g2_nand2_1 _10641_ (.Y(_03032_),
    .A(net2582),
    .B(net2135));
 sg13g2_xor2_1 _10642_ (.B(_03032_),
    .A(_03006_),
    .X(_03033_));
 sg13g2_nand2b_1 _10643_ (.Y(_03034_),
    .B(_03033_),
    .A_N(_03030_));
 sg13g2_xnor2_1 _10644_ (.Y(_03035_),
    .A(_03030_),
    .B(_03033_));
 sg13g2_nand2_1 _10645_ (.Y(_03036_),
    .A(_03029_),
    .B(_03035_));
 sg13g2_xnor2_1 _10646_ (.Y(_03037_),
    .A(_03029_),
    .B(_03035_));
 sg13g2_xor2_1 _10647_ (.B(_03037_),
    .A(_03028_),
    .X(_03038_));
 sg13g2_nand2_1 _10648_ (.Y(_03039_),
    .A(_03027_),
    .B(_03038_));
 sg13g2_xnor2_1 _10649_ (.Y(_03040_),
    .A(_03027_),
    .B(_03038_));
 sg13g2_xnor2_1 _10650_ (.Y(_03041_),
    .A(_02056_),
    .B(_03040_));
 sg13g2_nor2b_1 _10651_ (.A(_03026_),
    .B_N(_03041_),
    .Y(_03042_));
 sg13g2_nand2b_1 _10652_ (.Y(_03043_),
    .B(_03026_),
    .A_N(_03041_));
 sg13g2_nand2b_1 _10653_ (.Y(_03044_),
    .B(_03043_),
    .A_N(_03042_));
 sg13g2_a21o_1 _10654_ (.A2(_03025_),
    .A1(_03020_),
    .B1(_03018_),
    .X(_03045_));
 sg13g2_xnor2_1 _10655_ (.Y(_00009_),
    .A(_03044_),
    .B(_03045_));
 sg13g2_o21ai_1 _10656_ (.B1(_03036_),
    .Y(_03046_),
    .A1(_03028_),
    .A2(_03037_));
 sg13g2_nand2_1 _10657_ (.Y(_03047_),
    .A(net2579),
    .B(net2132));
 sg13g2_o21ai_1 _10658_ (.B1(_03034_),
    .Y(_03048_),
    .A1(_03006_),
    .A2(_03032_));
 sg13g2_nand2_1 _10659_ (.Y(_03049_),
    .A(net2580),
    .B(net2126));
 sg13g2_nand2_1 _10660_ (.Y(_03050_),
    .A(net2581),
    .B(net2129));
 sg13g2_nand2_1 _10661_ (.Y(_03051_),
    .A(net2581),
    .B(net2135));
 sg13g2_xor2_1 _10662_ (.B(_03051_),
    .A(_03031_),
    .X(_03052_));
 sg13g2_nand2b_1 _10663_ (.Y(_03053_),
    .B(_03052_),
    .A_N(_03049_));
 sg13g2_xnor2_1 _10664_ (.Y(_03054_),
    .A(_03049_),
    .B(_03052_));
 sg13g2_nand2_1 _10665_ (.Y(_03055_),
    .A(_03048_),
    .B(_03054_));
 sg13g2_xnor2_1 _10666_ (.Y(_03056_),
    .A(_03048_),
    .B(_03054_));
 sg13g2_xor2_1 _10667_ (.B(_03056_),
    .A(_03047_),
    .X(_03057_));
 sg13g2_nand2_1 _10668_ (.Y(_03058_),
    .A(_03046_),
    .B(_03057_));
 sg13g2_xnor2_1 _10669_ (.Y(_03059_),
    .A(_03046_),
    .B(_03057_));
 sg13g2_xnor2_1 _10670_ (.Y(_03060_),
    .A(_02057_),
    .B(_03059_));
 sg13g2_o21ai_1 _10671_ (.B1(_03039_),
    .Y(_03061_),
    .A1(_02056_),
    .A2(_03040_));
 sg13g2_nor2b_1 _10672_ (.A(_03060_),
    .B_N(_03061_),
    .Y(_03062_));
 sg13g2_inv_1 _10673_ (.Y(_03063_),
    .A(_03062_));
 sg13g2_xnor2_1 _10674_ (.Y(_03064_),
    .A(_03060_),
    .B(_03061_));
 sg13g2_nand3b_1 _10675_ (.B(_03043_),
    .C(_03020_),
    .Y(_03065_),
    .A_N(_03042_));
 sg13g2_a21oi_1 _10676_ (.A1(_03022_),
    .A2(_03024_),
    .Y(_03066_),
    .B1(_03065_));
 sg13g2_o21ai_1 _10677_ (.B1(_03043_),
    .Y(_03067_),
    .A1(_03019_),
    .A2(_03042_));
 sg13g2_nor2_1 _10678_ (.A(_03066_),
    .B(_03067_),
    .Y(_03068_));
 sg13g2_o21ai_1 _10679_ (.B1(_03064_),
    .Y(_03069_),
    .A1(_03066_),
    .A2(_03067_));
 sg13g2_xnor2_1 _10680_ (.Y(_00010_),
    .A(_03064_),
    .B(_03068_));
 sg13g2_o21ai_1 _10681_ (.B1(_03055_),
    .Y(_03070_),
    .A1(_03047_),
    .A2(_03056_));
 sg13g2_nand2_1 _10682_ (.Y(_03071_),
    .A(net2578),
    .B(net2132));
 sg13g2_o21ai_1 _10683_ (.B1(_03053_),
    .Y(_03072_),
    .A1(_03031_),
    .A2(_03051_));
 sg13g2_nand2_1 _10684_ (.Y(_03073_),
    .A(net2579),
    .B(net2126));
 sg13g2_nand2_1 _10685_ (.Y(_03074_),
    .A(net2580),
    .B(net2129));
 sg13g2_nand2_1 _10686_ (.Y(_03075_),
    .A(net2580),
    .B(net2135));
 sg13g2_xor2_1 _10687_ (.B(_03075_),
    .A(_03050_),
    .X(_03076_));
 sg13g2_nand2b_1 _10688_ (.Y(_03077_),
    .B(_03076_),
    .A_N(_03073_));
 sg13g2_xnor2_1 _10689_ (.Y(_03078_),
    .A(_03073_),
    .B(_03076_));
 sg13g2_nand2_1 _10690_ (.Y(_03079_),
    .A(_03072_),
    .B(_03078_));
 sg13g2_xnor2_1 _10691_ (.Y(_03080_),
    .A(_03072_),
    .B(_03078_));
 sg13g2_xor2_1 _10692_ (.B(_03080_),
    .A(_03071_),
    .X(_03081_));
 sg13g2_nand2_1 _10693_ (.Y(_03082_),
    .A(_03070_),
    .B(_03081_));
 sg13g2_xnor2_1 _10694_ (.Y(_03083_),
    .A(_03070_),
    .B(_03081_));
 sg13g2_xnor2_1 _10695_ (.Y(_03084_),
    .A(_02058_),
    .B(_03083_));
 sg13g2_o21ai_1 _10696_ (.B1(_03058_),
    .Y(_03085_),
    .A1(_02057_),
    .A2(_03059_));
 sg13g2_nor2b_1 _10697_ (.A(_03084_),
    .B_N(_03085_),
    .Y(_03086_));
 sg13g2_xnor2_1 _10698_ (.Y(_03087_),
    .A(_03084_),
    .B(_03085_));
 sg13g2_inv_1 _10699_ (.Y(_03088_),
    .A(_03087_));
 sg13g2_a21oi_1 _10700_ (.A1(_03063_),
    .A2(_03069_),
    .Y(_03089_),
    .B1(_03088_));
 sg13g2_nand3_1 _10701_ (.B(_03069_),
    .C(_03088_),
    .A(_03063_),
    .Y(_03090_));
 sg13g2_nor2b_1 _10702_ (.A(_03089_),
    .B_N(_03090_),
    .Y(_00011_));
 sg13g2_o21ai_1 _10703_ (.B1(_03079_),
    .Y(_03091_),
    .A1(_03071_),
    .A2(_03080_));
 sg13g2_nand2_1 _10704_ (.Y(_03092_),
    .A(net2577),
    .B(net2132));
 sg13g2_o21ai_1 _10705_ (.B1(_03077_),
    .Y(_03093_),
    .A1(_03050_),
    .A2(_03075_));
 sg13g2_nand2_1 _10706_ (.Y(_03094_),
    .A(net2578),
    .B(net2126));
 sg13g2_nand2_2 _10707_ (.Y(_03095_),
    .A(net2579),
    .B(net2135));
 sg13g2_xor2_1 _10708_ (.B(_03095_),
    .A(_03074_),
    .X(_03096_));
 sg13g2_nand2b_1 _10709_ (.Y(_03097_),
    .B(_03096_),
    .A_N(_03094_));
 sg13g2_xnor2_1 _10710_ (.Y(_03098_),
    .A(_03094_),
    .B(_03096_));
 sg13g2_nand2_1 _10711_ (.Y(_03099_),
    .A(_03093_),
    .B(_03098_));
 sg13g2_xnor2_1 _10712_ (.Y(_03100_),
    .A(_03093_),
    .B(_03098_));
 sg13g2_xor2_1 _10713_ (.B(_03100_),
    .A(_03092_),
    .X(_03101_));
 sg13g2_nand2_1 _10714_ (.Y(_03102_),
    .A(_03091_),
    .B(_03101_));
 sg13g2_xnor2_1 _10715_ (.Y(_03103_),
    .A(_03091_),
    .B(_03101_));
 sg13g2_xnor2_1 _10716_ (.Y(_03104_),
    .A(_02059_),
    .B(_03103_));
 sg13g2_o21ai_1 _10717_ (.B1(_03082_),
    .Y(_03105_),
    .A1(_02058_),
    .A2(_03083_));
 sg13g2_nand2b_1 _10718_ (.Y(_03106_),
    .B(_03105_),
    .A_N(_03104_));
 sg13g2_xnor2_1 _10719_ (.Y(_03107_),
    .A(_03104_),
    .B(_03105_));
 sg13g2_o21ai_1 _10720_ (.B1(_03107_),
    .Y(_03108_),
    .A1(_03086_),
    .A2(_03089_));
 sg13g2_or3_1 _10721_ (.A(_03086_),
    .B(_03089_),
    .C(_03107_),
    .X(_03109_));
 sg13g2_and2_1 _10722_ (.A(_03108_),
    .B(_03109_),
    .X(_00001_));
 sg13g2_o21ai_1 _10723_ (.B1(_03099_),
    .Y(_03110_),
    .A1(_03092_),
    .A2(_03100_));
 sg13g2_nand2_1 _10724_ (.Y(_03111_),
    .A(net2576),
    .B(net2132));
 sg13g2_o21ai_1 _10725_ (.B1(_03097_),
    .Y(_03112_),
    .A1(_03074_),
    .A2(_03095_));
 sg13g2_nand2_1 _10726_ (.Y(_03113_),
    .A(net2577),
    .B(net2126));
 sg13g2_nand2_2 _10727_ (.Y(_03114_),
    .A(net2578),
    .B(net2129));
 sg13g2_nor2_1 _10728_ (.A(_03095_),
    .B(_03114_),
    .Y(_03115_));
 sg13g2_or2_1 _10729_ (.X(_03116_),
    .B(_03114_),
    .A(_03095_));
 sg13g2_a22oi_1 _10730_ (.Y(_03117_),
    .B1(net2129),
    .B2(net2579),
    .A2(net2135),
    .A1(net2578));
 sg13g2_or2_1 _10731_ (.X(_03118_),
    .B(_03117_),
    .A(_03115_));
 sg13g2_xor2_1 _10732_ (.B(_03118_),
    .A(_03113_),
    .X(_03119_));
 sg13g2_nand2_1 _10733_ (.Y(_03120_),
    .A(_03112_),
    .B(_03119_));
 sg13g2_xnor2_1 _10734_ (.Y(_03121_),
    .A(_03112_),
    .B(_03119_));
 sg13g2_xor2_1 _10735_ (.B(_03121_),
    .A(_03111_),
    .X(_03122_));
 sg13g2_nand2_1 _10736_ (.Y(_03123_),
    .A(_03110_),
    .B(_03122_));
 sg13g2_xnor2_1 _10737_ (.Y(_03124_),
    .A(_03110_),
    .B(_03122_));
 sg13g2_xnor2_1 _10738_ (.Y(_03125_),
    .A(_02060_),
    .B(_03124_));
 sg13g2_o21ai_1 _10739_ (.B1(_03102_),
    .Y(_03126_),
    .A1(_02059_),
    .A2(_03103_));
 sg13g2_nor2b_1 _10740_ (.A(_03125_),
    .B_N(_03126_),
    .Y(_03127_));
 sg13g2_xor2_1 _10741_ (.B(_03126_),
    .A(_03125_),
    .X(_03128_));
 sg13g2_a21oi_1 _10742_ (.A1(_03106_),
    .A2(_03108_),
    .Y(_03129_),
    .B1(_03128_));
 sg13g2_nand3_1 _10743_ (.B(_03108_),
    .C(_03128_),
    .A(_03106_),
    .Y(_03130_));
 sg13g2_nor2b_1 _10744_ (.A(_03129_),
    .B_N(_03130_),
    .Y(_00002_));
 sg13g2_a21oi_1 _10745_ (.A1(\i_tinyqv.mem.q_ctrl.data_ready ),
    .A2(_02763_),
    .Y(_03131_),
    .B1(\i_tinyqv.mem.qspi_write_done ));
 sg13g2_nor2_2 _10746_ (.A(net2611),
    .B(_03131_),
    .Y(_03132_));
 sg13g2_or2_1 _10747_ (.X(_03133_),
    .B(_03131_),
    .A(net2611));
 sg13g2_a22oi_1 _10748_ (.Y(_03134_),
    .B1(net2390),
    .B2(_03133_),
    .A2(_02020_),
    .A1(net2472));
 sg13g2_nor3_2 _10749_ (.A(\i_tinyqv.cpu.data_ready_latch ),
    .B(net2318),
    .C(_03134_),
    .Y(_03135_));
 sg13g2_nor2_1 _10750_ (.A(net4309),
    .B(net2320),
    .Y(_03136_));
 sg13g2_nor2_1 _10751_ (.A(_03135_),
    .B(_03136_),
    .Y(_03137_));
 sg13g2_nand3_1 _10752_ (.B(_02765_),
    .C(_03137_),
    .A(\i_tinyqv.cpu.is_load ),
    .Y(_03138_));
 sg13g2_o21ai_1 _10753_ (.B1(_02809_),
    .Y(_03139_),
    .A1(net2528),
    .A2(net2530));
 sg13g2_nand2_1 _10754_ (.Y(_03140_),
    .A(_02792_),
    .B(_03139_));
 sg13g2_nor2_1 _10755_ (.A(_02806_),
    .B(_03140_),
    .Y(_03141_));
 sg13g2_and2_1 _10756_ (.A(_02496_),
    .B(_02792_),
    .X(_03142_));
 sg13g2_nand2_1 _10757_ (.Y(_03143_),
    .A(_02496_),
    .B(_02792_));
 sg13g2_nor2_1 _10758_ (.A(_01991_),
    .B(_02796_),
    .Y(_03144_));
 sg13g2_nand2_2 _10759_ (.Y(_03145_),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .B(_02795_));
 sg13g2_nor2_1 _10760_ (.A(_03142_),
    .B(_03145_),
    .Y(_03146_));
 sg13g2_a22oi_1 _10761_ (.Y(_03147_),
    .B1(_03146_),
    .B2(_01962_),
    .A2(_03141_),
    .A1(_03138_));
 sg13g2_and2_1 _10762_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .X(_03148_));
 sg13g2_nand2_1 _10763_ (.Y(_03149_),
    .A(net2505),
    .B(_03148_));
 sg13g2_nand4_1 _10764_ (.B(net2504),
    .C(net1889),
    .A(net2505),
    .Y(_03150_),
    .D(_03148_));
 sg13g2_nand2b_2 _10765_ (.Y(_03151_),
    .B(\i_tinyqv.cpu.i_core.cycle[0] ),
    .A_N(\i_tinyqv.cpu.i_core.cycle[1] ));
 sg13g2_nor2_2 _10766_ (.A(net2365),
    .B(_03151_),
    .Y(_03152_));
 sg13g2_nor3_2 _10767_ (.A(net2527),
    .B(net2524),
    .C(net2529),
    .Y(_03153_));
 sg13g2_or3_1 _10768_ (.A(net2527),
    .B(net2525),
    .C(net2529),
    .X(_03154_));
 sg13g2_xnor2_1 _10769_ (.Y(_03155_),
    .A(_02738_),
    .B(_02742_));
 sg13g2_and3_2 _10770_ (.X(_03156_),
    .A(net2525),
    .B(_02559_),
    .C(_02794_));
 sg13g2_nor2_2 _10771_ (.A(net2434),
    .B(_02559_),
    .Y(_03157_));
 sg13g2_a21o_1 _10772_ (.A2(_02733_),
    .A1(_02713_),
    .B1(net2529),
    .X(_03158_));
 sg13g2_o21ai_1 _10773_ (.B1(_03158_),
    .Y(_03159_),
    .A1(_02713_),
    .A2(_02733_));
 sg13g2_and2_1 _10774_ (.A(_03157_),
    .B(_03159_),
    .X(_03160_));
 sg13g2_a221oi_1 _10775_ (.B2(_02774_),
    .C1(_03160_),
    .B1(_03156_),
    .A1(_03153_),
    .Y(_03161_),
    .A2(_03155_));
 sg13g2_a21oi_1 _10776_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .A2(net2134),
    .Y(_03162_),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[0] ));
 sg13g2_nand2_1 _10777_ (.Y(_03163_),
    .A(_02867_),
    .B(_03144_));
 sg13g2_o21ai_1 _10778_ (.B1(_03161_),
    .Y(_03164_),
    .A1(_03162_),
    .A2(_03163_));
 sg13g2_nor4_1 _10779_ (.A(\i_tinyqv.cpu.alu_op[3] ),
    .B(net2319),
    .C(_02796_),
    .D(_03151_),
    .Y(_03165_));
 sg13g2_nor2_1 _10780_ (.A(_02794_),
    .B(_03151_),
    .Y(_03166_));
 sg13g2_or2_1 _10781_ (.X(_03167_),
    .B(_03151_),
    .A(_02794_));
 sg13g2_nand2_1 _10782_ (.Y(_03168_),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sg13g2_xnor2_1 _10783_ (.Y(_03169_),
    .A(net2533),
    .B(net2522));
 sg13g2_nor2_1 _10784_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_03169_),
    .Y(_03170_));
 sg13g2_nand2_1 _10785_ (.Y(_03171_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_03169_));
 sg13g2_xor2_1 _10786_ (.B(net2524),
    .A(\i_tinyqv.cpu.counter[3] ),
    .X(_03172_));
 sg13g2_nor2b_1 _10787_ (.A(_03172_),
    .B_N(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .Y(_03173_));
 sg13g2_xnor2_1 _10788_ (.Y(_03174_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .B(_03172_));
 sg13g2_xnor2_1 _10789_ (.Y(_03175_),
    .A(net2540),
    .B(net2522));
 sg13g2_and2_1 _10790_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_03175_),
    .X(_03176_));
 sg13g2_a21oi_1 _10791_ (.A1(_03174_),
    .A2(_03176_),
    .Y(_03177_),
    .B1(_03173_));
 sg13g2_o21ai_1 _10792_ (.B1(_03171_),
    .Y(_03178_),
    .A1(_03170_),
    .A2(_03177_));
 sg13g2_and2_1 _10793_ (.A(_03168_),
    .B(_03178_),
    .X(_03179_));
 sg13g2_nor2_1 _10794_ (.A(net2518),
    .B(net2581),
    .Y(_03180_));
 sg13g2_nand2b_1 _10795_ (.Y(_03181_),
    .B(net2526),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[21] ));
 sg13g2_nor2b_1 _10796_ (.A(_03180_),
    .B_N(_03181_),
    .Y(_03182_));
 sg13g2_nand2b_1 _10797_ (.Y(_03183_),
    .B(_03181_),
    .A_N(_03180_));
 sg13g2_mux2_1 _10798_ (.A0(net2582),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(net2518),
    .X(_03184_));
 sg13g2_inv_1 _10799_ (.Y(_03185_),
    .A(_03184_));
 sg13g2_xor2_1 _10800_ (.B(_03175_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .X(_03186_));
 sg13g2_xnor2_1 _10801_ (.Y(_03187_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_03175_));
 sg13g2_or2_1 _10802_ (.X(_03188_),
    .B(net2579),
    .A(net2518));
 sg13g2_o21ai_1 _10803_ (.B1(_03188_),
    .Y(_03189_),
    .A1(net2432),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[19] ));
 sg13g2_or2_1 _10804_ (.X(_03190_),
    .B(net2580),
    .A(net2519));
 sg13g2_o21ai_1 _10805_ (.B1(_03190_),
    .Y(_03191_),
    .A1(net2432),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[20] ));
 sg13g2_mux4_1 _10806_ (.S0(net2477),
    .A0(_03183_),
    .A1(_03185_),
    .A2(_03189_),
    .A3(_03191_),
    .S1(net2407),
    .X(_03192_));
 sg13g2_nand2b_1 _10807_ (.Y(_03193_),
    .B(_03171_),
    .A_N(_03170_));
 sg13g2_and2_1 _10808_ (.A(_03177_),
    .B(_03193_),
    .X(_03194_));
 sg13g2_nand2_2 _10809_ (.Y(_03195_),
    .A(_03177_),
    .B(_03193_));
 sg13g2_or2_1 _10810_ (.X(_03196_),
    .B(net2583),
    .A(net2518));
 sg13g2_o21ai_1 _10811_ (.B1(_03196_),
    .Y(_03197_),
    .A1(net2432),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[23] ));
 sg13g2_inv_1 _10812_ (.Y(_03198_),
    .A(_03197_));
 sg13g2_mux2_1 _10813_ (.A0(net2584),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(net2518),
    .X(_03199_));
 sg13g2_mux2_1 _10814_ (.A0(net2585),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S(net2519),
    .X(_03200_));
 sg13g2_mux2_1 _10815_ (.A0(net2586),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(net2519),
    .X(_03201_));
 sg13g2_nand2b_1 _10816_ (.Y(_03202_),
    .B(net2483),
    .A_N(_03201_));
 sg13g2_or2_1 _10817_ (.X(_03203_),
    .B(_03200_),
    .A(net2481));
 sg13g2_mux4_1 _10818_ (.S0(net2478),
    .A0(_03198_),
    .A1(_03199_),
    .A2(_03200_),
    .A3(_03201_),
    .S1(net2474),
    .X(_03204_));
 sg13g2_a21oi_1 _10819_ (.A1(net2313),
    .A2(_03204_),
    .Y(_03205_),
    .B1(net2178));
 sg13g2_o21ai_1 _10820_ (.B1(_03205_),
    .Y(_03206_),
    .A1(net2313),
    .A2(_03192_));
 sg13g2_or2_1 _10821_ (.X(_03207_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A(net2519));
 sg13g2_o21ai_1 _10822_ (.B1(_03207_),
    .Y(_03208_),
    .A1(net2432),
    .A2(net2584));
 sg13g2_mux2_1 _10823_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(net2583),
    .S(net2518),
    .X(_03209_));
 sg13g2_nand2_1 _10824_ (.Y(_03210_),
    .A(net2481),
    .B(_03209_));
 sg13g2_o21ai_1 _10825_ (.B1(_03210_),
    .Y(_03211_),
    .A1(net2481),
    .A2(_03208_));
 sg13g2_or2_1 _10826_ (.X(_03212_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A(net2518));
 sg13g2_o21ai_1 _10827_ (.B1(_03212_),
    .Y(_03213_),
    .A1(net2432),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[9] ));
 sg13g2_nor2_1 _10828_ (.A(net2479),
    .B(_03213_),
    .Y(_03214_));
 sg13g2_mux2_1 _10829_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .S(net2518),
    .X(_03215_));
 sg13g2_a21oi_1 _10830_ (.A1(net2479),
    .A2(_03215_),
    .Y(_03216_),
    .B1(_03214_));
 sg13g2_a21oi_1 _10831_ (.A1(net2473),
    .A2(_03216_),
    .Y(_03217_),
    .B1(net2311));
 sg13g2_o21ai_1 _10832_ (.B1(_03217_),
    .Y(_03218_),
    .A1(net2473),
    .A2(_03211_));
 sg13g2_or2_1 _10833_ (.X(_03219_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A(net2523));
 sg13g2_o21ai_1 _10834_ (.B1(_03219_),
    .Y(_03220_),
    .A1(net2433),
    .A2(net2586));
 sg13g2_nor2_1 _10835_ (.A(net2483),
    .B(_03220_),
    .Y(_03221_));
 sg13g2_mux2_1 _10836_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(net2585),
    .S(net2523),
    .X(_03222_));
 sg13g2_a21oi_1 _10837_ (.A1(net2483),
    .A2(_03222_),
    .Y(_03223_),
    .B1(_03221_));
 sg13g2_nand2_1 _10838_ (.Y(_03224_),
    .A(net2475),
    .B(_03223_));
 sg13g2_mux2_1 _10839_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .S(net2523),
    .X(_03225_));
 sg13g2_nor2b_1 _10840_ (.A(net2484),
    .B_N(_03225_),
    .Y(_03226_));
 sg13g2_mux2_1 _10841_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(net2587),
    .S(net2523),
    .X(_03227_));
 sg13g2_a21oi_1 _10842_ (.A1(net2484),
    .A2(_03227_),
    .Y(_03228_),
    .B1(_03226_));
 sg13g2_a21oi_1 _10843_ (.A1(net2408),
    .A2(_03228_),
    .Y(_03229_),
    .B1(net2314));
 sg13g2_nand2_1 _10844_ (.Y(_03230_),
    .A(_03224_),
    .B(_03229_));
 sg13g2_nand3_1 _10845_ (.B(_03218_),
    .C(_03230_),
    .A(net2178),
    .Y(_03231_));
 sg13g2_xnor2_1 _10846_ (.Y(_03232_),
    .A(_03174_),
    .B(_03176_));
 sg13g2_nand3_1 _10847_ (.B(_03231_),
    .C(_03232_),
    .A(_03206_),
    .Y(_03233_));
 sg13g2_or2_1 _10848_ (.X(_03234_),
    .B(net2587),
    .A(net2521));
 sg13g2_o21ai_1 _10849_ (.B1(_03234_),
    .Y(_03235_),
    .A1(net2433),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[27] ));
 sg13g2_mux2_1 _10850_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .S(net2523),
    .X(_03236_));
 sg13g2_nand2_1 _10851_ (.Y(_03237_),
    .A(net2485),
    .B(_03236_));
 sg13g2_o21ai_1 _10852_ (.B1(_03237_),
    .Y(_03238_),
    .A1(net2485),
    .A2(_03235_));
 sg13g2_or2_1 _10853_ (.X(_03239_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .A(net2521));
 sg13g2_o21ai_1 _10854_ (.B1(_03239_),
    .Y(_03240_),
    .A1(net2433),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[29] ));
 sg13g2_nand2_1 _10855_ (.Y(_03241_),
    .A(net2521),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[30] ));
 sg13g2_o21ai_1 _10856_ (.B1(_03241_),
    .Y(_03242_),
    .A1(net2521),
    .A2(_02047_));
 sg13g2_nand2_1 _10857_ (.Y(_03243_),
    .A(net2485),
    .B(_03242_));
 sg13g2_o21ai_1 _10858_ (.B1(_03243_),
    .Y(_03244_),
    .A1(net2485),
    .A2(_03240_));
 sg13g2_mux2_1 _10859_ (.A0(_03238_),
    .A1(_03244_),
    .S(net2476),
    .X(_03245_));
 sg13g2_nand2_1 _10860_ (.Y(_03246_),
    .A(net2521),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sg13g2_o21ai_1 _10861_ (.B1(_03246_),
    .Y(_03247_),
    .A1(net2522),
    .A2(_02048_));
 sg13g2_nor2_1 _10862_ (.A(net2486),
    .B(_03247_),
    .Y(_03248_));
 sg13g2_a21oi_1 _10863_ (.A1(net2486),
    .A2(_03168_),
    .Y(_03249_),
    .B1(_03248_));
 sg13g2_a21oi_1 _10864_ (.A1(net2476),
    .A2(_03168_),
    .Y(_03250_),
    .B1(net2312));
 sg13g2_o21ai_1 _10865_ (.B1(_03250_),
    .Y(_03251_),
    .A1(net2476),
    .A2(_03249_));
 sg13g2_a21oi_1 _10866_ (.A1(net2312),
    .A2(_03245_),
    .Y(_03252_),
    .B1(net2178));
 sg13g2_or2_1 _10867_ (.X(_03253_),
    .B(net2577),
    .A(net2519));
 sg13g2_o21ai_1 _10868_ (.B1(_03253_),
    .Y(_03254_),
    .A1(net2432),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sg13g2_mux2_1 _10869_ (.A0(net2578),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(net2520),
    .X(_03255_));
 sg13g2_inv_1 _10870_ (.Y(_03256_),
    .A(_03255_));
 sg13g2_nand2_1 _10871_ (.Y(_03257_),
    .A(net2479),
    .B(_03255_));
 sg13g2_o21ai_1 _10872_ (.B1(_03257_),
    .Y(_03258_),
    .A1(net2479),
    .A2(_03254_));
 sg13g2_mux2_1 _10873_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(net2576),
    .S(net2520),
    .X(_03259_));
 sg13g2_nor2b_1 _10874_ (.A(net2482),
    .B_N(_03259_),
    .Y(_03260_));
 sg13g2_mux2_1 _10875_ (.A0(net2576),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net2520),
    .X(_03261_));
 sg13g2_a21oi_1 _10876_ (.A1(net2481),
    .A2(_03261_),
    .Y(_03262_),
    .B1(_03260_));
 sg13g2_nand2_1 _10877_ (.Y(_03263_),
    .A(net2406),
    .B(_03262_));
 sg13g2_o21ai_1 _10878_ (.B1(_03263_),
    .Y(_03264_),
    .A1(net2406),
    .A2(_03258_));
 sg13g2_or2_1 _10879_ (.X(_03265_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A(net2520));
 sg13g2_o21ai_1 _10880_ (.B1(_03265_),
    .Y(_03266_),
    .A1(net2432),
    .A2(net2578));
 sg13g2_nor2_1 _10881_ (.A(net2481),
    .B(_03266_),
    .Y(_03267_));
 sg13g2_mux2_1 _10882_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .S(net2520),
    .X(_03268_));
 sg13g2_a21oi_1 _10883_ (.A1(net2482),
    .A2(_03268_),
    .Y(_03269_),
    .B1(_03267_));
 sg13g2_or2_1 _10884_ (.X(_03270_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A(net2520));
 sg13g2_o21ai_1 _10885_ (.B1(_03270_),
    .Y(_03271_),
    .A1(net2432),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[11] ));
 sg13g2_mux2_1 _10886_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .S(net2520),
    .X(_03272_));
 sg13g2_nand2_1 _10887_ (.Y(_03273_),
    .A(net2480),
    .B(_03272_));
 sg13g2_o21ai_1 _10888_ (.B1(_03273_),
    .Y(_03274_),
    .A1(net2481),
    .A2(_03271_));
 sg13g2_o21ai_1 _10889_ (.B1(net2311),
    .Y(_03275_),
    .A1(net2474),
    .A2(_03274_));
 sg13g2_a21oi_1 _10890_ (.A1(net2473),
    .A2(_03269_),
    .Y(_03276_),
    .B1(_03275_));
 sg13g2_nor2_1 _10891_ (.A(_03195_),
    .B(_03276_),
    .Y(_03277_));
 sg13g2_o21ai_1 _10892_ (.B1(_03277_),
    .Y(_03278_),
    .A1(net2312),
    .A2(_03264_));
 sg13g2_a21oi_1 _10893_ (.A1(_03251_),
    .A2(_03252_),
    .Y(_03279_),
    .B1(_03232_));
 sg13g2_a21oi_1 _10894_ (.A1(_03278_),
    .A2(_03279_),
    .Y(_03280_),
    .B1(_03178_));
 sg13g2_a21oi_1 _10895_ (.A1(_03233_),
    .A2(_03280_),
    .Y(_03281_),
    .B1(_03179_));
 sg13g2_mux2_1 _10896_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .S(net2523),
    .X(_03282_));
 sg13g2_mux2_1 _10897_ (.A0(_03282_),
    .A1(_03225_),
    .S(net2484),
    .X(_03283_));
 sg13g2_nor2_1 _10898_ (.A(net2408),
    .B(_03283_),
    .Y(_03284_));
 sg13g2_nor2_1 _10899_ (.A(net2521),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .Y(_03285_));
 sg13g2_a21oi_1 _10900_ (.A1(net2521),
    .A2(_02047_),
    .Y(_03286_),
    .B1(_03285_));
 sg13g2_nor2_1 _10901_ (.A(net2522),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .Y(_03287_));
 sg13g2_a21oi_1 _10902_ (.A1(net2522),
    .A2(_02048_),
    .Y(_03288_),
    .B1(_03287_));
 sg13g2_nand2b_1 _10903_ (.Y(_03289_),
    .B(_03288_),
    .A_N(net2486));
 sg13g2_a21oi_1 _10904_ (.A1(net2485),
    .A2(_03286_),
    .Y(_03290_),
    .B1(net2476));
 sg13g2_a21oi_1 _10905_ (.A1(_03289_),
    .A2(_03290_),
    .Y(_03291_),
    .B1(_03284_));
 sg13g2_nor2_1 _10906_ (.A(net2483),
    .B(_03227_),
    .Y(_03292_));
 sg13g2_a21oi_1 _10907_ (.A1(net2484),
    .A2(_03220_),
    .Y(_03293_),
    .B1(_03292_));
 sg13g2_nor2_1 _10908_ (.A(net2483),
    .B(_03222_),
    .Y(_03294_));
 sg13g2_a21oi_1 _10909_ (.A1(net2483),
    .A2(_03208_),
    .Y(_03295_),
    .B1(_03294_));
 sg13g2_inv_1 _10910_ (.Y(_03296_),
    .A(_03295_));
 sg13g2_a21oi_1 _10911_ (.A1(net2475),
    .A2(_03296_),
    .Y(_03297_),
    .B1(net2312));
 sg13g2_o21ai_1 _10912_ (.B1(_03297_),
    .Y(_03298_),
    .A1(net2475),
    .A2(_03293_));
 sg13g2_nor2_1 _10913_ (.A(net2479),
    .B(_03215_),
    .Y(_03299_));
 sg13g2_a21oi_1 _10914_ (.A1(net2479),
    .A2(_03271_),
    .Y(_03300_),
    .B1(_03299_));
 sg13g2_inv_1 _10915_ (.Y(_03301_),
    .A(_03300_));
 sg13g2_nor2_1 _10916_ (.A(net2478),
    .B(_03209_),
    .Y(_03302_));
 sg13g2_a21oi_1 _10917_ (.A1(net2478),
    .A2(_03213_),
    .Y(_03303_),
    .B1(_03302_));
 sg13g2_a21oi_1 _10918_ (.A1(net2473),
    .A2(_03301_),
    .Y(_03304_),
    .B1(net2313));
 sg13g2_o21ai_1 _10919_ (.B1(_03304_),
    .Y(_03305_),
    .A1(net2473),
    .A2(_03303_));
 sg13g2_mux2_1 _10920_ (.A0(_03268_),
    .A1(_03259_),
    .S(net2479),
    .X(_03306_));
 sg13g2_inv_1 _10921_ (.Y(_03307_),
    .A(_03306_));
 sg13g2_nor2_1 _10922_ (.A(net2480),
    .B(_03272_),
    .Y(_03308_));
 sg13g2_a21oi_1 _10923_ (.A1(net2481),
    .A2(_03266_),
    .Y(_03309_),
    .B1(_03308_));
 sg13g2_a21oi_1 _10924_ (.A1(net2474),
    .A2(_03307_),
    .Y(_03310_),
    .B1(net2311));
 sg13g2_o21ai_1 _10925_ (.B1(_03310_),
    .Y(_03311_),
    .A1(net2473),
    .A2(_03309_));
 sg13g2_nor2_1 _10926_ (.A(net2483),
    .B(_03201_),
    .Y(_03312_));
 sg13g2_a21oi_1 _10927_ (.A1(net2484),
    .A2(_03235_),
    .Y(_03313_),
    .B1(_03312_));
 sg13g2_mux2_1 _10928_ (.A0(_03199_),
    .A1(_03200_),
    .S(net2478),
    .X(_03314_));
 sg13g2_nor2_1 _10929_ (.A(net2473),
    .B(_03314_),
    .Y(_03315_));
 sg13g2_nor2_1 _10930_ (.A(net2313),
    .B(_03315_),
    .Y(_03316_));
 sg13g2_o21ai_1 _10931_ (.B1(_03316_),
    .Y(_03317_),
    .A1(net2408),
    .A2(_03313_));
 sg13g2_mux2_1 _10932_ (.A0(_03242_),
    .A1(_03247_),
    .S(net2486),
    .X(_03318_));
 sg13g2_nor2_1 _10933_ (.A(net2485),
    .B(_03236_),
    .Y(_03319_));
 sg13g2_a21oi_1 _10934_ (.A1(net2485),
    .A2(_03240_),
    .Y(_03320_),
    .B1(_03319_));
 sg13g2_mux2_1 _10935_ (.A0(_03318_),
    .A1(_03320_),
    .S(net2408),
    .X(_03321_));
 sg13g2_nand2_1 _10936_ (.Y(_03322_),
    .A(net2477),
    .B(_03182_));
 sg13g2_o21ai_1 _10937_ (.B1(_03322_),
    .Y(_03323_),
    .A1(net2477),
    .A2(_03191_));
 sg13g2_nor2_1 _10938_ (.A(net2477),
    .B(_03184_),
    .Y(_03324_));
 sg13g2_a21oi_1 _10939_ (.A1(net2477),
    .A2(_03197_),
    .Y(_03325_),
    .B1(_03324_));
 sg13g2_nor2_1 _10940_ (.A(net2477),
    .B(_03255_),
    .Y(_03326_));
 sg13g2_a21oi_1 _10941_ (.A1(net2478),
    .A2(_03189_),
    .Y(_03327_),
    .B1(_03326_));
 sg13g2_nor2_1 _10942_ (.A(net2479),
    .B(_03261_),
    .Y(_03328_));
 sg13g2_a21oi_1 _10943_ (.A1(net2481),
    .A2(_03254_),
    .Y(_03329_),
    .B1(_03328_));
 sg13g2_mux4_1 _10944_ (.S0(net2474),
    .A0(_03323_),
    .A1(_03325_),
    .A2(_03329_),
    .A3(_03327_),
    .S1(net2311),
    .X(_03330_));
 sg13g2_a21oi_1 _10945_ (.A1(net2312),
    .A2(_03291_),
    .Y(_03331_),
    .B1(_03195_));
 sg13g2_nor2_1 _10946_ (.A(net2178),
    .B(_03330_),
    .Y(_03332_));
 sg13g2_a21oi_1 _10947_ (.A1(_03298_),
    .A2(_03331_),
    .Y(_03333_),
    .B1(_03332_));
 sg13g2_nand3_1 _10948_ (.B(_03305_),
    .C(_03311_),
    .A(net2178),
    .Y(_03334_));
 sg13g2_a21oi_1 _10949_ (.A1(net2314),
    .A2(_03321_),
    .Y(_03335_),
    .B1(_03194_));
 sg13g2_a21oi_1 _10950_ (.A1(_03317_),
    .A2(_03335_),
    .Y(_03336_),
    .B1(_03232_));
 sg13g2_a221oi_1 _10951_ (.B2(_03336_),
    .C1(_03178_),
    .B1(_03334_),
    .A1(_03232_),
    .Y(_03337_),
    .A2(_03333_));
 sg13g2_nor3_1 _10952_ (.A(net2433),
    .B(_03179_),
    .C(_03337_),
    .Y(_03338_));
 sg13g2_a21oi_1 _10953_ (.A1(net2433),
    .A2(_03281_),
    .Y(_03339_),
    .B1(_03338_));
 sg13g2_nor2_1 _10954_ (.A(_03167_),
    .B(_03339_),
    .Y(_03340_));
 sg13g2_or3_1 _10955_ (.A(_03164_),
    .B(_03165_),
    .C(_03340_),
    .X(_03341_));
 sg13g2_nor2_2 _10956_ (.A(_02554_),
    .B(_03165_),
    .Y(_03342_));
 sg13g2_a21o_1 _10957_ (.A2(net2365),
    .A1(\i_tinyqv.cpu.i_core.cmp ),
    .B1(_03342_),
    .X(_03343_));
 sg13g2_a22oi_1 _10958_ (.Y(_03344_),
    .B1(_03341_),
    .B2(_03343_),
    .A2(_03152_),
    .A1(net2589));
 sg13g2_nand2_1 _10959_ (.Y(_03345_),
    .A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ));
 sg13g2_xnor2_1 _10960_ (.Y(_03346_),
    .A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ));
 sg13g2_nand2_1 _10961_ (.Y(_03347_),
    .A(\i_tinyqv.cpu.instr_len[1] ),
    .B(\i_tinyqv.cpu.pc[1] ));
 sg13g2_o21ai_1 _10962_ (.B1(_03345_),
    .Y(_03348_),
    .A1(_03346_),
    .A2(_03347_));
 sg13g2_nand3_1 _10963_ (.B(net2574),
    .C(_03348_),
    .A(net2573),
    .Y(_03349_));
 sg13g2_nand4_1 _10964_ (.B(net2573),
    .C(net2575),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .Y(_03350_),
    .D(_03348_));
 sg13g2_nor2_1 _10965_ (.A(_01977_),
    .B(_03350_),
    .Y(_03351_));
 sg13g2_nand3_1 _10966_ (.B(net2572),
    .C(_03351_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .Y(_03352_));
 sg13g2_nor2_1 _10967_ (.A(_01975_),
    .B(_03352_),
    .Y(_03353_));
 sg13g2_nand3_1 _10968_ (.B(net2571),
    .C(_03353_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .Y(_03354_));
 sg13g2_nor2_1 _10969_ (.A(_01974_),
    .B(_03354_),
    .Y(_03355_));
 sg13g2_nand3_1 _10970_ (.B(net2569),
    .C(_03355_),
    .A(net2568),
    .Y(_03356_));
 sg13g2_nor2_1 _10971_ (.A(_01972_),
    .B(_03356_),
    .Y(_03357_));
 sg13g2_nand3_1 _10972_ (.B(net2567),
    .C(_03357_),
    .A(\i_tinyqv.cpu.instr_data_start[17] ),
    .Y(_03358_));
 sg13g2_nor2_1 _10973_ (.A(_01971_),
    .B(_03358_),
    .Y(_03359_));
 sg13g2_nand3_1 _10974_ (.B(\i_tinyqv.cpu.instr_data_start[19] ),
    .C(_03359_),
    .A(\i_tinyqv.cpu.instr_data_start[20] ),
    .Y(_03360_));
 sg13g2_a21o_1 _10975_ (.A2(_03359_),
    .A1(net2565),
    .B1(\i_tinyqv.cpu.instr_data_start[20] ),
    .X(_03361_));
 sg13g2_nand2_1 _10976_ (.Y(_03362_),
    .A(_03360_),
    .B(_03361_));
 sg13g2_xor2_1 _10977_ (.B(_03357_),
    .A(net2567),
    .X(_03363_));
 sg13g2_a21o_1 _10978_ (.A2(_03348_),
    .A1(net2575),
    .B1(net2573),
    .X(_03364_));
 sg13g2_and2_1 _10979_ (.A(_03349_),
    .B(_03364_),
    .X(_03365_));
 sg13g2_a21o_1 _10980_ (.A2(_03351_),
    .A1(net2572),
    .B1(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(_03366_));
 sg13g2_and2_1 _10981_ (.A(_03352_),
    .B(_03366_),
    .X(_03367_));
 sg13g2_a22oi_1 _10982_ (.Y(_03368_),
    .B1(_03367_),
    .B2(net2382),
    .A2(_03365_),
    .A1(net2368));
 sg13g2_xnor2_1 _10983_ (.Y(_03369_),
    .A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(_03354_));
 sg13g2_nor2_1 _10984_ (.A(net2533),
    .B(_03368_),
    .Y(_03370_));
 sg13g2_a221oi_1 _10985_ (.B2(_02705_),
    .C1(_03370_),
    .B1(_03369_),
    .A1(net2323),
    .Y(_03371_),
    .A2(_03363_));
 sg13g2_o21ai_1 _10986_ (.B1(_03371_),
    .Y(_03372_),
    .A1(_02551_),
    .A2(_03362_));
 sg13g2_nor3_2 _10987_ (.A(\i_tinyqv.cpu.is_jal ),
    .B(\i_tinyqv.cpu.is_jalr ),
    .C(_03139_),
    .Y(_03373_));
 sg13g2_nand2_2 _10988_ (.Y(_03374_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_nor3_1 _10989_ (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .B(net2531),
    .C(_03374_),
    .Y(_03375_));
 sg13g2_nor3_1 _10990_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .Y(_03376_));
 sg13g2_nand3_1 _10991_ (.B(_03375_),
    .C(_03376_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .Y(_03377_));
 sg13g2_nor3_1 _10992_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .Y(_03378_));
 sg13g2_nand2_2 _10993_ (.Y(_03379_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .B(_03378_));
 sg13g2_or2_1 _10994_ (.X(_03380_),
    .B(_03379_),
    .A(_03377_));
 sg13g2_nor2_1 _10995_ (.A(_02549_),
    .B(_03380_),
    .Y(_03381_));
 sg13g2_nand2_1 _10996_ (.Y(_03382_),
    .A(\i_tinyqv.cpu.i_core.mip[0] ),
    .B(_03381_));
 sg13g2_nor2_1 _10997_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .Y(_03383_));
 sg13g2_nor3_1 _10998_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .Y(_03384_));
 sg13g2_nand2_2 _10999_ (.Y(_03385_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .B(_03384_));
 sg13g2_nand2_1 _11000_ (.Y(_03386_),
    .A(net2534),
    .B(_02539_));
 sg13g2_nor2_2 _11001_ (.A(net2369),
    .B(_03386_),
    .Y(_03387_));
 sg13g2_nand2_1 _11002_ (.Y(_03388_),
    .A(net4440),
    .B(net2533));
 sg13g2_nor3_1 _11003_ (.A(_03377_),
    .B(_03385_),
    .C(_03387_),
    .Y(_03389_));
 sg13g2_and2_1 _11004_ (.A(\i_tinyqv.cpu.i_core.mepc[0] ),
    .B(_03389_),
    .X(_03390_));
 sg13g2_nand2_1 _11005_ (.Y(_03391_),
    .A(_01997_),
    .B(_03376_));
 sg13g2_nor4_2 _11006_ (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .B(net2531),
    .C(_03374_),
    .Y(_03392_),
    .D(_03391_));
 sg13g2_nand2b_2 _11007_ (.Y(_03393_),
    .B(_03392_),
    .A_N(_03379_));
 sg13g2_nor2_1 _11008_ (.A(_02549_),
    .B(_03393_),
    .Y(_03394_));
 sg13g2_nor2b_1 _11009_ (.A(_03385_),
    .B_N(_03392_),
    .Y(_03395_));
 sg13g2_nand3b_1 _11010_ (.B(_03383_),
    .C(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .Y(_03396_),
    .A_N(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sg13g2_nor2_1 _11011_ (.A(_03377_),
    .B(_03396_),
    .Y(_03397_));
 sg13g2_nand2_1 _11012_ (.Y(_03398_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .B(net2531));
 sg13g2_or4_1 _11013_ (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .C(_03391_),
    .D(_03398_),
    .X(_03399_));
 sg13g2_nor2_2 _11014_ (.A(_03396_),
    .B(_03399_),
    .Y(_03400_));
 sg13g2_nor2b_2 _11015_ (.A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .B_N(_03384_),
    .Y(_03401_));
 sg13g2_nor2b_2 _11016_ (.A(_03399_),
    .B_N(_03401_),
    .Y(_03402_));
 sg13g2_nor2_2 _11017_ (.A(_03385_),
    .B(_03399_),
    .Y(_03403_));
 sg13g2_a221oi_1 _11018_ (.B2(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .C1(_03390_),
    .B1(_03400_),
    .A1(net2322),
    .Y(_03404_),
    .A2(_03395_));
 sg13g2_a22oi_1 _11019_ (.Y(_03405_),
    .B1(_03403_),
    .B2(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .A2(_03394_),
    .A1(\i_tinyqv.cpu.i_core.mie[0] ));
 sg13g2_a22oi_1 _11020_ (.Y(_03406_),
    .B1(net2320),
    .B2(\i_tinyqv.cpu.i_core.mcause[0] ),
    .A2(net2322),
    .A1(\i_tinyqv.cpu.i_core.mcause[4] ));
 sg13g2_inv_1 _11021_ (.Y(_03407_),
    .A(_03406_));
 sg13g2_a22oi_1 _11022_ (.Y(_03408_),
    .B1(_03407_),
    .B2(_03397_),
    .A2(_03402_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[0] ));
 sg13g2_nand4_1 _11023_ (.B(_03404_),
    .C(_03405_),
    .A(_03382_),
    .Y(_03409_),
    .D(_03408_));
 sg13g2_a22oi_1 _11024_ (.Y(_03410_),
    .B1(_03373_),
    .B2(_03409_),
    .A2(_03372_),
    .A1(_02803_));
 sg13g2_nand2_1 _11025_ (.Y(_03411_),
    .A(_02804_),
    .B(_03410_));
 sg13g2_o21ai_1 _11026_ (.B1(_03411_),
    .Y(_03412_),
    .A1(_02719_),
    .A2(_02804_));
 sg13g2_nor2b_1 _11027_ (.A(net2534),
    .B_N(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .Y(_03413_));
 sg13g2_nor3_1 _11028_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(_02707_),
    .C(_03413_),
    .Y(_03414_));
 sg13g2_or3_1 _11029_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(_02707_),
    .C(_03413_),
    .X(_03415_));
 sg13g2_a21oi_2 _11030_ (.B1(_03138_),
    .Y(_03416_),
    .A2(_03414_),
    .A1(\i_tinyqv.cpu.i_core.load_top_bit ));
 sg13g2_nand2_2 _11031_ (.Y(_03417_),
    .A(_02758_),
    .B(_03132_));
 sg13g2_mux2_1 _11032_ (.A0(net2596),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(net1908),
    .X(_03418_));
 sg13g2_o21ai_1 _11033_ (.B1(net2377),
    .Y(_03419_),
    .A1(\i_tinyqv.cpu.instr_data_in[8] ),
    .A2(net1908));
 sg13g2_a21oi_2 _11034_ (.B1(_03419_),
    .Y(_03420_),
    .A2(net1908),
    .A1(_02035_));
 sg13g2_nand4_1 _11035_ (.B(\i_tinyqv.cpu.data_write_n[0] ),
    .C(_02757_),
    .A(\i_tinyqv.cpu.data_read_n[0] ),
    .Y(_03421_),
    .D(_03132_));
 sg13g2_nand2b_1 _11036_ (.Y(_03422_),
    .B(net2410),
    .A_N(net1906));
 sg13g2_a21oi_1 _11037_ (.A1(_02063_),
    .A2(net1906),
    .Y(_03423_),
    .B1(net2379));
 sg13g2_a221oi_1 _11038_ (.B2(_03423_),
    .C1(_03420_),
    .B1(_03422_),
    .A1(net2369),
    .Y(_03424_),
    .A2(_03418_));
 sg13g2_a21oi_1 _11039_ (.A1(_02064_),
    .A2(net1907),
    .Y(_03425_),
    .B1(net2371));
 sg13g2_o21ai_1 _11040_ (.B1(_03425_),
    .Y(_03426_),
    .A1(net2596),
    .A2(net1907));
 sg13g2_nand3_1 _11041_ (.B(_03424_),
    .C(_03426_),
    .A(net2390),
    .Y(_03427_));
 sg13g2_o21ai_1 _11042_ (.B1(net2378),
    .Y(_03428_),
    .A1(_01807_),
    .A2(\i_latch_mem.data_out[0] ));
 sg13g2_nor2b_2 _11043_ (.A(\addr[5] ),
    .B_N(_02485_),
    .Y(_03429_));
 sg13g2_nand3_1 _11044_ (.B(\addr[5] ),
    .C(_02485_),
    .A(\addr[4] ),
    .Y(_03430_));
 sg13g2_nand2_2 _11045_ (.Y(_03431_),
    .A(_02013_),
    .B(_02474_));
 sg13g2_nor2_2 _11046_ (.A(_03430_),
    .B(_03431_),
    .Y(_03432_));
 sg13g2_nor2_2 _11047_ (.A(_02475_),
    .B(_03430_),
    .Y(_03433_));
 sg13g2_and2_1 _11048_ (.A(_02015_),
    .B(_02485_),
    .X(_03434_));
 sg13g2_nand2_1 _11049_ (.Y(_03435_),
    .A(_02015_),
    .B(_02485_));
 sg13g2_nand2_2 _11050_ (.Y(_03436_),
    .A(_02014_),
    .B(_03429_));
 sg13g2_nor2_2 _11051_ (.A(_03431_),
    .B(_03436_),
    .Y(_03437_));
 sg13g2_a21o_2 _11052_ (.A2(_03437_),
    .A1(uo_out[0]),
    .B1(net2174),
    .X(_03438_));
 sg13g2_a221oi_1 _11053_ (.B2(\i_wdt.counter[0] ),
    .C1(_03438_),
    .B1(net2116),
    .A1(\timer_count[0] ),
    .Y(_03439_),
    .A2(net2122));
 sg13g2_nand3_1 _11054_ (.B(net2466),
    .C(_03434_),
    .A(_02013_),
    .Y(_03440_));
 sg13g2_nor2_2 _11055_ (.A(_02487_),
    .B(_03440_),
    .Y(_03441_));
 sg13g2_nand2_2 _11056_ (.Y(_03442_),
    .A(\addr[4] ),
    .B(_03429_));
 sg13g2_nor2_1 _11057_ (.A(_03440_),
    .B(_03442_),
    .Y(_03443_));
 sg13g2_inv_1 _11058_ (.Y(_03444_),
    .A(net2083));
 sg13g2_a22oi_1 _11059_ (.Y(_03445_),
    .B1(net2083),
    .B2(\i2c_data_out[0] ),
    .A2(net2085),
    .A1(\i_rtc.seconds_out[0] ));
 sg13g2_nor2_1 _11060_ (.A(_02487_),
    .B(_03431_),
    .Y(_03446_));
 sg13g2_nor3_1 _11061_ (.A(net4715),
    .B(net4762),
    .C(net4021),
    .Y(_03447_));
 sg13g2_or3_1 _11062_ (.A(net4715),
    .B(net4762),
    .C(net4021),
    .X(_03448_));
 sg13g2_nand2_2 _11063_ (.Y(_03449_),
    .A(_01754_),
    .B(_03447_));
 sg13g2_nor2_2 _11064_ (.A(_02475_),
    .B(_03442_),
    .Y(_03450_));
 sg13g2_a22oi_1 _11065_ (.Y(_03451_),
    .B1(_03449_),
    .B2(_03450_),
    .A2(net2082),
    .A1(\i_spi.data[0] ));
 sg13g2_nand2b_2 _11066_ (.Y(_03452_),
    .B(_03434_),
    .A_N(_02095_));
 sg13g2_nor2_2 _11067_ (.A(_03436_),
    .B(_03452_),
    .Y(_03453_));
 sg13g2_a22oi_1 _11068_ (.Y(_03454_),
    .B1(_03453_),
    .B2(\gpio_out_sel[0] ),
    .A2(_02488_),
    .A1(net2457));
 sg13g2_nor2_2 _11069_ (.A(_03436_),
    .B(_03440_),
    .Y(_03455_));
 sg13g2_nor2_2 _11070_ (.A(_02095_),
    .B(_02487_),
    .Y(_03456_));
 sg13g2_nor2b_2 _11071_ (.A(net2488),
    .B_N(\i_seal.read_seq[0] ),
    .Y(_03457_));
 sg13g2_inv_1 _11072_ (.Y(_03458_),
    .A(net2351));
 sg13g2_nor2_1 _11073_ (.A(net2488),
    .B(\i_seal.read_seq[0] ),
    .Y(_03459_));
 sg13g2_a22oi_1 _11074_ (.Y(_03460_),
    .B1(net2345),
    .B2(\i_seal.sealed_value[0] ),
    .A2(net2351),
    .A1(\i_seal.sealed_mono[0] ));
 sg13g2_inv_1 _11075_ (.Y(_03461_),
    .A(_03460_));
 sg13g2_a22oi_1 _11076_ (.Y(_03462_),
    .B1(_03456_),
    .B2(_03461_),
    .A2(net2080),
    .A1(\crc16_read[0] ));
 sg13g2_nor2_2 _11077_ (.A(\i_seal.state[1] ),
    .B(\i_seal.state[0] ),
    .Y(_03463_));
 sg13g2_or2_1 _11078_ (.X(_03464_),
    .B(\i_seal.state[0] ),
    .A(\i_seal.state[1] ));
 sg13g2_nor3_2 _11079_ (.A(_02486_),
    .B(_03429_),
    .C(_03440_),
    .Y(_03465_));
 sg13g2_nor2_1 _11080_ (.A(_03442_),
    .B(_03452_),
    .Y(_03466_));
 sg13g2_a22oi_1 _11081_ (.Y(_03467_),
    .B1(net2078),
    .B2(\i2c_config_out[0] ),
    .A2(_03465_),
    .A1(net2341));
 sg13g2_nor2_2 _11082_ (.A(_03431_),
    .B(_03442_),
    .Y(_03468_));
 sg13g2_inv_2 _11083_ (.Y(_03469_),
    .A(net2076));
 sg13g2_nor2_2 _11084_ (.A(_02475_),
    .B(_03436_),
    .Y(_03470_));
 sg13g2_a22oi_1 _11085_ (.Y(_03471_),
    .B1(_03470_),
    .B2(net2),
    .A2(_03468_),
    .A1(\i_uart_rx.recieved_data[0] ));
 sg13g2_and4_1 _11086_ (.A(_03454_),
    .B(_03462_),
    .C(_03467_),
    .D(_03471_),
    .X(_03472_));
 sg13g2_nand4_1 _11087_ (.B(_03445_),
    .C(_03451_),
    .A(_03439_),
    .Y(_03473_),
    .D(_03472_));
 sg13g2_nand2b_2 _11088_ (.Y(_03474_),
    .B(_02489_),
    .A_N(\addr[5] ));
 sg13g2_nand4_1 _11089_ (.B(net2466),
    .C(_02015_),
    .A(_02013_),
    .Y(_03475_),
    .D(_02489_));
 sg13g2_nand3_1 _11090_ (.B(\addr[5] ),
    .C(_02489_),
    .A(\addr[4] ),
    .Y(_03476_));
 sg13g2_a21oi_1 _11091_ (.A1(_02095_),
    .A2(_02485_),
    .Y(_03477_),
    .B1(\addr[6] ));
 sg13g2_nor2b_2 _11092_ (.A(_02487_),
    .B_N(_03477_),
    .Y(_03478_));
 sg13g2_nand2b_1 _11093_ (.Y(_03479_),
    .B(_02486_),
    .A_N(\addr[5] ));
 sg13g2_nor2_2 _11094_ (.A(_03440_),
    .B(_03479_),
    .Y(_03480_));
 sg13g2_nand2b_1 _11095_ (.Y(_03481_),
    .B(_03473_),
    .A_N(_03428_));
 sg13g2_nor3_1 _11096_ (.A(_02486_),
    .B(_03429_),
    .C(_03452_),
    .Y(_03482_));
 sg13g2_nor2_1 _11097_ (.A(net2174),
    .B(net2074),
    .Y(_03483_));
 sg13g2_a22oi_1 _11098_ (.Y(_03484_),
    .B1(net2080),
    .B2(\crc16_read[8] ),
    .A2(net2083),
    .A1(\i2c_data_out[8] ));
 sg13g2_a22oi_1 _11099_ (.Y(_03485_),
    .B1(net2116),
    .B2(\i_wdt.counter[8] ),
    .A2(net2121),
    .A1(\timer_count[8] ));
 sg13g2_nand2_1 _11100_ (.Y(_03486_),
    .A(net2488),
    .B(\i_seal.sealed_crc[0] ));
 sg13g2_a22oi_1 _11101_ (.Y(_03487_),
    .B1(net2346),
    .B2(\i_seal.sealed_value[8] ),
    .A2(net2350),
    .A1(\i_seal.sealed_mono[8] ));
 sg13g2_nand2_1 _11102_ (.Y(_03488_),
    .A(_02015_),
    .B(_03456_));
 sg13g2_a21oi_2 _11103_ (.B1(net2005),
    .Y(_03489_),
    .A2(_03487_),
    .A1(_03486_));
 sg13g2_a221oi_1 _11104_ (.B2(\i2c_config_out[8] ),
    .C1(_03489_),
    .B1(net2077),
    .A1(\i_rtc.seconds_out[8] ),
    .Y(_03490_),
    .A2(net2085));
 sg13g2_nand4_1 _11105_ (.B(_03484_),
    .C(_03485_),
    .A(_03483_),
    .Y(_03491_),
    .D(_03490_));
 sg13g2_o21ai_1 _11106_ (.B1(net2384),
    .Y(_03492_),
    .A1(_01807_),
    .A2(\i_latch_mem.data_out[8] ));
 sg13g2_nand2b_1 _11107_ (.Y(_03493_),
    .B(_03491_),
    .A_N(_03492_));
 sg13g2_a21oi_1 _11108_ (.A1(net2468),
    .A2(_02065_),
    .Y(_03494_),
    .B1(net2370));
 sg13g2_a22oi_1 _11109_ (.Y(_03495_),
    .B1(net2345),
    .B2(\i_seal.sealed_value[12] ),
    .A2(\i_seal.sealed_crc[4] ),
    .A1(net2488));
 sg13g2_o21ai_1 _11110_ (.B1(_03495_),
    .Y(_03496_),
    .A1(_01935_),
    .A2(net2310));
 sg13g2_a22oi_1 _11111_ (.Y(_03497_),
    .B1(net2118),
    .B2(\i_wdt.counter[12] ),
    .A2(net2123),
    .A1(\timer_count[12] ));
 sg13g2_a22oi_1 _11112_ (.Y(_03498_),
    .B1(net2075),
    .B2(_03496_),
    .A2(net2085),
    .A1(\i_rtc.seconds_out[12] ));
 sg13g2_a22oi_1 _11113_ (.Y(_03499_),
    .B1(_03480_),
    .B2(\crc16_read[12] ),
    .A2(net2077),
    .A1(\i2c_config_out[12] ));
 sg13g2_nand4_1 _11114_ (.B(_03497_),
    .C(_03498_),
    .A(_03434_),
    .Y(_03500_),
    .D(_03499_));
 sg13g2_a21oi_1 _11115_ (.A1(net2467),
    .A2(_02062_),
    .Y(_03501_),
    .B1(net2366));
 sg13g2_nand2_1 _11116_ (.Y(_03502_),
    .A(\timer_count[4] ),
    .B(net2121));
 sg13g2_nand2_1 _11117_ (.Y(_03503_),
    .A(net6),
    .B(_03470_));
 sg13g2_nand3_1 _11118_ (.B(_03502_),
    .C(_03503_),
    .A(_03483_),
    .Y(_03504_));
 sg13g2_nand2_1 _11119_ (.Y(_03505_),
    .A(\i_wdt.counter[4] ),
    .B(net2117));
 sg13g2_a22oi_1 _11120_ (.Y(_03506_),
    .B1(net2347),
    .B2(\i_seal.sealed_value[4] ),
    .A2(net2350),
    .A1(\i_seal.sealed_mono[4] ));
 sg13g2_o21ai_1 _11121_ (.B1(_03505_),
    .Y(_03507_),
    .A1(net2002),
    .A2(_03506_));
 sg13g2_a22oi_1 _11122_ (.Y(_03508_),
    .B1(net2080),
    .B2(\crc16_read[4] ),
    .A2(net2082),
    .A1(\i_spi.data[4] ));
 sg13g2_a22oi_1 _11123_ (.Y(_03509_),
    .B1(net2076),
    .B2(\i_uart_rx.recieved_data[4] ),
    .A2(net2086),
    .A1(\i_rtc.seconds_out[4] ));
 sg13g2_a22oi_1 _11124_ (.Y(_03510_),
    .B1(_03453_),
    .B2(\gpio_out_sel[4] ),
    .A2(_03437_),
    .A1(uo_out[4]));
 sg13g2_a22oi_1 _11125_ (.Y(_03511_),
    .B1(net2079),
    .B2(\i2c_config_out[4] ),
    .A2(net2083),
    .A1(\i2c_data_out[4] ));
 sg13g2_nand4_1 _11126_ (.B(_03509_),
    .C(_03510_),
    .A(_03508_),
    .Y(_03512_),
    .D(_03511_));
 sg13g2_or3_1 _11127_ (.A(_03504_),
    .B(_03507_),
    .C(_03512_),
    .X(_03513_));
 sg13g2_a22oi_1 _11128_ (.Y(_03514_),
    .B1(_03501_),
    .B2(_03513_),
    .A2(_03500_),
    .A1(_03494_));
 sg13g2_nand4_1 _11129_ (.B(_03481_),
    .C(_03493_),
    .A(net2388),
    .Y(_03515_),
    .D(_03514_));
 sg13g2_and2_1 _11130_ (.A(net2435),
    .B(_03515_),
    .X(_03516_));
 sg13g2_a221oi_1 _11131_ (.B2(\pps_count[12] ),
    .C1(net2176),
    .B1(net2073),
    .A1(\i_rtc.seconds_out[28] ),
    .Y(_03517_),
    .A2(net2089));
 sg13g2_nand2_1 _11132_ (.Y(_03518_),
    .A(\i_seal.sealed_value[28] ),
    .B(net2342));
 sg13g2_a22oi_1 _11133_ (.Y(_03519_),
    .B1(net2348),
    .B2(\i_seal.sealed_sid[4] ),
    .A2(\i_seal.sealed_mono[28] ),
    .A1(net2491));
 sg13g2_a21oi_2 _11134_ (.B1(net2003),
    .Y(_03520_),
    .A2(_03519_),
    .A1(_03518_));
 sg13g2_a221oi_1 _11135_ (.B2(\i_wdt.counter[28] ),
    .C1(_03520_),
    .B1(net2120),
    .A1(\timer_count[28] ),
    .Y(_03521_),
    .A2(net2125));
 sg13g2_a221oi_1 _11136_ (.B2(_03521_),
    .C1(net2370),
    .B1(_03517_),
    .A1(net2470),
    .Y(_03522_),
    .A2(_02067_));
 sg13g2_o21ai_1 _11137_ (.B1(net2384),
    .Y(_03523_),
    .A1(_01807_),
    .A2(\i_latch_mem.data_out[24] ));
 sg13g2_a221oi_1 _11138_ (.B2(\pps_count[8] ),
    .C1(net2176),
    .B1(net2072),
    .A1(\i_rtc.seconds_out[24] ),
    .Y(_03524_),
    .A2(net2088));
 sg13g2_nand2_1 _11139_ (.Y(_03525_),
    .A(\i_seal.sealed_value[24] ),
    .B(net2342));
 sg13g2_a22oi_1 _11140_ (.Y(_03526_),
    .B1(net2348),
    .B2(\i_seal.sealed_sid[0] ),
    .A2(\i_seal.sealed_mono[24] ),
    .A1(net2491));
 sg13g2_a21oi_1 _11141_ (.A1(_03525_),
    .A2(_03526_),
    .Y(_03527_),
    .B1(net2003));
 sg13g2_a221oi_1 _11142_ (.B2(\i_wdt.counter[24] ),
    .C1(_03527_),
    .B1(net2119),
    .A1(\timer_count[24] ),
    .Y(_03528_),
    .A2(net2124));
 sg13g2_a21oi_1 _11143_ (.A1(_03524_),
    .A2(_03528_),
    .Y(_03529_),
    .B1(_03523_));
 sg13g2_nor3_2 _11144_ (.A(net2389),
    .B(_03522_),
    .C(_03529_),
    .Y(_03530_));
 sg13g2_mux2_1 _11145_ (.A0(net2597),
    .A1(\i_tinyqv.mem.qspi_data_buf[28] ),
    .S(_03133_),
    .X(_03531_));
 sg13g2_nor2_1 _11146_ (.A(\i_tinyqv.mem.qspi_data_buf[24] ),
    .B(_03132_),
    .Y(_03532_));
 sg13g2_a21oi_1 _11147_ (.A1(net2410),
    .A2(_03132_),
    .Y(_03533_),
    .B1(_03532_));
 sg13g2_a221oi_1 _11148_ (.B2(net2382),
    .C1(net2387),
    .B1(_03533_),
    .A1(net2374),
    .Y(_03534_),
    .A2(_03531_));
 sg13g2_nor3_1 _11149_ (.A(net2435),
    .B(_03530_),
    .C(_03534_),
    .Y(_03535_));
 sg13g2_nor3_2 _11150_ (.A(\i_crc16.bit_cnt[2] ),
    .B(net4280),
    .C(net3481),
    .Y(_03536_));
 sg13g2_nor2b_2 _11151_ (.A(net4170),
    .B_N(_03536_),
    .Y(_03537_));
 sg13g2_nand2b_2 _11152_ (.Y(_03538_),
    .B(_03536_),
    .A_N(net4170));
 sg13g2_nand2_1 _11153_ (.Y(_03539_),
    .A(_03463_),
    .B(net2308));
 sg13g2_a22oi_1 _11154_ (.Y(_03540_),
    .B1(net2345),
    .B2(\i_seal.sealed_value[16] ),
    .A2(\i_seal.sealed_crc[8] ),
    .A1(net2489));
 sg13g2_o21ai_1 _11155_ (.B1(_03540_),
    .Y(_03541_),
    .A1(_01931_),
    .A2(net2310));
 sg13g2_a22oi_1 _11156_ (.Y(_03542_),
    .B1(net2072),
    .B2(\pps_count[4] ),
    .A2(net2088),
    .A1(\i_rtc.seconds_out[20] ));
 sg13g2_a22oi_1 _11157_ (.Y(_03543_),
    .B1(net2343),
    .B2(\i_seal.sealed_value[20] ),
    .A2(net2349),
    .A1(\i_seal.sealed_mono[20] ));
 sg13g2_o21ai_1 _11158_ (.B1(_03543_),
    .Y(_03544_),
    .A1(_01809_),
    .A2(_01942_));
 sg13g2_a22oi_1 _11159_ (.Y(_03545_),
    .B1(_03541_),
    .B2(net2075),
    .A2(_03539_),
    .A1(_03480_));
 sg13g2_a22oi_1 _11160_ (.Y(_03546_),
    .B1(net2073),
    .B2(\pps_count[0] ),
    .A2(net2089),
    .A1(\i_rtc.seconds_out[16] ));
 sg13g2_a22oi_1 _11161_ (.Y(_03547_),
    .B1(net2118),
    .B2(\i_wdt.counter[16] ),
    .A2(net2125),
    .A1(\timer_count[16] ));
 sg13g2_nand4_1 _11162_ (.B(_03545_),
    .C(_03546_),
    .A(net2438),
    .Y(_03548_),
    .D(_03547_));
 sg13g2_nand2_1 _11163_ (.Y(_03549_),
    .A(net2075),
    .B(_03544_));
 sg13g2_a22oi_1 _11164_ (.Y(_03550_),
    .B1(net2119),
    .B2(\i_wdt.counter[20] ),
    .A2(net2124),
    .A1(\timer_count[20] ));
 sg13g2_nand4_1 _11165_ (.B(_03542_),
    .C(_03549_),
    .A(net2542),
    .Y(_03551_),
    .D(_03550_));
 sg13g2_a21oi_1 _11166_ (.A1(_03548_),
    .A2(_03551_),
    .Y(_03552_),
    .B1(net2177));
 sg13g2_o21ai_1 _11167_ (.B1(net2470),
    .Y(_03553_),
    .A1(net2541),
    .A2(\i_latch_mem.data_out[16] ));
 sg13g2_a21oi_1 _11168_ (.A1(net2541),
    .A2(_02066_),
    .Y(_03554_),
    .B1(_03553_));
 sg13g2_nor2_1 _11169_ (.A(net2389),
    .B(_03554_),
    .Y(_03555_));
 sg13g2_o21ai_1 _11170_ (.B1(_03555_),
    .Y(_03556_),
    .A1(net2471),
    .A2(_03552_));
 sg13g2_nand2_1 _11171_ (.Y(_03557_),
    .A(net2540),
    .B(\i_tinyqv.mem.data_from_read[20] ));
 sg13g2_a21oi_1 _11172_ (.A1(net2438),
    .A2(\i_tinyqv.mem.data_from_read[16] ),
    .Y(_03558_),
    .B1(net2387));
 sg13g2_a21oi_1 _11173_ (.A1(_03557_),
    .A2(_03558_),
    .Y(_03559_),
    .B1(_02547_));
 sg13g2_a221oi_1 _11174_ (.B2(_03559_),
    .C1(_03535_),
    .B1(_03556_),
    .A1(_03427_),
    .Y(_03560_),
    .A2(_03516_));
 sg13g2_or2_1 _11175_ (.X(_03561_),
    .B(_03560_),
    .A(_03414_));
 sg13g2_a221oi_1 _11176_ (.B2(_03561_),
    .C1(_03143_),
    .B1(_03416_),
    .A1(_03138_),
    .Y(_03562_),
    .A2(_03412_));
 sg13g2_inv_1 _11177_ (.Y(_03563_),
    .A(_03562_));
 sg13g2_o21ai_1 _11178_ (.B1(_03563_),
    .Y(_03564_),
    .A1(_03142_),
    .A2(_03344_));
 sg13g2_mux2_1 _11179_ (.A0(net1816),
    .A1(net4802),
    .S(_03150_),
    .X(_00066_));
 sg13g2_xor2_1 _11180_ (.B(_02744_),
    .A(_02743_),
    .X(_03565_));
 sg13g2_and2_1 _11181_ (.A(_02776_),
    .B(_03156_),
    .X(_03566_));
 sg13g2_o21ai_1 _11182_ (.B1(_02001_),
    .Y(_03567_),
    .A1(_02674_),
    .A2(_02690_));
 sg13g2_nand2_1 _11183_ (.Y(_03568_),
    .A(_02775_),
    .B(_03567_));
 sg13g2_a221oi_1 _11184_ (.B2(_03157_),
    .C1(_03566_),
    .B1(_03568_),
    .A1(_03153_),
    .Y(_03569_),
    .A2(_03565_));
 sg13g2_nand2_1 _11185_ (.Y(_03570_),
    .A(_03145_),
    .B(_03569_));
 sg13g2_xor2_1 _11186_ (.B(_02868_),
    .A(_02867_),
    .X(_03571_));
 sg13g2_o21ai_1 _11187_ (.B1(_03570_),
    .Y(_03572_),
    .A1(_03145_),
    .A2(_03571_));
 sg13g2_nor2_1 _11188_ (.A(net2474),
    .B(_03327_),
    .Y(_03573_));
 sg13g2_o21ai_1 _11189_ (.B1(net2311),
    .Y(_03574_),
    .A1(net2407),
    .A2(_03323_));
 sg13g2_mux2_1 _11190_ (.A0(_03314_),
    .A1(_03325_),
    .S(net2407),
    .X(_03575_));
 sg13g2_a21oi_1 _11191_ (.A1(net2313),
    .A2(_03575_),
    .Y(_03576_),
    .B1(net2178));
 sg13g2_o21ai_1 _11192_ (.B1(_03576_),
    .Y(_03577_),
    .A1(_03573_),
    .A2(_03574_));
 sg13g2_nor2_1 _11193_ (.A(net2408),
    .B(_03293_),
    .Y(_03578_));
 sg13g2_o21ai_1 _11194_ (.B1(net2312),
    .Y(_03579_),
    .A1(net2475),
    .A2(_03283_));
 sg13g2_nor2_1 _11195_ (.A(net2407),
    .B(_03303_),
    .Y(_03580_));
 sg13g2_a21oi_1 _11196_ (.A1(net2408),
    .A2(_03296_),
    .Y(_03581_),
    .B1(_03580_));
 sg13g2_a21oi_1 _11197_ (.A1(net2314),
    .A2(_03581_),
    .Y(_03582_),
    .B1(_03195_));
 sg13g2_o21ai_1 _11198_ (.B1(_03582_),
    .Y(_03583_),
    .A1(_03578_),
    .A2(_03579_));
 sg13g2_nand3_1 _11199_ (.B(_03577_),
    .C(_03583_),
    .A(_03232_),
    .Y(_03584_));
 sg13g2_mux2_1 _11200_ (.A0(_03313_),
    .A1(_03320_),
    .S(net2475),
    .X(_03585_));
 sg13g2_nand2b_1 _11201_ (.Y(_03586_),
    .B(net2409),
    .A_N(_03318_));
 sg13g2_a22oi_1 _11202_ (.Y(_03587_),
    .B1(_03586_),
    .B2(_03250_),
    .A2(_03585_),
    .A1(_03187_));
 sg13g2_a21oi_1 _11203_ (.A1(net2406),
    .A2(_03307_),
    .Y(_03588_),
    .B1(net2311));
 sg13g2_o21ai_1 _11204_ (.B1(_03588_),
    .Y(_03589_),
    .A1(net2406),
    .A2(_03329_));
 sg13g2_nor2_1 _11205_ (.A(net2406),
    .B(_03309_),
    .Y(_03590_));
 sg13g2_a21oi_1 _11206_ (.A1(net2407),
    .A2(_03301_),
    .Y(_03591_),
    .B1(_03590_));
 sg13g2_a21oi_1 _11207_ (.A1(net2312),
    .A2(_03591_),
    .Y(_03592_),
    .B1(_03195_));
 sg13g2_a221oi_1 _11208_ (.B2(_03592_),
    .C1(_03232_),
    .B1(_03589_),
    .A1(_03195_),
    .Y(_03593_),
    .A2(_03587_));
 sg13g2_nor2_1 _11209_ (.A(_03178_),
    .B(_03593_),
    .Y(_03594_));
 sg13g2_a21oi_1 _11210_ (.A1(_03584_),
    .A2(_03594_),
    .Y(_03595_),
    .B1(_03179_));
 sg13g2_mux4_1 _11211_ (.S0(net2477),
    .A0(_03189_),
    .A1(_03191_),
    .A2(_03254_),
    .A3(_03256_),
    .S1(net2407),
    .X(_03596_));
 sg13g2_mux4_1 _11212_ (.S0(net2477),
    .A0(_03182_),
    .A1(_03184_),
    .A2(_03198_),
    .A3(_03199_),
    .S1(net2474),
    .X(_03597_));
 sg13g2_mux2_1 _11213_ (.A0(_03244_),
    .A1(_03249_),
    .S(net2476),
    .X(_03598_));
 sg13g2_or2_1 _11214_ (.X(_03599_),
    .B(_03238_),
    .A(net2409));
 sg13g2_a21oi_1 _11215_ (.A1(_03202_),
    .A2(_03203_),
    .Y(_03600_),
    .B1(net2473));
 sg13g2_nor2_1 _11216_ (.A(net2314),
    .B(_03600_),
    .Y(_03601_));
 sg13g2_nand2b_1 _11217_ (.Y(_03602_),
    .B(_03286_),
    .A_N(net2485));
 sg13g2_a21oi_1 _11218_ (.A1(net2483),
    .A2(_03282_),
    .Y(_03603_),
    .B1(net2475));
 sg13g2_a21o_1 _11219_ (.A2(_03262_),
    .A1(net2474),
    .B1(net2311),
    .X(_03604_));
 sg13g2_a21o_1 _11220_ (.A2(_03269_),
    .A1(net2406),
    .B1(_03604_),
    .X(_03605_));
 sg13g2_and2_1 _11221_ (.A(net2406),
    .B(_03216_),
    .X(_03606_));
 sg13g2_o21ai_1 _11222_ (.B1(net2311),
    .Y(_03607_),
    .A1(net2406),
    .A2(_03274_));
 sg13g2_a21oi_1 _11223_ (.A1(net2313),
    .A2(_03597_),
    .Y(_03608_),
    .B1(net2178));
 sg13g2_o21ai_1 _11224_ (.B1(_03608_),
    .Y(_03609_),
    .A1(net2313),
    .A2(_03596_));
 sg13g2_a221oi_1 _11225_ (.B2(_03603_),
    .C1(net2313),
    .B1(_03602_),
    .A1(net2475),
    .Y(_03610_),
    .A2(_03228_));
 sg13g2_nor2_1 _11226_ (.A(net2408),
    .B(_03211_),
    .Y(_03611_));
 sg13g2_a21o_1 _11227_ (.A2(_03223_),
    .A1(net2408),
    .B1(_03187_),
    .X(_03612_));
 sg13g2_nor2_1 _11228_ (.A(_03611_),
    .B(_03612_),
    .Y(_03613_));
 sg13g2_or3_1 _11229_ (.A(_03195_),
    .B(_03610_),
    .C(_03613_),
    .X(_03614_));
 sg13g2_nand3_1 _11230_ (.B(_03609_),
    .C(_03614_),
    .A(_03232_),
    .Y(_03615_));
 sg13g2_and2_1 _11231_ (.A(net2178),
    .B(_03605_),
    .X(_03616_));
 sg13g2_o21ai_1 _11232_ (.B1(_03616_),
    .Y(_03617_),
    .A1(_03606_),
    .A2(_03607_));
 sg13g2_a221oi_1 _11233_ (.B2(_03601_),
    .C1(_03194_),
    .B1(_03599_),
    .A1(net2314),
    .Y(_03618_),
    .A2(_03598_));
 sg13g2_nor2_1 _11234_ (.A(_03232_),
    .B(_03618_),
    .Y(_03619_));
 sg13g2_a21oi_1 _11235_ (.A1(_03617_),
    .A2(_03619_),
    .Y(_03620_),
    .B1(_03178_));
 sg13g2_a21oi_1 _11236_ (.A1(_03615_),
    .A2(_03620_),
    .Y(_03621_),
    .B1(_03179_));
 sg13g2_nor2_1 _11237_ (.A(net2524),
    .B(_03595_),
    .Y(_03622_));
 sg13g2_o21ai_1 _11238_ (.B1(_03166_),
    .Y(_03623_),
    .A1(net2434),
    .A2(_03621_));
 sg13g2_o21ai_1 _11239_ (.B1(_03572_),
    .Y(_03624_),
    .A1(_03622_),
    .A2(_03623_));
 sg13g2_a22oi_1 _11240_ (.Y(_03625_),
    .B1(_03342_),
    .B2(_03624_),
    .A2(_03152_),
    .A1(net2588));
 sg13g2_or2_1 _11241_ (.X(_03626_),
    .B(_03360_),
    .A(_01969_));
 sg13g2_xnor2_1 _11242_ (.Y(_03627_),
    .A(_01969_),
    .B(_03360_));
 sg13g2_xnor2_1 _11243_ (.Y(_03628_),
    .A(net2569),
    .B(_03355_));
 sg13g2_xor2_1 _11244_ (.B(_03349_),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(_03629_));
 sg13g2_xnor2_1 _11245_ (.Y(_03630_),
    .A(\i_tinyqv.cpu.instr_len[1] ),
    .B(\i_tinyqv.cpu.pc[1] ));
 sg13g2_a221oi_1 _11246_ (.B2(net2378),
    .C1(net2532),
    .B1(_03630_),
    .A1(net2368),
    .Y(_03631_),
    .A2(_03629_));
 sg13g2_xnor2_1 _11247_ (.Y(_03632_),
    .A(_01975_),
    .B(_03352_));
 sg13g2_a22oi_1 _11248_ (.Y(_03633_),
    .B1(_03632_),
    .B2(net2382),
    .A2(_03628_),
    .A1(net2373));
 sg13g2_a21o_1 _11249_ (.A2(_03357_),
    .A1(\i_tinyqv.cpu.instr_data_start[16] ),
    .B1(net2566),
    .X(_03634_));
 sg13g2_nand2_1 _11250_ (.Y(_03635_),
    .A(_03358_),
    .B(_03634_));
 sg13g2_inv_1 _11251_ (.Y(_03636_),
    .A(_03635_));
 sg13g2_a22oi_1 _11252_ (.Y(_03637_),
    .B1(_03636_),
    .B2(net2323),
    .A2(_03633_),
    .A1(_03631_));
 sg13g2_o21ai_1 _11253_ (.B1(_03637_),
    .Y(_03638_),
    .A1(_02551_),
    .A2(_03627_));
 sg13g2_and2_1 _11254_ (.A(\i_tinyqv.cpu.i_core.mepc[1] ),
    .B(_03389_),
    .X(_03639_));
 sg13g2_a22oi_1 _11255_ (.Y(_03640_),
    .B1(_03394_),
    .B2(\i_tinyqv.cpu.i_core.mie[1] ),
    .A2(_03381_),
    .A1(\i_tinyqv.cpu.i_core.mip[1] ));
 sg13g2_and4_1 _11256_ (.A(_01997_),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .D(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .X(_03641_));
 sg13g2_nand3_1 _11257_ (.B(net2531),
    .C(_03383_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .Y(_03642_));
 sg13g2_nor4_1 _11258_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .C(_03374_),
    .D(_03642_),
    .Y(_03643_));
 sg13g2_a22oi_1 _11259_ (.Y(_03644_),
    .B1(_03641_),
    .B2(_03643_),
    .A2(_03397_),
    .A1(\i_tinyqv.cpu.i_core.mcause[1] ));
 sg13g2_nand2b_1 _11260_ (.Y(_03645_),
    .B(net2321),
    .A_N(_03644_));
 sg13g2_mux2_1 _11261_ (.A0(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .S(net2316),
    .X(_03646_));
 sg13g2_nand2_1 _11262_ (.Y(_03647_),
    .A(_03403_),
    .B(_03646_));
 sg13g2_a221oi_1 _11263_ (.B2(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .C1(_03639_),
    .B1(_03402_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .Y(_03648_),
    .A2(_03400_));
 sg13g2_nand4_1 _11264_ (.B(_03645_),
    .C(_03647_),
    .A(_03640_),
    .Y(_03649_),
    .D(_03648_));
 sg13g2_a22oi_1 _11265_ (.Y(_03650_),
    .B1(_03649_),
    .B2(_03373_),
    .A2(_03638_),
    .A1(_02803_));
 sg13g2_nand2_1 _11266_ (.Y(_03651_),
    .A(_02804_),
    .B(_03650_));
 sg13g2_o21ai_1 _11267_ (.B1(_03651_),
    .Y(_03652_),
    .A1(_02689_),
    .A2(_02804_));
 sg13g2_nand2_1 _11268_ (.Y(_03653_),
    .A(_03138_),
    .B(_03652_));
 sg13g2_nand2_1 _11269_ (.Y(_03654_),
    .A(\i_rtc.seconds_out[9] ),
    .B(net2085));
 sg13g2_a22oi_1 _11270_ (.Y(_03655_),
    .B1(net2346),
    .B2(\i_seal.sealed_value[9] ),
    .A2(\i_seal.sealed_crc[1] ),
    .A1(net2488));
 sg13g2_o21ai_1 _11271_ (.B1(_03655_),
    .Y(_03656_),
    .A1(_01938_),
    .A2(net2310));
 sg13g2_a22oi_1 _11272_ (.Y(_03657_),
    .B1(net2075),
    .B2(_03656_),
    .A2(net2084),
    .A1(\i_i2c_peri.i_i2c.busy_reg ));
 sg13g2_a22oi_1 _11273_ (.Y(_03658_),
    .B1(_03480_),
    .B2(\crc16_read[9] ),
    .A2(net2077),
    .A1(\i2c_config_out[9] ));
 sg13g2_a221oi_1 _11274_ (.B2(\i_wdt.counter[9] ),
    .C1(net2174),
    .B1(net2116),
    .A1(\timer_count[9] ),
    .Y(_03659_),
    .A2(net2121));
 sg13g2_nand4_1 _11275_ (.B(_03657_),
    .C(_03658_),
    .A(_03654_),
    .Y(_03660_),
    .D(_03659_));
 sg13g2_o21ai_1 _11276_ (.B1(_03660_),
    .Y(_03661_),
    .A1(_01807_),
    .A2(\i_latch_mem.data_out[9] ));
 sg13g2_nor3_1 _11277_ (.A(net2389),
    .B(net2380),
    .C(_03661_),
    .Y(_03662_));
 sg13g2_a21oi_1 _11278_ (.A1(net2472),
    .A2(_02069_),
    .Y(_03663_),
    .B1(_02539_));
 sg13g2_a22oi_1 _11279_ (.Y(_03664_),
    .B1(net2346),
    .B2(\i_seal.sealed_value[1] ),
    .A2(net2351),
    .A1(\i_seal.sealed_mono[1] ));
 sg13g2_nor2_1 _11280_ (.A(net2002),
    .B(_03664_),
    .Y(_03665_));
 sg13g2_a221oi_1 _11281_ (.B2(\i_wdt.counter[1] ),
    .C1(_03665_),
    .B1(net2117),
    .A1(\timer_count[1] ),
    .Y(_03666_),
    .A2(net2122));
 sg13g2_nor2b_1 _11282_ (.A(net4787),
    .B_N(\i_uart_rx.fsm_state[3] ),
    .Y(_03667_));
 sg13g2_nand2_1 _11283_ (.Y(_03668_),
    .A(net5236),
    .B(_01750_));
 sg13g2_and2_1 _11284_ (.A(net2459),
    .B(_03667_),
    .X(_03669_));
 sg13g2_nand2_1 _11285_ (.Y(_03670_),
    .A(net2459),
    .B(_03667_));
 sg13g2_and2_1 _11286_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_03669_),
    .X(_03671_));
 sg13g2_a22oi_1 _11287_ (.Y(_03672_),
    .B1(_03671_),
    .B2(_03450_),
    .A2(net2080),
    .A1(\crc16_read[1] ));
 sg13g2_a22oi_1 _11288_ (.Y(_03673_),
    .B1(net2086),
    .B2(\i_rtc.seconds_out[1] ),
    .A2(_03437_),
    .A1(uo_out[1]));
 sg13g2_a22oi_1 _11289_ (.Y(_03674_),
    .B1(net2076),
    .B2(\i_uart_rx.recieved_data[1] ),
    .A2(_03453_),
    .A1(\gpio_out_sel[1] ));
 sg13g2_a22oi_1 _11290_ (.Y(_03675_),
    .B1(net2078),
    .B2(\i2c_config_out[1] ),
    .A2(net2082),
    .A1(\i_spi.data[1] ));
 sg13g2_a21oi_1 _11291_ (.A1(_03463_),
    .A2(_03465_),
    .Y(_03676_),
    .B1(net2174));
 sg13g2_a22oi_1 _11292_ (.Y(_03677_),
    .B1(_03470_),
    .B2(net3),
    .A2(net2083),
    .A1(\i2c_data_out[1] ));
 sg13g2_and4_1 _11293_ (.A(_03674_),
    .B(_03675_),
    .C(_03676_),
    .D(_03677_),
    .X(_03678_));
 sg13g2_nand4_1 _11294_ (.B(_03672_),
    .C(_03673_),
    .A(_03666_),
    .Y(_03679_),
    .D(_03678_));
 sg13g2_nand2b_1 _11295_ (.Y(_03680_),
    .B(net2467),
    .A_N(\i_latch_mem.data_out[13] ));
 sg13g2_a22oi_1 _11296_ (.Y(_03681_),
    .B1(net2346),
    .B2(\i_seal.sealed_value[13] ),
    .A2(\i_seal.sealed_crc[5] ),
    .A1(net2489));
 sg13g2_o21ai_1 _11297_ (.B1(_03681_),
    .Y(_03682_),
    .A1(_01934_),
    .A2(net2310));
 sg13g2_a22oi_1 _11298_ (.Y(_03683_),
    .B1(net2118),
    .B2(\i_wdt.counter[13] ),
    .A2(net2123),
    .A1(\timer_count[13] ));
 sg13g2_a22oi_1 _11299_ (.Y(_03684_),
    .B1(_03682_),
    .B2(net2075),
    .A2(_03480_),
    .A1(\crc16_read[13] ));
 sg13g2_a22oi_1 _11300_ (.Y(_03685_),
    .B1(net2077),
    .B2(\i2c_config_out[13] ),
    .A2(net2086),
    .A1(\i_rtc.seconds_out[13] ));
 sg13g2_nand4_1 _11301_ (.B(_03683_),
    .C(_03684_),
    .A(_03434_),
    .Y(_03686_),
    .D(_03685_));
 sg13g2_nand3_1 _11302_ (.B(_03680_),
    .C(_03686_),
    .A(net2374),
    .Y(_03687_));
 sg13g2_a21oi_1 _11303_ (.A1(net2467),
    .A2(_02070_),
    .Y(_03688_),
    .B1(net2366));
 sg13g2_a22oi_1 _11304_ (.Y(_03689_),
    .B1(net2116),
    .B2(\i_wdt.counter[5] ),
    .A2(net2121),
    .A1(\timer_count[5] ));
 sg13g2_a21oi_1 _11305_ (.A1(\i_spi.data[5] ),
    .A2(net2082),
    .Y(_03690_),
    .B1(net2174));
 sg13g2_a22oi_1 _11306_ (.Y(_03691_),
    .B1(net2346),
    .B2(\i_seal.sealed_value[5] ),
    .A2(net2350),
    .A1(\i_seal.sealed_mono[5] ));
 sg13g2_inv_1 _11307_ (.Y(_03692_),
    .A(_03691_));
 sg13g2_a22oi_1 _11308_ (.Y(_03693_),
    .B1(_03456_),
    .B2(_03692_),
    .A2(net2085),
    .A1(\i_rtc.seconds_out[5] ));
 sg13g2_nand2_2 _11309_ (.Y(_03694_),
    .A(\crc16_read[5] ),
    .B(net2081));
 sg13g2_a22oi_1 _11310_ (.Y(_03695_),
    .B1(net2076),
    .B2(\i_uart_rx.recieved_data[5] ),
    .A2(_03453_),
    .A1(\gpio_out_sel[5] ));
 sg13g2_a22oi_1 _11311_ (.Y(_03696_),
    .B1(net2079),
    .B2(\i2c_config_out[5] ),
    .A2(net2083),
    .A1(\i2c_data_out[5] ));
 sg13g2_a22oi_1 _11312_ (.Y(_03697_),
    .B1(_03470_),
    .B2(net7),
    .A2(_03437_),
    .A1(uo_out[5]));
 sg13g2_and4_1 _11313_ (.A(_03694_),
    .B(_03695_),
    .C(_03696_),
    .D(_03697_),
    .X(_03698_));
 sg13g2_nand4_1 _11314_ (.B(_03690_),
    .C(_03693_),
    .A(_03689_),
    .Y(_03699_),
    .D(_03698_));
 sg13g2_nor2_1 _11315_ (.A(net2602),
    .B(net1908),
    .Y(_03700_));
 sg13g2_a21oi_1 _11316_ (.A1(_02036_),
    .A2(net1908),
    .Y(_03701_),
    .B1(_03700_));
 sg13g2_mux2_1 _11317_ (.A0(net2594),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(net1908),
    .X(_03702_));
 sg13g2_o21ai_1 _11318_ (.B1(net2383),
    .Y(_03703_),
    .A1(net2602),
    .A2(net1906));
 sg13g2_a21oi_2 _11319_ (.B1(_03703_),
    .Y(_03704_),
    .A2(net1906),
    .A1(_02071_));
 sg13g2_a21oi_1 _11320_ (.A1(_02072_),
    .A2(net1907),
    .Y(_03705_),
    .B1(net2371));
 sg13g2_o21ai_1 _11321_ (.B1(_03705_),
    .Y(_03706_),
    .A1(net2594),
    .A2(net1907));
 sg13g2_a22oi_1 _11322_ (.Y(_03707_),
    .B1(_03688_),
    .B2(_03699_),
    .A2(_03679_),
    .A1(_03663_));
 sg13g2_a21oi_1 _11323_ (.A1(_03687_),
    .A2(_03707_),
    .Y(_03708_),
    .B1(net2389));
 sg13g2_a221oi_1 _11324_ (.B2(net2368),
    .C1(_03704_),
    .B1(_03702_),
    .A1(net2377),
    .Y(_03709_),
    .A2(_03701_));
 sg13g2_a21oi_1 _11325_ (.A1(_03706_),
    .A2(_03709_),
    .Y(_03710_),
    .B1(net2387));
 sg13g2_nor4_1 _11326_ (.A(net2534),
    .B(_03662_),
    .C(_03708_),
    .D(_03710_),
    .Y(_03711_));
 sg13g2_a221oi_1 _11327_ (.B2(\pps_count[9] ),
    .C1(net2176),
    .B1(net2072),
    .A1(\i_rtc.seconds_out[25] ),
    .Y(_03712_),
    .A2(net2088));
 sg13g2_nand2_1 _11328_ (.Y(_03713_),
    .A(\i_seal.sealed_value[25] ),
    .B(net2342));
 sg13g2_a22oi_1 _11329_ (.Y(_03714_),
    .B1(net2348),
    .B2(\i_seal.sealed_sid[1] ),
    .A2(\i_seal.sealed_mono[25] ),
    .A1(net2491));
 sg13g2_a21oi_2 _11330_ (.B1(net2003),
    .Y(_03715_),
    .A2(_03714_),
    .A1(_03713_));
 sg13g2_a221oi_1 _11331_ (.B2(\i_wdt.counter[25] ),
    .C1(_03715_),
    .B1(net2120),
    .A1(\timer_count[25] ),
    .Y(_03716_),
    .A2(net2124));
 sg13g2_a221oi_1 _11332_ (.B2(_03716_),
    .C1(net2379),
    .B1(_03712_),
    .A1(net2470),
    .Y(_03717_),
    .A2(_02073_));
 sg13g2_a221oi_1 _11333_ (.B2(\pps_count[13] ),
    .C1(net2176),
    .B1(net2073),
    .A1(\i_rtc.seconds_out[29] ),
    .Y(_03718_),
    .A2(net2089));
 sg13g2_nand2_1 _11334_ (.Y(_03719_),
    .A(\i_seal.sealed_value[29] ),
    .B(net2342));
 sg13g2_a22oi_1 _11335_ (.Y(_03720_),
    .B1(net2348),
    .B2(\i_seal.sealed_sid[5] ),
    .A2(\i_seal.sealed_mono[29] ),
    .A1(net2491));
 sg13g2_a21oi_2 _11336_ (.B1(net2003),
    .Y(_03721_),
    .A2(_03720_),
    .A1(_03719_));
 sg13g2_a221oi_1 _11337_ (.B2(\i_wdt.counter[29] ),
    .C1(_03721_),
    .B1(net2120),
    .A1(\timer_count[29] ),
    .Y(_03722_),
    .A2(net2125));
 sg13g2_a221oi_1 _11338_ (.B2(_03722_),
    .C1(net2370),
    .B1(_03718_),
    .A1(net2470),
    .Y(_03723_),
    .A2(_02074_));
 sg13g2_nor3_1 _11339_ (.A(net2389),
    .B(_03717_),
    .C(_03723_),
    .Y(_03724_));
 sg13g2_mux2_1 _11340_ (.A0(net2603),
    .A1(\i_tinyqv.mem.qspi_data_buf[25] ),
    .S(_03133_),
    .X(_03725_));
 sg13g2_mux2_1 _11341_ (.A0(net2595),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .S(_03133_),
    .X(_03726_));
 sg13g2_a221oi_1 _11342_ (.B2(net2374),
    .C1(net2387),
    .B1(_03726_),
    .A1(net2382),
    .Y(_03727_),
    .A2(_03725_));
 sg13g2_and2_1 _11343_ (.A(net2541),
    .B(\i_latch_mem.data_out[21] ),
    .X(_03728_));
 sg13g2_a21oi_1 _11344_ (.A1(net2438),
    .A2(\i_latch_mem.data_out[17] ),
    .Y(_03729_),
    .B1(_03728_));
 sg13g2_and2_1 _11345_ (.A(net2540),
    .B(\i_tinyqv.mem.data_from_read[21] ),
    .X(_03730_));
 sg13g2_a21oi_1 _11346_ (.A1(net2438),
    .A2(\i_tinyqv.mem.data_from_read[17] ),
    .Y(_03731_),
    .B1(_03730_));
 sg13g2_a221oi_1 _11347_ (.B2(net2389),
    .C1(net2537),
    .B1(_03731_),
    .A1(net2469),
    .Y(_03732_),
    .A2(_03729_));
 sg13g2_a221oi_1 _11348_ (.B2(\pps_count[1] ),
    .C1(net2542),
    .B1(net2073),
    .A1(\i_rtc.seconds_out[17] ),
    .Y(_03733_),
    .A2(net2089));
 sg13g2_nand2_1 _11349_ (.Y(_03734_),
    .A(\i_seal.sealed_mono[17] ),
    .B(net2350));
 sg13g2_a22oi_1 _11350_ (.Y(_03735_),
    .B1(net2343),
    .B2(\i_seal.sealed_value[17] ),
    .A2(\i_seal.sealed_crc[9] ),
    .A1(net2491));
 sg13g2_a21oi_2 _11351_ (.B1(net2003),
    .Y(_03736_),
    .A2(_03735_),
    .A1(_03734_));
 sg13g2_a221oi_1 _11352_ (.B2(\i_wdt.counter[17] ),
    .C1(_03736_),
    .B1(net2120),
    .A1(\timer_count[17] ),
    .Y(_03737_),
    .A2(net2125));
 sg13g2_a221oi_1 _11353_ (.B2(\pps_count[5] ),
    .C1(net2438),
    .B1(net2072),
    .A1(\i_rtc.seconds_out[21] ),
    .Y(_03738_),
    .A2(net2088));
 sg13g2_nand2_1 _11354_ (.Y(_03739_),
    .A(\i_seal.sealed_value[21] ),
    .B(net2344));
 sg13g2_a22oi_1 _11355_ (.Y(_03740_),
    .B1(net2351),
    .B2(\i_seal.sealed_mono[21] ),
    .A2(\i_seal.sealed_crc[13] ),
    .A1(net2490));
 sg13g2_a21oi_1 _11356_ (.A1(_03739_),
    .A2(_03740_),
    .Y(_03741_),
    .B1(net2004));
 sg13g2_a221oi_1 _11357_ (.B2(\i_wdt.counter[21] ),
    .C1(_03741_),
    .B1(net2119),
    .A1(\timer_count[21] ),
    .Y(_03742_),
    .A2(net2124));
 sg13g2_a22oi_1 _11358_ (.Y(_03743_),
    .B1(_03738_),
    .B2(_03742_),
    .A2(_03737_),
    .A1(_03733_));
 sg13g2_o21ai_1 _11359_ (.B1(_03732_),
    .Y(_03744_),
    .A1(net2175),
    .A2(_03743_));
 sg13g2_o21ai_1 _11360_ (.B1(_03744_),
    .Y(_03745_),
    .A1(_03724_),
    .A2(_03727_));
 sg13g2_o21ai_1 _11361_ (.B1(_03415_),
    .Y(_03746_),
    .A1(net2435),
    .A2(_03745_));
 sg13g2_o21ai_1 _11362_ (.B1(_03416_),
    .Y(_03747_),
    .A1(_03711_),
    .A2(_03746_));
 sg13g2_nand3_1 _11363_ (.B(_03653_),
    .C(_03747_),
    .A(_03142_),
    .Y(_03748_));
 sg13g2_o21ai_1 _11364_ (.B1(_03748_),
    .Y(_03749_),
    .A1(_03142_),
    .A2(_03625_));
 sg13g2_mux2_1 _11365_ (.A0(net1815),
    .A1(net5168),
    .S(_03150_),
    .X(_00067_));
 sg13g2_nor2_1 _11366_ (.A(_01968_),
    .B(_03626_),
    .Y(_03750_));
 sg13g2_xnor2_1 _11367_ (.Y(_03751_),
    .A(_01968_),
    .B(_03626_));
 sg13g2_xnor2_1 _11368_ (.Y(_03752_),
    .A(_01971_),
    .B(_03358_));
 sg13g2_inv_1 _11369_ (.Y(_03753_),
    .A(_03752_));
 sg13g2_a21o_1 _11370_ (.A2(_03355_),
    .A1(\i_tinyqv.cpu.instr_data_start[13] ),
    .B1(\i_tinyqv.cpu.instr_data_start[14] ),
    .X(_03754_));
 sg13g2_nand2_1 _11371_ (.Y(_03755_),
    .A(_03356_),
    .B(_03754_));
 sg13g2_xnor2_1 _11372_ (.Y(_03756_),
    .A(net2571),
    .B(_03353_));
 sg13g2_nor2_1 _11373_ (.A(net2379),
    .B(_03756_),
    .Y(_03757_));
 sg13g2_xnor2_1 _11374_ (.Y(_03758_),
    .A(_01977_),
    .B(_03350_));
 sg13g2_nor2_1 _11375_ (.A(_02544_),
    .B(_03758_),
    .Y(_03759_));
 sg13g2_xnor2_1 _11376_ (.Y(_03760_),
    .A(_03346_),
    .B(_03347_));
 sg13g2_nor2_1 _11377_ (.A(_02539_),
    .B(_03760_),
    .Y(_03761_));
 sg13g2_nor3_1 _11378_ (.A(_03757_),
    .B(_03759_),
    .C(_03761_),
    .Y(_03762_));
 sg13g2_o21ai_1 _11379_ (.B1(_03762_),
    .Y(_03763_),
    .A1(net2371),
    .A2(_03755_));
 sg13g2_a22oi_1 _11380_ (.Y(_03764_),
    .B1(_03763_),
    .B2(net2437),
    .A2(_03753_),
    .A1(net2323));
 sg13g2_o21ai_1 _11381_ (.B1(_03764_),
    .Y(_03765_),
    .A1(_02551_),
    .A2(_03751_));
 sg13g2_mux2_1 _11382_ (.A0(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .S(net2316),
    .X(_03766_));
 sg13g2_a22oi_1 _11383_ (.Y(_03767_),
    .B1(_03403_),
    .B2(_03766_),
    .A2(_03400_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[2] ));
 sg13g2_nand2_1 _11384_ (.Y(_03768_),
    .A(net2318),
    .B(net2315));
 sg13g2_a22oi_1 _11385_ (.Y(_03769_),
    .B1(_03768_),
    .B2(_03395_),
    .A2(_03402_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[2] ));
 sg13g2_nand2_1 _11386_ (.Y(_03770_),
    .A(_03392_),
    .B(_03401_));
 sg13g2_nor2_1 _11387_ (.A(net2318),
    .B(_03770_),
    .Y(_03771_));
 sg13g2_a22oi_1 _11388_ (.Y(_03772_),
    .B1(_03671_),
    .B2(_03381_),
    .A2(_03394_),
    .A1(\i_tinyqv.cpu.i_core.mie[2] ));
 sg13g2_a22oi_1 _11389_ (.Y(_03773_),
    .B1(_03771_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .A2(_03389_),
    .A1(\i_tinyqv.cpu.i_core.mepc[2] ));
 sg13g2_nand4_1 _11390_ (.B(_03769_),
    .C(_03772_),
    .A(_03767_),
    .Y(_03774_),
    .D(_03773_));
 sg13g2_a22oi_1 _11391_ (.Y(_03775_),
    .B1(_03774_),
    .B2(_03373_),
    .A2(_03765_),
    .A1(_02803_));
 sg13g2_nand2_1 _11392_ (.Y(_03776_),
    .A(_02804_),
    .B(_03775_));
 sg13g2_o21ai_1 _11393_ (.B1(_03776_),
    .Y(_03777_),
    .A1(_02640_),
    .A2(_02804_));
 sg13g2_nand2_1 _11394_ (.Y(_03778_),
    .A(_03138_),
    .B(_03777_));
 sg13g2_nor2b_1 _11395_ (.A(\i_latch_mem.data_out[10] ),
    .B_N(net2467),
    .Y(_03779_));
 sg13g2_nor3_1 _11396_ (.A(net2389),
    .B(net2380),
    .C(_03779_),
    .Y(_03780_));
 sg13g2_a22oi_1 _11397_ (.Y(_03781_),
    .B1(net2077),
    .B2(\i2c_config_out[10] ),
    .A2(net2080),
    .A1(\crc16_read[10] ));
 sg13g2_a22oi_1 _11398_ (.Y(_03782_),
    .B1(net2084),
    .B2(\i_i2c_peri.rx_has_data ),
    .A2(net2086),
    .A1(\i_rtc.seconds_out[10] ));
 sg13g2_nand2_1 _11399_ (.Y(_03783_),
    .A(\timer_count[10] ),
    .B(net2121));
 sg13g2_a22oi_1 _11400_ (.Y(_03784_),
    .B1(net2345),
    .B2(\i_seal.sealed_value[10] ),
    .A2(\i_seal.sealed_crc[2] ),
    .A1(net2488));
 sg13g2_o21ai_1 _11401_ (.B1(_03784_),
    .Y(_03785_),
    .A1(_01937_),
    .A2(net2310));
 sg13g2_a221oi_1 _11402_ (.B2(_03785_),
    .C1(net2177),
    .B1(_03456_),
    .A1(\i_wdt.counter[10] ),
    .Y(_03786_),
    .A2(net2116));
 sg13g2_nand4_1 _11403_ (.B(_03782_),
    .C(_03783_),
    .A(_03781_),
    .Y(_03787_),
    .D(_03786_));
 sg13g2_nand2b_1 _11404_ (.Y(_03788_),
    .B(net2467),
    .A_N(\i_latch_mem.data_out[2] ));
 sg13g2_a22oi_1 _11405_ (.Y(_03789_),
    .B1(net2347),
    .B2(\i_seal.sealed_value[2] ),
    .A2(net2350),
    .A1(\i_seal.sealed_mono[2] ));
 sg13g2_nor2_1 _11406_ (.A(net2002),
    .B(_03789_),
    .Y(_03790_));
 sg13g2_a221oi_1 _11407_ (.B2(\i_wdt.counter[2] ),
    .C1(_03790_),
    .B1(net2117),
    .A1(\timer_count[2] ),
    .Y(_03791_),
    .A2(net2122));
 sg13g2_nand2_1 _11408_ (.Y(_03792_),
    .A(\i2c_data_out[2] ),
    .B(net2084));
 sg13g2_a22oi_1 _11409_ (.Y(_03793_),
    .B1(net2076),
    .B2(\i_uart_rx.recieved_data[2] ),
    .A2(net2082),
    .A1(\i_spi.data[2] ));
 sg13g2_a22oi_1 _11410_ (.Y(_03794_),
    .B1(net2081),
    .B2(\crc16_read[2] ),
    .A2(net2087),
    .A1(\i_rtc.seconds_out[2] ));
 sg13g2_a22oi_1 _11411_ (.Y(_03795_),
    .B1(net2078),
    .B2(\i2c_config_out[2] ),
    .A2(_03465_),
    .A1(\i_seal.commit_dropped ));
 sg13g2_a21oi_1 _11412_ (.A1(net4),
    .A2(_03470_),
    .Y(_03796_),
    .B1(net2174));
 sg13g2_a22oi_1 _11413_ (.Y(_03797_),
    .B1(_03453_),
    .B2(\gpio_out_sel[2] ),
    .A2(_03437_),
    .A1(uo_out[2]));
 sg13g2_and4_1 _11414_ (.A(_03794_),
    .B(_03795_),
    .C(_03796_),
    .D(_03797_),
    .X(_03798_));
 sg13g2_nand4_1 _11415_ (.B(_03792_),
    .C(_03793_),
    .A(_03791_),
    .Y(_03799_),
    .D(_03798_));
 sg13g2_nand3_1 _11416_ (.B(_03788_),
    .C(_03799_),
    .A(net2378),
    .Y(_03800_));
 sg13g2_nand2b_1 _11417_ (.Y(_03801_),
    .B(net2467),
    .A_N(\i_latch_mem.data_out[14] ));
 sg13g2_a22oi_1 _11418_ (.Y(_03802_),
    .B1(net2345),
    .B2(\i_seal.sealed_value[14] ),
    .A2(\i_seal.sealed_crc[6] ),
    .A1(net2488));
 sg13g2_o21ai_1 _11419_ (.B1(_03802_),
    .Y(_03803_),
    .A1(_01933_),
    .A2(net2310));
 sg13g2_a22oi_1 _11420_ (.Y(_03804_),
    .B1(net2118),
    .B2(\i_wdt.counter[14] ),
    .A2(net2123),
    .A1(\timer_count[14] ));
 sg13g2_a22oi_1 _11421_ (.Y(_03805_),
    .B1(_03803_),
    .B2(net2075),
    .A2(_03480_),
    .A1(\crc16_read[14] ));
 sg13g2_a22oi_1 _11422_ (.Y(_03806_),
    .B1(net2077),
    .B2(\i2c_config_out[14] ),
    .A2(net2085),
    .A1(\i_rtc.seconds_out[14] ));
 sg13g2_nand4_1 _11423_ (.B(_03804_),
    .C(_03805_),
    .A(_03434_),
    .Y(_03807_),
    .D(_03806_));
 sg13g2_nand3_1 _11424_ (.B(_03801_),
    .C(_03807_),
    .A(net2374),
    .Y(_03808_));
 sg13g2_a21oi_2 _11425_ (.B1(net2366),
    .Y(_03809_),
    .A2(_02076_),
    .A1(net2467));
 sg13g2_a221oi_1 _11426_ (.B2(net8),
    .C1(net2175),
    .B1(_03470_),
    .A1(\timer_count[6] ),
    .Y(_03810_),
    .A2(net2122));
 sg13g2_a22oi_1 _11427_ (.Y(_03811_),
    .B1(net2347),
    .B2(\i_seal.sealed_value[6] ),
    .A2(net2350),
    .A1(\i_seal.sealed_mono[6] ));
 sg13g2_nor2_1 _11428_ (.A(net2002),
    .B(_03811_),
    .Y(_03812_));
 sg13g2_a21oi_1 _11429_ (.A1(\i_wdt.counter[6] ),
    .A2(net2117),
    .Y(_03813_),
    .B1(_03812_));
 sg13g2_nand2_1 _11430_ (.Y(_03814_),
    .A(_03810_),
    .B(_03813_));
 sg13g2_a22oi_1 _11431_ (.Y(_03815_),
    .B1(net2076),
    .B2(\i_uart_rx.recieved_data[6] ),
    .A2(net2084),
    .A1(\i2c_data_out[6] ));
 sg13g2_a22oi_1 _11432_ (.Y(_03816_),
    .B1(net2079),
    .B2(\i2c_config_out[6] ),
    .A2(_03437_),
    .A1(uo_out[6]));
 sg13g2_a22oi_1 _11433_ (.Y(_03817_),
    .B1(_03453_),
    .B2(\gpio_out_sel[6] ),
    .A2(net2086),
    .A1(\i_rtc.seconds_out[6] ));
 sg13g2_a22oi_1 _11434_ (.Y(_03818_),
    .B1(net2080),
    .B2(\crc16_read[6] ),
    .A2(net2082),
    .A1(\i_spi.data[6] ));
 sg13g2_nand4_1 _11435_ (.B(_03816_),
    .C(_03817_),
    .A(_03815_),
    .Y(_03819_),
    .D(_03818_));
 sg13g2_o21ai_1 _11436_ (.B1(_03809_),
    .Y(_03820_),
    .A1(_03814_),
    .A2(_03819_));
 sg13g2_nand4_1 _11437_ (.B(_03800_),
    .C(_03808_),
    .A(net2388),
    .Y(_03821_),
    .D(_03820_));
 sg13g2_a21oi_1 _11438_ (.A1(_02077_),
    .A2(net1907),
    .Y(_03822_),
    .B1(net2379));
 sg13g2_o21ai_1 _11439_ (.B1(_03822_),
    .Y(_03823_),
    .A1(net2600),
    .A2(net1907));
 sg13g2_mux2_1 _11440_ (.A0(net2592),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net1908),
    .X(_03824_));
 sg13g2_mux2_1 _11441_ (.A0(net2600),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net1908),
    .X(_03825_));
 sg13g2_a22oi_1 _11442_ (.Y(_03826_),
    .B1(_03825_),
    .B2(net2377),
    .A2(_03824_),
    .A1(net2368));
 sg13g2_a21oi_1 _11443_ (.A1(_02078_),
    .A2(net1907),
    .Y(_03827_),
    .B1(net2371));
 sg13g2_o21ai_1 _11444_ (.B1(_03827_),
    .Y(_03828_),
    .A1(net2592),
    .A2(net1907));
 sg13g2_nand4_1 _11445_ (.B(_03823_),
    .C(_03826_),
    .A(net2390),
    .Y(_03829_),
    .D(_03828_));
 sg13g2_a221oi_1 _11446_ (.B2(_03829_),
    .C1(net2535),
    .B1(_03821_),
    .A1(_03780_),
    .Y(_03830_),
    .A2(_03787_));
 sg13g2_a221oi_1 _11447_ (.B2(\pps_count[14] ),
    .C1(net2176),
    .B1(net2073),
    .A1(\i_rtc.seconds_out[30] ),
    .Y(_03831_),
    .A2(net2089));
 sg13g2_nand2_1 _11448_ (.Y(_03832_),
    .A(\i_seal.sealed_sid[6] ),
    .B(net2348));
 sg13g2_a22oi_1 _11449_ (.Y(_03833_),
    .B1(net2342),
    .B2(\i_seal.sealed_value[30] ),
    .A2(\i_seal.sealed_mono[30] ),
    .A1(net2491));
 sg13g2_a21oi_2 _11450_ (.B1(net2003),
    .Y(_03834_),
    .A2(_03833_),
    .A1(_03832_));
 sg13g2_a221oi_1 _11451_ (.B2(\i_wdt.counter[30] ),
    .C1(_03834_),
    .B1(net2120),
    .A1(\timer_count[30] ),
    .Y(_03835_),
    .A2(net2125));
 sg13g2_a221oi_1 _11452_ (.B2(_03835_),
    .C1(net2371),
    .B1(_03831_),
    .A1(net2470),
    .Y(_03836_),
    .A2(_02080_));
 sg13g2_and2_1 _11453_ (.A(net2491),
    .B(\i_seal.sealed_mono[26] ),
    .X(_03837_));
 sg13g2_a221oi_1 _11454_ (.B2(\i_seal.sealed_value[26] ),
    .C1(_03837_),
    .B1(net2342),
    .A1(\i_seal.sealed_sid[2] ),
    .Y(_03838_),
    .A2(net2348));
 sg13g2_a221oi_1 _11455_ (.B2(\i_wdt.counter[26] ),
    .C1(net2176),
    .B1(net2119),
    .A1(\timer_count[26] ),
    .Y(_03839_),
    .A2(net2124));
 sg13g2_nor2b_1 _11456_ (.A(_03838_),
    .B_N(net2075),
    .Y(_03840_));
 sg13g2_a221oi_1 _11457_ (.B2(\pps_count[10] ),
    .C1(_03840_),
    .B1(net2072),
    .A1(\i_rtc.seconds_out[26] ),
    .Y(_03841_),
    .A2(net2088));
 sg13g2_a221oi_1 _11458_ (.B2(_03841_),
    .C1(net2380),
    .B1(_03839_),
    .A1(net2470),
    .Y(_03842_),
    .A2(_02079_));
 sg13g2_nor3_1 _11459_ (.A(_02470_),
    .B(_03836_),
    .C(_03842_),
    .Y(_03843_));
 sg13g2_mux2_1 _11460_ (.A0(net2600),
    .A1(\i_tinyqv.mem.qspi_data_buf[26] ),
    .S(_03133_),
    .X(_03844_));
 sg13g2_mux2_1 _11461_ (.A0(net2593),
    .A1(\i_tinyqv.mem.qspi_data_buf[30] ),
    .S(_03133_),
    .X(_03845_));
 sg13g2_a221oi_1 _11462_ (.B2(net2374),
    .C1(net2388),
    .B1(_03845_),
    .A1(net2382),
    .Y(_03846_),
    .A2(_03844_));
 sg13g2_a221oi_1 _11463_ (.B2(\pps_count[6] ),
    .C1(_01989_),
    .B1(net2072),
    .A1(\i_rtc.seconds_out[22] ),
    .Y(_03847_),
    .A2(net2088));
 sg13g2_nand2_1 _11464_ (.Y(_03848_),
    .A(net2490),
    .B(\i_seal.sealed_crc[14] ));
 sg13g2_a22oi_1 _11465_ (.Y(_03849_),
    .B1(net2343),
    .B2(\i_seal.sealed_value[22] ),
    .A2(net2349),
    .A1(\i_seal.sealed_mono[22] ));
 sg13g2_a21oi_1 _11466_ (.A1(_03848_),
    .A2(_03849_),
    .Y(_03850_),
    .B1(net2004));
 sg13g2_a221oi_1 _11467_ (.B2(\i_wdt.counter[22] ),
    .C1(_03850_),
    .B1(net2119),
    .A1(\timer_count[22] ),
    .Y(_03851_),
    .A2(net2124));
 sg13g2_a221oi_1 _11468_ (.B2(\pps_count[2] ),
    .C1(net2542),
    .B1(net2072),
    .A1(\i_rtc.seconds_out[18] ),
    .Y(_03852_),
    .A2(net2088));
 sg13g2_nand2_1 _11469_ (.Y(_03853_),
    .A(\i_seal.sealed_value[18] ),
    .B(net2343));
 sg13g2_a22oi_1 _11470_ (.Y(_03854_),
    .B1(net2350),
    .B2(\i_seal.sealed_mono[18] ),
    .A2(\i_seal.sealed_crc[10] ),
    .A1(net2492));
 sg13g2_a21oi_2 _11471_ (.B1(net2003),
    .Y(_03855_),
    .A2(_03854_),
    .A1(_03853_));
 sg13g2_a221oi_1 _11472_ (.B2(\i_wdt.counter[18] ),
    .C1(_03855_),
    .B1(net2120),
    .A1(\timer_count[18] ),
    .Y(_03856_),
    .A2(net2125));
 sg13g2_a22oi_1 _11473_ (.Y(_03857_),
    .B1(_03852_),
    .B2(_03856_),
    .A2(_03851_),
    .A1(_03847_));
 sg13g2_or2_1 _11474_ (.X(_03858_),
    .B(\i_tinyqv.mem.data_from_read[18] ),
    .A(net2539));
 sg13g2_o21ai_1 _11475_ (.B1(_03858_),
    .Y(_03859_),
    .A1(net2438),
    .A2(\i_tinyqv.mem.data_from_read[22] ));
 sg13g2_and2_1 _11476_ (.A(net2541),
    .B(\i_latch_mem.data_out[22] ),
    .X(_03860_));
 sg13g2_a21oi_1 _11477_ (.A1(net2438),
    .A2(\i_latch_mem.data_out[18] ),
    .Y(_03861_),
    .B1(_03860_));
 sg13g2_a221oi_1 _11478_ (.B2(net2469),
    .C1(net2537),
    .B1(_03861_),
    .A1(net2389),
    .Y(_03862_),
    .A2(_03859_));
 sg13g2_o21ai_1 _11479_ (.B1(_03862_),
    .Y(_03863_),
    .A1(net2175),
    .A2(_03857_));
 sg13g2_o21ai_1 _11480_ (.B1(_03863_),
    .Y(_03864_),
    .A1(_03843_),
    .A2(_03846_));
 sg13g2_o21ai_1 _11481_ (.B1(_03415_),
    .Y(_03865_),
    .A1(net2436),
    .A2(_03864_));
 sg13g2_o21ai_1 _11482_ (.B1(_03416_),
    .Y(_03866_),
    .A1(_03830_),
    .A2(_03865_));
 sg13g2_nand2_1 _11483_ (.Y(_03867_),
    .A(_03778_),
    .B(_03866_));
 sg13g2_xnor2_1 _11484_ (.Y(_03868_),
    .A(_02745_),
    .B(_02747_));
 sg13g2_nand2_1 _11485_ (.Y(_03869_),
    .A(_03153_),
    .B(_03868_));
 sg13g2_o21ai_1 _11486_ (.B1(_02780_),
    .Y(_03870_),
    .A1(net2529),
    .A2(_02781_));
 sg13g2_a22oi_1 _11487_ (.Y(_03871_),
    .B1(_03157_),
    .B2(_03870_),
    .A2(_03156_),
    .A1(_02782_));
 sg13g2_nand2_1 _11488_ (.Y(_03872_),
    .A(_02870_),
    .B(_02871_));
 sg13g2_nand3_1 _11489_ (.B(_03144_),
    .C(_03872_),
    .A(_02872_),
    .Y(_03873_));
 sg13g2_nand4_1 _11490_ (.B(_03869_),
    .C(_03871_),
    .A(_03167_),
    .Y(_03874_),
    .D(_03873_));
 sg13g2_nor2_1 _11491_ (.A(net2434),
    .B(_03595_),
    .Y(_03875_));
 sg13g2_nor2_1 _11492_ (.A(net2524),
    .B(_03621_),
    .Y(_03876_));
 sg13g2_o21ai_1 _11493_ (.B1(_03166_),
    .Y(_03877_),
    .A1(_03875_),
    .A2(_03876_));
 sg13g2_nand3_1 _11494_ (.B(_03874_),
    .C(_03877_),
    .A(_03342_),
    .Y(_03878_));
 sg13g2_a21oi_1 _11495_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .A2(_03152_),
    .Y(_03879_),
    .B1(_03142_));
 sg13g2_a22oi_1 _11496_ (.Y(_03880_),
    .B1(_03878_),
    .B2(_03879_),
    .A2(_03867_),
    .A1(_03142_));
 sg13g2_mux2_1 _11497_ (.A0(net1798),
    .A1(net5242),
    .S(_03150_),
    .X(_00068_));
 sg13g2_and2_1 _11498_ (.A(\gpio_out[7] ),
    .B(\gpio_out_sel[7] ),
    .X(uo_out[7]));
 sg13g2_xnor2_1 _11499_ (.Y(_03881_),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .B(_03750_));
 sg13g2_xnor2_1 _11500_ (.Y(_03882_),
    .A(_01972_),
    .B(_03356_));
 sg13g2_xnor2_1 _11501_ (.Y(_03883_),
    .A(net2572),
    .B(_03351_));
 sg13g2_xor2_1 _11502_ (.B(_03348_),
    .A(net2575),
    .X(_03884_));
 sg13g2_inv_1 _11503_ (.Y(_03885_),
    .A(_03884_));
 sg13g2_a221oi_1 _11504_ (.B2(net2377),
    .C1(net2533),
    .B1(_03885_),
    .A1(net2369),
    .Y(_03886_),
    .A2(_03883_));
 sg13g2_a21o_1 _11505_ (.A2(_03353_),
    .A1(net2571),
    .B1(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(_03887_));
 sg13g2_nand2_1 _11506_ (.Y(_03888_),
    .A(_03354_),
    .B(_03887_));
 sg13g2_a22oi_1 _11507_ (.Y(_03889_),
    .B1(_03888_),
    .B2(net2382),
    .A2(_03882_),
    .A1(net2373));
 sg13g2_xnor2_1 _11508_ (.Y(_03890_),
    .A(\i_tinyqv.cpu.instr_data_start[19] ),
    .B(_03359_));
 sg13g2_inv_1 _11509_ (.Y(_03891_),
    .A(_03890_));
 sg13g2_a22oi_1 _11510_ (.Y(_03892_),
    .B1(_03891_),
    .B2(net2323),
    .A2(_03889_),
    .A1(_03886_));
 sg13g2_o21ai_1 _11511_ (.B1(_03892_),
    .Y(_03893_),
    .A1(_02551_),
    .A2(_03881_));
 sg13g2_nor2_1 _11512_ (.A(net2321),
    .B(_03770_),
    .Y(_03894_));
 sg13g2_nand2_1 _11513_ (.Y(_03895_),
    .A(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .B(net2316));
 sg13g2_o21ai_1 _11514_ (.B1(_03895_),
    .Y(_03896_),
    .A1(_01961_),
    .A2(net2316));
 sg13g2_nand2_1 _11515_ (.Y(_03897_),
    .A(\i_tinyqv.cpu.i_core.mepc[3] ),
    .B(_03389_));
 sg13g2_a22oi_1 _11516_ (.Y(_03898_),
    .B1(_02769_),
    .B2(\i_tinyqv.cpu.i_core.mcause[4] ),
    .A2(net2320),
    .A1(\i_tinyqv.cpu.i_core.mcause[3] ));
 sg13g2_nor3_1 _11517_ (.A(_03377_),
    .B(_03396_),
    .C(_03898_),
    .Y(_03899_));
 sg13g2_a22oi_1 _11518_ (.Y(_03900_),
    .B1(net2322),
    .B2(\i_tinyqv.cpu.i_core.mie[4] ),
    .A2(net2324),
    .A1(\i_tinyqv.cpu.i_core.mie[3] ));
 sg13g2_nor2_1 _11519_ (.A(_03393_),
    .B(_03900_),
    .Y(_03901_));
 sg13g2_a221oi_1 _11520_ (.B2(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .C1(_03901_),
    .B1(_03771_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .Y(_03902_),
    .A2(_03400_));
 sg13g2_nand3_1 _11521_ (.B(net2322),
    .C(_03894_),
    .A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .Y(_03903_));
 sg13g2_a221oi_1 _11522_ (.B2(_03896_),
    .C1(_03899_),
    .B1(_03403_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .Y(_03904_),
    .A2(_03402_));
 sg13g2_nand4_1 _11523_ (.B(_03902_),
    .C(_03903_),
    .A(_03897_),
    .Y(_03905_),
    .D(_03904_));
 sg13g2_a22oi_1 _11524_ (.Y(_03906_),
    .B1(_03905_),
    .B2(_03373_),
    .A2(_03893_),
    .A1(_02803_));
 sg13g2_mux2_1 _11525_ (.A0(_02571_),
    .A1(_03906_),
    .S(_02804_),
    .X(_03907_));
 sg13g2_nand2_1 _11526_ (.Y(_03908_),
    .A(_03138_),
    .B(_03907_));
 sg13g2_o21ai_1 _11527_ (.B1(net2374),
    .Y(_03909_),
    .A1(net2590),
    .A2(net1906));
 sg13g2_a21oi_1 _11528_ (.A1(_02083_),
    .A2(net1906),
    .Y(_03910_),
    .B1(_03909_));
 sg13g2_mux2_1 _11529_ (.A0(net2590),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(_03417_),
    .X(_03911_));
 sg13g2_a21oi_1 _11530_ (.A1(_02037_),
    .A2(_03417_),
    .Y(_03912_),
    .B1(_02539_));
 sg13g2_o21ai_1 _11531_ (.B1(_03912_),
    .Y(_03913_),
    .A1(net2598),
    .A2(_03417_));
 sg13g2_a21oi_1 _11532_ (.A1(_02082_),
    .A2(net1906),
    .Y(_03914_),
    .B1(net2379));
 sg13g2_o21ai_1 _11533_ (.B1(_03914_),
    .Y(_03915_),
    .A1(net2598),
    .A2(net1906));
 sg13g2_a21oi_1 _11534_ (.A1(net2369),
    .A2(_03911_),
    .Y(_03916_),
    .B1(_03910_));
 sg13g2_nand4_1 _11535_ (.B(_03913_),
    .C(_03915_),
    .A(net2390),
    .Y(_03917_),
    .D(_03916_));
 sg13g2_nand2b_1 _11536_ (.Y(_03918_),
    .B(net2468),
    .A_N(\i_latch_mem.data_out[11] ));
 sg13g2_a22oi_1 _11537_ (.Y(_03919_),
    .B1(net2077),
    .B2(\i2c_config_out[11] ),
    .A2(net2086),
    .A1(\i_rtc.seconds_out[11] ));
 sg13g2_a22oi_1 _11538_ (.Y(_03920_),
    .B1(net2346),
    .B2(\i_seal.sealed_value[11] ),
    .A2(\i_seal.sealed_crc[3] ),
    .A1(net2489));
 sg13g2_o21ai_1 _11539_ (.B1(_03920_),
    .Y(_03921_),
    .A1(_01936_),
    .A2(_03458_));
 sg13g2_a22oi_1 _11540_ (.Y(_03922_),
    .B1(_03456_),
    .B2(_03921_),
    .A2(net2084),
    .A1(\i_i2c_peri.tx_pending ));
 sg13g2_nand2_1 _11541_ (.Y(_03923_),
    .A(\i_wdt.counter[11] ),
    .B(net2116));
 sg13g2_a221oi_1 _11542_ (.B2(\crc16_read[11] ),
    .C1(net2174),
    .B1(net2081),
    .A1(\timer_count[11] ),
    .Y(_03924_),
    .A2(net2121));
 sg13g2_nand4_1 _11543_ (.B(_03922_),
    .C(_03923_),
    .A(_03919_),
    .Y(_03925_),
    .D(_03924_));
 sg13g2_nand3_1 _11544_ (.B(_03918_),
    .C(_03925_),
    .A(net2384),
    .Y(_03926_));
 sg13g2_nand2b_1 _11545_ (.Y(_03927_),
    .B(net2468),
    .A_N(\i_latch_mem.data_out[3] ));
 sg13g2_a221oi_1 _11546_ (.B2(net5),
    .C1(net2175),
    .B1(_03470_),
    .A1(\i_wdt.counter[3] ),
    .Y(_03928_),
    .A2(net2116));
 sg13g2_a22oi_1 _11547_ (.Y(_03929_),
    .B1(net2345),
    .B2(\i_seal.sealed_value[3] ),
    .A2(net2351),
    .A1(\i_seal.sealed_mono[3] ));
 sg13g2_nor2_2 _11548_ (.A(net2002),
    .B(_03929_),
    .Y(_03930_));
 sg13g2_a21oi_1 _11549_ (.A1(\timer_count[3] ),
    .A2(net2122),
    .Y(_03931_),
    .B1(_03930_));
 sg13g2_a22oi_1 _11550_ (.Y(_03932_),
    .B1(_03468_),
    .B2(\i_uart_rx.recieved_data[3] ),
    .A2(net2080),
    .A1(\crc16_read[3] ));
 sg13g2_a22oi_1 _11551_ (.Y(_03933_),
    .B1(net2079),
    .B2(\i2c_config_out[3] ),
    .A2(_03437_),
    .A1(uo_out[3]));
 sg13g2_a22oi_1 _11552_ (.Y(_03934_),
    .B1(_03453_),
    .B2(\gpio_out_sel[3] ),
    .A2(net2083),
    .A1(\i2c_data_out[3] ));
 sg13g2_a22oi_1 _11553_ (.Y(_03935_),
    .B1(_03446_),
    .B2(\i_spi.data[3] ),
    .A2(net2086),
    .A1(\i_rtc.seconds_out[3] ));
 sg13g2_and4_1 _11554_ (.A(_03932_),
    .B(_03933_),
    .C(_03934_),
    .D(_03935_),
    .X(_03936_));
 sg13g2_nand3_1 _11555_ (.B(_03931_),
    .C(_03936_),
    .A(_03928_),
    .Y(_03937_));
 sg13g2_nand3_1 _11556_ (.B(_03927_),
    .C(_03937_),
    .A(net2378),
    .Y(_03938_));
 sg13g2_nand2b_1 _11557_ (.Y(_03939_),
    .B(net2468),
    .A_N(\i_latch_mem.data_out[15] ));
 sg13g2_a22oi_1 _11558_ (.Y(_03940_),
    .B1(net2118),
    .B2(\i_wdt.counter[15] ),
    .A2(net2123),
    .A1(\timer_count[15] ));
 sg13g2_a22oi_1 _11559_ (.Y(_03941_),
    .B1(net2345),
    .B2(\i_seal.sealed_value[15] ),
    .A2(\i_seal.sealed_crc[7] ),
    .A1(net2488));
 sg13g2_o21ai_1 _11560_ (.B1(_03941_),
    .Y(_03942_),
    .A1(_01932_),
    .A2(net2310));
 sg13g2_a22oi_1 _11561_ (.Y(_03943_),
    .B1(net2077),
    .B2(\i2c_config_out[15] ),
    .A2(net2085),
    .A1(\i_rtc.seconds_out[15] ));
 sg13g2_a22oi_1 _11562_ (.Y(_03944_),
    .B1(_03942_),
    .B2(_03478_),
    .A2(_03480_),
    .A1(\crc16_read[15] ));
 sg13g2_nand4_1 _11563_ (.B(_03940_),
    .C(_03943_),
    .A(_03434_),
    .Y(_03945_),
    .D(_03944_));
 sg13g2_nand3_1 _11564_ (.B(_03939_),
    .C(_03945_),
    .A(net2375),
    .Y(_03946_));
 sg13g2_nand2b_1 _11565_ (.Y(_03947_),
    .B(net2468),
    .A_N(\i_latch_mem.data_out[7] ));
 sg13g2_a221oi_1 _11566_ (.B2(\i_uart_rx.recieved_data[7] ),
    .C1(net2174),
    .B1(net2076),
    .A1(\timer_count[7] ),
    .Y(_03948_),
    .A2(net2121));
 sg13g2_a22oi_1 _11567_ (.Y(_03949_),
    .B1(net2346),
    .B2(\i_seal.sealed_value[7] ),
    .A2(net2350),
    .A1(\i_seal.sealed_mono[7] ));
 sg13g2_nor2_1 _11568_ (.A(net2005),
    .B(_03949_),
    .Y(_03950_));
 sg13g2_a21oi_1 _11569_ (.A1(\i_wdt.counter[7] ),
    .A2(net2116),
    .Y(_03951_),
    .B1(_03950_));
 sg13g2_a22oi_1 _11570_ (.Y(_03952_),
    .B1(uo_out[7]),
    .B2(_03437_),
    .A2(net2086),
    .A1(\i_rtc.seconds_out[7] ));
 sg13g2_a22oi_1 _11571_ (.Y(_03953_),
    .B1(net2079),
    .B2(\i2c_config_out[7] ),
    .A2(net2083),
    .A1(\i2c_data_out[7] ));
 sg13g2_a22oi_1 _11572_ (.Y(_03954_),
    .B1(_03470_),
    .B2(net9),
    .A2(net2082),
    .A1(\i_spi.data[7] ));
 sg13g2_a22oi_1 _11573_ (.Y(_03955_),
    .B1(net2080),
    .B2(\crc16_read[7] ),
    .A2(_03453_),
    .A1(\gpio_out_sel[7] ));
 sg13g2_and4_1 _11574_ (.A(_03952_),
    .B(_03953_),
    .C(_03954_),
    .D(_03955_),
    .X(_03956_));
 sg13g2_nand3_1 _11575_ (.B(_03951_),
    .C(_03956_),
    .A(_03948_),
    .Y(_03957_));
 sg13g2_nand3_1 _11576_ (.B(_03947_),
    .C(_03957_),
    .A(net2369),
    .Y(_03958_));
 sg13g2_nand4_1 _11577_ (.B(_03938_),
    .C(_03946_),
    .A(_03926_),
    .Y(_03959_),
    .D(_03958_));
 sg13g2_nand3_1 _11578_ (.B(_03917_),
    .C(_03959_),
    .A(net2436),
    .Y(_03960_));
 sg13g2_nor2b_1 _11579_ (.A(net2541),
    .B_N(\i_latch_mem.data_out[19] ),
    .Y(_03961_));
 sg13g2_a21oi_1 _11580_ (.A1(net2542),
    .A2(\i_latch_mem.data_out[23] ),
    .Y(_03962_),
    .B1(_03961_));
 sg13g2_or2_1 _11581_ (.X(_03963_),
    .B(\i_tinyqv.mem.data_from_read[19] ),
    .A(net2539));
 sg13g2_o21ai_1 _11582_ (.B1(_03963_),
    .Y(_03964_),
    .A1(net2438),
    .A2(\i_tinyqv.mem.data_from_read[23] ));
 sg13g2_a221oi_1 _11583_ (.B2(net2390),
    .C1(_02547_),
    .B1(_03964_),
    .A1(net2472),
    .Y(_03965_),
    .A2(_03962_));
 sg13g2_a221oi_1 _11584_ (.B2(\pps_count[3] ),
    .C1(net2542),
    .B1(net2073),
    .A1(\i_rtc.seconds_out[19] ),
    .Y(_03966_),
    .A2(net2088));
 sg13g2_nand2_1 _11585_ (.Y(_03967_),
    .A(\i_seal.sealed_value[19] ),
    .B(net2343));
 sg13g2_a22oi_1 _11586_ (.Y(_03968_),
    .B1(net2351),
    .B2(\i_seal.sealed_mono[19] ),
    .A2(\i_seal.sealed_crc[11] ),
    .A1(net2492));
 sg13g2_a21oi_1 _11587_ (.A1(_03967_),
    .A2(_03968_),
    .Y(_03969_),
    .B1(net2004));
 sg13g2_a221oi_1 _11588_ (.B2(\i_wdt.counter[19] ),
    .C1(_03969_),
    .B1(net2119),
    .A1(\timer_count[19] ),
    .Y(_03970_),
    .A2(net2124));
 sg13g2_a221oi_1 _11589_ (.B2(\pps_count[7] ),
    .C1(_01989_),
    .B1(net2072),
    .A1(\i_rtc.seconds_out[23] ),
    .Y(_03971_),
    .A2(net2089));
 sg13g2_nand2_1 _11590_ (.Y(_03972_),
    .A(\i_seal.sealed_mono[23] ),
    .B(net2349));
 sg13g2_a22oi_1 _11591_ (.Y(_03973_),
    .B1(net2344),
    .B2(\i_seal.sealed_value[23] ),
    .A2(\i_seal.sealed_crc[15] ),
    .A1(net2490));
 sg13g2_a21oi_1 _11592_ (.A1(_03972_),
    .A2(_03973_),
    .Y(_03974_),
    .B1(net2004));
 sg13g2_a221oi_1 _11593_ (.B2(\i_wdt.counter[23] ),
    .C1(_03974_),
    .B1(net2119),
    .A1(\timer_count[23] ),
    .Y(_03975_),
    .A2(net2125));
 sg13g2_a22oi_1 _11594_ (.Y(_03976_),
    .B1(_03971_),
    .B2(_03975_),
    .A2(_03970_),
    .A1(_03966_));
 sg13g2_o21ai_1 _11595_ (.B1(_03965_),
    .Y(_03977_),
    .A1(net2175),
    .A2(_03976_));
 sg13g2_a22oi_1 _11596_ (.Y(_03978_),
    .B1(net2119),
    .B2(\i_wdt.counter[27] ),
    .A2(net2124),
    .A1(\timer_count[27] ));
 sg13g2_a22oi_1 _11597_ (.Y(_03979_),
    .B1(net2342),
    .B2(\i_seal.sealed_value[27] ),
    .A2(net2348),
    .A1(\i_seal.sealed_sid[3] ));
 sg13g2_o21ai_1 _11598_ (.B1(_03979_),
    .Y(_03980_),
    .A1(_01809_),
    .A2(_01930_));
 sg13g2_a21o_1 _11599_ (.A2(_03980_),
    .A1(net2075),
    .B1(net2176),
    .X(_03981_));
 sg13g2_a221oi_1 _11600_ (.B2(\pps_count[11] ),
    .C1(_03981_),
    .B1(net2073),
    .A1(\i_rtc.seconds_out[27] ),
    .Y(_03982_),
    .A2(net2089));
 sg13g2_a22oi_1 _11601_ (.Y(_03983_),
    .B1(_03978_),
    .B2(_03982_),
    .A2(_02084_),
    .A1(net2470));
 sg13g2_nor3_1 _11602_ (.A(\i_tinyqv.mem.qspi_data_buf[27] ),
    .B(net2387),
    .C(_03132_),
    .Y(_03984_));
 sg13g2_nor3_1 _11603_ (.A(net2598),
    .B(net2387),
    .C(_03133_),
    .Y(_03985_));
 sg13g2_nor3_1 _11604_ (.A(_02524_),
    .B(_03984_),
    .C(_03985_),
    .Y(_03986_));
 sg13g2_a21oi_1 _11605_ (.A1(net2591),
    .A2(_03132_),
    .Y(_03987_),
    .B1(net2388));
 sg13g2_o21ai_1 _11606_ (.B1(_03987_),
    .Y(_03988_),
    .A1(_02085_),
    .A2(_03132_));
 sg13g2_a221oi_1 _11607_ (.B2(\pps_count[15] ),
    .C1(net2176),
    .B1(net2074),
    .A1(\i_rtc.seconds_out[31] ),
    .Y(_03989_),
    .A2(net2089));
 sg13g2_nand2_1 _11608_ (.Y(_03990_),
    .A(\i_seal.sealed_sid[7] ),
    .B(net2348));
 sg13g2_a22oi_1 _11609_ (.Y(_03991_),
    .B1(net2342),
    .B2(\i_seal.sealed_value[31] ),
    .A2(\i_seal.sealed_mono[31] ),
    .A1(net2491));
 sg13g2_a21oi_2 _11610_ (.B1(net2003),
    .Y(_03992_),
    .A2(_03991_),
    .A1(_03990_));
 sg13g2_a221oi_1 _11611_ (.B2(\i_wdt.counter[31] ),
    .C1(_03992_),
    .B1(net2120),
    .A1(\timer_count[31] ),
    .Y(_03993_),
    .A2(net2125));
 sg13g2_a221oi_1 _11612_ (.B2(_03993_),
    .C1(net2316),
    .B1(_03989_),
    .A1(net2470),
    .Y(_03994_),
    .A2(_02086_));
 sg13g2_a22oi_1 _11613_ (.Y(_03995_),
    .B1(_03988_),
    .B2(_03994_),
    .A2(_03986_),
    .A1(_03983_));
 sg13g2_and3_2 _11614_ (.X(_03996_),
    .A(_03960_),
    .B(_03977_),
    .C(_03995_));
 sg13g2_o21ai_1 _11615_ (.B1(_03416_),
    .Y(_03997_),
    .A1(_03414_),
    .A2(_03996_));
 sg13g2_nand2_1 _11616_ (.Y(_03998_),
    .A(_03908_),
    .B(_03997_));
 sg13g2_a21oi_1 _11617_ (.A1(_02872_),
    .A2(_02874_),
    .Y(_03999_),
    .B1(_03145_));
 sg13g2_nand2b_1 _11618_ (.Y(_04000_),
    .B(_03999_),
    .A_N(_02875_));
 sg13g2_nand2_1 _11619_ (.Y(_04001_),
    .A(_02748_),
    .B(_02749_));
 sg13g2_nor2_1 _11620_ (.A(_02750_),
    .B(_03154_),
    .Y(_04002_));
 sg13g2_o21ai_1 _11621_ (.B1(_02778_),
    .Y(_04003_),
    .A1(net2529),
    .A2(_02777_));
 sg13g2_nor2b_1 _11622_ (.A(_02779_),
    .B_N(_03156_),
    .Y(_04004_));
 sg13g2_a221oi_1 _11623_ (.B2(_03157_),
    .C1(_04004_),
    .B1(_04003_),
    .A1(_04001_),
    .Y(_04005_),
    .A2(_04002_));
 sg13g2_nand3_1 _11624_ (.B(_04000_),
    .C(_04005_),
    .A(_03167_),
    .Y(_04006_));
 sg13g2_nor3_1 _11625_ (.A(net2523),
    .B(_03179_),
    .C(_03337_),
    .Y(_04007_));
 sg13g2_a21oi_1 _11626_ (.A1(net2521),
    .A2(_03281_),
    .Y(_04008_),
    .B1(_04007_));
 sg13g2_nand2_1 _11627_ (.Y(_04009_),
    .A(_03166_),
    .B(_04008_));
 sg13g2_nand3_1 _11628_ (.B(_04006_),
    .C(_04009_),
    .A(_03342_),
    .Y(_04010_));
 sg13g2_a21oi_1 _11629_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A2(_03152_),
    .Y(_04011_),
    .B1(_03142_));
 sg13g2_a22oi_1 _11630_ (.Y(_04012_),
    .B1(_04010_),
    .B2(_04011_),
    .A2(_03998_),
    .A1(_03142_));
 sg13g2_mux2_1 _11631_ (.A0(net1796),
    .A1(net4988),
    .S(_03150_),
    .X(_00069_));
 sg13g2_nor2b_2 _11632_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .Y(_04013_));
 sg13g2_nand4_1 _11633_ (.B(net2504),
    .C(net1889),
    .A(net2505),
    .Y(_04014_),
    .D(_04013_));
 sg13g2_mux2_1 _11634_ (.A0(net1817),
    .A1(net5243),
    .S(_04014_),
    .X(_00062_));
 sg13g2_mux2_1 _11635_ (.A0(net1815),
    .A1(net5043),
    .S(_04014_),
    .X(_00063_));
 sg13g2_mux2_1 _11636_ (.A0(net1799),
    .A1(net4956),
    .S(_04014_),
    .X(_00064_));
 sg13g2_mux2_1 _11637_ (.A0(net1796),
    .A1(net5082),
    .S(_04014_),
    .X(_00065_));
 sg13g2_nor2b_2 _11638_ (.A(net4105),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .Y(_04015_));
 sg13g2_nand4_1 _11639_ (.B(net2504),
    .C(net1889),
    .A(net2505),
    .Y(_04016_),
    .D(_04015_));
 sg13g2_mux2_1 _11640_ (.A0(net1816),
    .A1(net5048),
    .S(_04016_),
    .X(_00058_));
 sg13g2_mux2_1 _11641_ (.A0(net1814),
    .A1(net4983),
    .S(_04016_),
    .X(_00059_));
 sg13g2_mux2_1 _11642_ (.A0(net1799),
    .A1(net4847),
    .S(_04016_),
    .X(_00060_));
 sg13g2_mux2_1 _11643_ (.A0(net1796),
    .A1(net4876),
    .S(_04016_),
    .X(_00061_));
 sg13g2_nor2_2 _11644_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .B(net4105),
    .Y(_04017_));
 sg13g2_and4_1 _11645_ (.A(net2505),
    .B(net2504),
    .C(net1889),
    .D(_04017_),
    .X(_04018_));
 sg13g2_mux2_1 _11646_ (.A0(net5039),
    .A1(net1816),
    .S(_04018_),
    .X(_00054_));
 sg13g2_mux2_1 _11647_ (.A0(net4959),
    .A1(net1814),
    .S(_04018_),
    .X(_00055_));
 sg13g2_mux2_1 _11648_ (.A0(net5023),
    .A1(net1798),
    .S(_04018_),
    .X(_00056_));
 sg13g2_mux2_1 _11649_ (.A0(net4967),
    .A1(net1797),
    .S(_04018_),
    .X(_00057_));
 sg13g2_nand2_1 _11650_ (.Y(_04019_),
    .A(net2504),
    .B(net1889));
 sg13g2_nor2_2 _11651_ (.A(net2505),
    .B(_04019_),
    .Y(_04020_));
 sg13g2_nand2_2 _11652_ (.Y(_04021_),
    .A(_03148_),
    .B(_04020_));
 sg13g2_nor2_1 _11653_ (.A(net1816),
    .B(_04021_),
    .Y(_04022_));
 sg13g2_a21oi_1 _11654_ (.A1(_01999_),
    .A2(_04021_),
    .Y(_00050_),
    .B1(_04022_));
 sg13g2_mux2_1 _11655_ (.A0(net1814),
    .A1(net5000),
    .S(_04021_),
    .X(_00051_));
 sg13g2_mux2_1 _11656_ (.A0(net1799),
    .A1(net5022),
    .S(_04021_),
    .X(_00052_));
 sg13g2_mux2_1 _11657_ (.A0(net1796),
    .A1(net4902),
    .S(_04021_),
    .X(_00053_));
 sg13g2_nand2_2 _11658_ (.Y(_04023_),
    .A(_04013_),
    .B(_04020_));
 sg13g2_mux2_1 _11659_ (.A0(net1817),
    .A1(net5203),
    .S(_04023_),
    .X(_00046_));
 sg13g2_mux2_1 _11660_ (.A0(net1815),
    .A1(net5208),
    .S(_04023_),
    .X(_00047_));
 sg13g2_mux2_1 _11661_ (.A0(net1799),
    .A1(net5164),
    .S(_04023_),
    .X(_00048_));
 sg13g2_mux2_1 _11662_ (.A0(net1796),
    .A1(net5133),
    .S(_04023_),
    .X(_00049_));
 sg13g2_nand2_2 _11663_ (.Y(_04024_),
    .A(_04015_),
    .B(_04020_));
 sg13g2_mux2_1 _11664_ (.A0(net1817),
    .A1(net5228),
    .S(_04024_),
    .X(_00094_));
 sg13g2_mux2_1 _11665_ (.A0(net1815),
    .A1(net5166),
    .S(_04024_),
    .X(_00095_));
 sg13g2_mux2_1 _11666_ (.A0(net1798),
    .A1(net5170),
    .S(_04024_),
    .X(_00096_));
 sg13g2_mux2_1 _11667_ (.A0(net1796),
    .A1(net4957),
    .S(_04024_),
    .X(_00097_));
 sg13g2_nand2_2 _11668_ (.Y(_04025_),
    .A(_04017_),
    .B(_04020_));
 sg13g2_mux2_1 _11669_ (.A0(net1817),
    .A1(net5165),
    .S(_04025_),
    .X(_00090_));
 sg13g2_mux2_1 _11670_ (.A0(net1814),
    .A1(net5171),
    .S(_04025_),
    .X(_00091_));
 sg13g2_mux2_1 _11671_ (.A0(net1799),
    .A1(net5221),
    .S(_04025_),
    .X(_00092_));
 sg13g2_mux2_1 _11672_ (.A0(net1797),
    .A1(net4678),
    .S(_04025_),
    .X(_00093_));
 sg13g2_nor2b_1 _11673_ (.A(net2504),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .Y(_04026_));
 sg13g2_nand3_1 _11674_ (.B(_03148_),
    .C(_04026_),
    .A(net1889),
    .Y(_04027_));
 sg13g2_mux2_1 _11675_ (.A0(net1816),
    .A1(net4989),
    .S(_04027_),
    .X(_00086_));
 sg13g2_mux2_1 _11676_ (.A0(net1814),
    .A1(net4807),
    .S(_04027_),
    .X(_00087_));
 sg13g2_mux2_1 _11677_ (.A0(net1798),
    .A1(net4968),
    .S(_04027_),
    .X(_00088_));
 sg13g2_mux2_1 _11678_ (.A0(net1797),
    .A1(net4980),
    .S(_04027_),
    .X(_00089_));
 sg13g2_nand3_1 _11679_ (.B(_04013_),
    .C(_04026_),
    .A(net1889),
    .Y(_04028_));
 sg13g2_nor2_1 _11680_ (.A(net1816),
    .B(_04028_),
    .Y(_04029_));
 sg13g2_a21oi_1 _11681_ (.A1(_02000_),
    .A2(_04028_),
    .Y(_00082_),
    .B1(_04029_));
 sg13g2_mux2_1 _11682_ (.A0(net1814),
    .A1(net4774),
    .S(_04028_),
    .X(_00083_));
 sg13g2_mux2_1 _11683_ (.A0(net1798),
    .A1(net4969),
    .S(_04028_),
    .X(_00084_));
 sg13g2_mux2_1 _11684_ (.A0(net1796),
    .A1(net4768),
    .S(_04028_),
    .X(_00085_));
 sg13g2_nand3_1 _11685_ (.B(_04015_),
    .C(_04026_),
    .A(_03147_),
    .Y(_04030_));
 sg13g2_mux2_1 _11686_ (.A0(net1816),
    .A1(net4987),
    .S(_04030_),
    .X(_00078_));
 sg13g2_mux2_1 _11687_ (.A0(net1814),
    .A1(net4706),
    .S(_04030_),
    .X(_00079_));
 sg13g2_mux2_1 _11688_ (.A0(net1798),
    .A1(net4901),
    .S(_04030_),
    .X(_00080_));
 sg13g2_mux2_1 _11689_ (.A0(net1796),
    .A1(net4837),
    .S(_04030_),
    .X(_00081_));
 sg13g2_nor2_1 _11690_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .B(net5382),
    .Y(_04031_));
 sg13g2_nand3_1 _11691_ (.B(_04013_),
    .C(_04031_),
    .A(net1889),
    .Y(_04032_));
 sg13g2_mux2_1 _11692_ (.A0(net1817),
    .A1(net5059),
    .S(_04032_),
    .X(_00074_));
 sg13g2_mux2_1 _11693_ (.A0(net1815),
    .A1(net4836),
    .S(_04032_),
    .X(_00075_));
 sg13g2_mux2_1 _11694_ (.A0(net1798),
    .A1(net4884),
    .S(_04032_),
    .X(_00076_));
 sg13g2_mux2_1 _11695_ (.A0(net1797),
    .A1(net4769),
    .S(_04032_),
    .X(_00077_));
 sg13g2_nand3_1 _11696_ (.B(_04015_),
    .C(net5383),
    .A(_03147_),
    .Y(_04033_));
 sg13g2_mux2_1 _11697_ (.A0(net1816),
    .A1(net4904),
    .S(_04033_),
    .X(_00070_));
 sg13g2_mux2_1 _11698_ (.A0(net1814),
    .A1(net5107),
    .S(_04033_),
    .X(_00071_));
 sg13g2_mux2_1 _11699_ (.A0(net1798),
    .A1(net4880),
    .S(_04033_),
    .X(_00072_));
 sg13g2_mux2_1 _11700_ (.A0(net1797),
    .A1(net5010),
    .S(_04033_),
    .X(_00073_));
 sg13g2_nor2_1 _11701_ (.A(net2606),
    .B(_01980_),
    .Y(_04034_));
 sg13g2_nor4_1 _11702_ (.A(net2604),
    .B(net2606),
    .C(_01980_),
    .D(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .Y(_04035_));
 sg13g2_nand2_1 _11703_ (.Y(_04036_),
    .A(net2439),
    .B(_04035_));
 sg13g2_and2_1 _11704_ (.A(net2604),
    .B(_04034_),
    .X(_04037_));
 sg13g2_nor2b_1 _11705_ (.A(net2604),
    .B_N(net2606),
    .Y(_04038_));
 sg13g2_nand2b_2 _11706_ (.Y(_04039_),
    .B(net2606),
    .A_N(net2604));
 sg13g2_nor2_2 _11707_ (.A(net2607),
    .B(_04039_),
    .Y(_04040_));
 sg13g2_nand2_1 _11708_ (.Y(_04041_),
    .A(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .B(_04040_));
 sg13g2_o21ai_1 _11709_ (.B1(_04037_),
    .Y(_04042_),
    .A1(net2439),
    .A2(net2596));
 sg13g2_nand3_1 _11710_ (.B(_04041_),
    .C(_04042_),
    .A(_04036_),
    .Y(uio_out[1]));
 sg13g2_nor2_1 _11711_ (.A(_04034_),
    .B(_04040_),
    .Y(_04043_));
 sg13g2_o21ai_1 _11712_ (.B1(_04037_),
    .Y(_04044_),
    .A1(net2439),
    .A2(net2594));
 sg13g2_a21oi_1 _11713_ (.A1(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .A2(_04040_),
    .Y(_04045_),
    .B1(_04043_));
 sg13g2_nand3b_1 _11714_ (.B(_04044_),
    .C(_04045_),
    .Y(uio_out[2]),
    .A_N(_04035_));
 sg13g2_nand2b_1 _11715_ (.Y(_04046_),
    .B(net2609),
    .A_N(net2592));
 sg13g2_a22oi_1 _11716_ (.Y(_04047_),
    .B1(_04046_),
    .B2(_04037_),
    .A2(_04040_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[22] ));
 sg13g2_inv_2 _11717_ (.Y(uio_out[4]),
    .A(_04047_));
 sg13g2_o21ai_1 _11718_ (.B1(_04037_),
    .Y(_04048_),
    .A1(net2439),
    .A2(net2590));
 sg13g2_a21oi_1 _11719_ (.A1(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .A2(_04040_),
    .Y(_04049_),
    .B1(_04043_));
 sg13g2_nand3_1 _11720_ (.B(_04048_),
    .C(_04049_),
    .A(_04036_),
    .Y(uio_out[5]));
 sg13g2_and2_1 _11721_ (.A(\i_latch_mem.genblk1[5].l_ram.data_out[0] ),
    .B(net2098),
    .X(_04050_));
 sg13g2_a22oi_1 _11722_ (.Y(_04051_),
    .B1(net2012),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[0] ),
    .A2(net2032),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11723_ (.Y(_04052_),
    .B1(net2011),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[0] ),
    .A2(net2031),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11724_ (.Y(_04053_),
    .B1(_02430_),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[0] ),
    .A2(net2090),
    .A1(\i_latch_mem.genblk1[23].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11725_ (.Y(_04054_),
    .B1(net2029),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[0] ),
    .A2(net2097),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11726_ (.Y(_04055_),
    .B1(_02370_),
    .B2(\i_latch_mem.genblk1[22].l_ram.data_out[0] ),
    .A2(net2094),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[0] ));
 sg13g2_nand3_1 _11727_ (.B(_04054_),
    .C(_04055_),
    .A(_04053_),
    .Y(_04056_));
 sg13g2_a221oi_1 _11728_ (.B2(\i_latch_mem.genblk1[30].l_ram.data_out[0] ),
    .C1(_04056_),
    .B1(net2008),
    .A1(\i_latch_mem.genblk1[21].l_ram.data_out[0] ),
    .Y(_04057_),
    .A2(net2092));
 sg13g2_a221oi_1 _11729_ (.B2(\i_latch_mem.genblk1[13].l_ram.data_out[0] ),
    .C1(_04050_),
    .B1(net2095),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[0] ),
    .Y(_04058_),
    .A2(net2099));
 sg13g2_a22oi_1 _11730_ (.Y(_04059_),
    .B1(net2093),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[0] ),
    .A2(_02288_),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11731_ (.Y(_04060_),
    .B1(net2100),
    .B2(\i_latch_mem.genblk1[31].l_ram.data_out[0] ),
    .A2(net2101),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[0] ));
 sg13g2_nand4_1 _11732_ (.B(_04058_),
    .C(_04059_),
    .A(_04057_),
    .Y(_04061_),
    .D(_04060_));
 sg13g2_a22oi_1 _11733_ (.Y(_04062_),
    .B1(net2022),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[0] ),
    .A2(net1993),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11734_ (.Y(_04063_),
    .B1(net1963),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[0] ),
    .A2(net2013),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11735_ (.Y(_04064_),
    .B1(net1977),
    .B2(\i_latch_mem.genblk1[18].l_ram.data_out[0] ),
    .A2(net1992),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[0] ));
 sg13g2_a22oi_1 _11736_ (.Y(_04065_),
    .B1(net2023),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[0] ),
    .A2(net1980),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[0] ));
 sg13g2_nand4_1 _11737_ (.B(_04063_),
    .C(_04064_),
    .A(_04062_),
    .Y(_04066_),
    .D(_04065_));
 sg13g2_a221oi_1 _11738_ (.B2(\i_latch_mem.genblk1[11].l_ram.data_out[0] ),
    .C1(_02235_),
    .B1(net2030),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[0] ),
    .Y(_04067_),
    .A2(net2096));
 sg13g2_a22oi_1 _11739_ (.Y(_04068_),
    .B1(net2007),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[0] ),
    .A2(net2010),
    .A1(\i_latch_mem.genblk1[27].l_ram.data_out[0] ));
 sg13g2_nand4_1 _11740_ (.B(_04052_),
    .C(_04067_),
    .A(_04051_),
    .Y(_04069_),
    .D(_04068_));
 sg13g2_or3_1 _11741_ (.A(_04061_),
    .B(_04066_),
    .C(_04069_),
    .X(_04070_));
 sg13g2_o21ai_1 _11742_ (.B1(_04070_),
    .Y(_04071_),
    .A1(\i_latch_mem.genblk1[0].l_ram.data_out[0] ),
    .A2(_02236_));
 sg13g2_nor2_1 _11743_ (.A(net3920),
    .B(net2392),
    .Y(_04072_));
 sg13g2_a21oi_1 _11744_ (.A1(net2392),
    .A2(_04071_),
    .Y(_00012_),
    .B1(_04072_));
 sg13g2_and2_1 _11745_ (.A(\i_latch_mem.genblk1[6].l_ram.data_out[1] ),
    .B(net2097),
    .X(_04073_));
 sg13g2_a22oi_1 _11746_ (.Y(_04074_),
    .B1(net1992),
    .B2(\i_latch_mem.genblk1[3].l_ram.data_out[1] ),
    .A2(net1993),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11747_ (.Y(_04075_),
    .B1(net2099),
    .B2(\i_latch_mem.genblk1[4].l_ram.data_out[1] ),
    .A2(net2100),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11748_ (.Y(_04076_),
    .B1(net2095),
    .B2(\i_latch_mem.genblk1[13].l_ram.data_out[1] ),
    .A2(_02192_),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11749_ (.Y(_04077_),
    .B1(net2093),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[1] ),
    .A2(net2094),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[1] ));
 sg13g2_nand3_1 _11750_ (.B(_04076_),
    .C(_04077_),
    .A(_04075_),
    .Y(_04078_));
 sg13g2_a221oi_1 _11751_ (.B2(\i_latch_mem.genblk1[28].l_ram.data_out[1] ),
    .C1(_04078_),
    .B1(net2009),
    .A1(\i_latch_mem.genblk1[12].l_ram.data_out[1] ),
    .Y(_04079_),
    .A2(net2029));
 sg13g2_a221oi_1 _11752_ (.B2(\i_latch_mem.genblk1[30].l_ram.data_out[1] ),
    .C1(_04073_),
    .B1(net2008),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[1] ),
    .Y(_04080_),
    .A2(net2096));
 sg13g2_a22oi_1 _11753_ (.Y(_04081_),
    .B1(net2092),
    .B2(\i_latch_mem.genblk1[21].l_ram.data_out[1] ),
    .A2(net2026),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11754_ (.Y(_04082_),
    .B1(net2090),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[1] ),
    .A2(net2091),
    .A1(\i_latch_mem.genblk1[22].l_ram.data_out[1] ));
 sg13g2_nand4_1 _11755_ (.B(_04080_),
    .C(_04081_),
    .A(_04079_),
    .Y(_04083_),
    .D(_04082_));
 sg13g2_a22oi_1 _11756_ (.Y(_04084_),
    .B1(net2013),
    .B2(\i_latch_mem.genblk1[24].l_ram.data_out[1] ),
    .A2(net2022),
    .A1(\i_latch_mem.genblk1[1].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11757_ (.Y(_04085_),
    .B1(_02330_),
    .B2(\i_latch_mem.genblk1[18].l_ram.data_out[1] ),
    .A2(net1980),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11758_ (.Y(_04086_),
    .B1(net2007),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[1] ),
    .A2(net2030),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11759_ (.Y(_04087_),
    .B1(net2023),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[1] ),
    .A2(net2032),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[1] ));
 sg13g2_nand4_1 _11760_ (.B(_04085_),
    .C(_04086_),
    .A(_04084_),
    .Y(_04088_),
    .D(_04087_));
 sg13g2_a221oi_1 _11761_ (.B2(\i_latch_mem.genblk1[10].l_ram.data_out[1] ),
    .C1(net1989),
    .B1(_02246_),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[1] ),
    .Y(_04089_),
    .A2(net2101));
 sg13g2_a22oi_1 _11762_ (.Y(_04090_),
    .B1(net1963),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[1] ),
    .A2(net2012),
    .A1(\i_latch_mem.genblk1[25].l_ram.data_out[1] ));
 sg13g2_a22oi_1 _11763_ (.Y(_04091_),
    .B1(net2010),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[1] ),
    .A2(net2011),
    .A1(\i_latch_mem.genblk1[26].l_ram.data_out[1] ));
 sg13g2_nand4_1 _11764_ (.B(_04089_),
    .C(_04090_),
    .A(_04074_),
    .Y(_04092_),
    .D(_04091_));
 sg13g2_or3_1 _11765_ (.A(_04083_),
    .B(_04088_),
    .C(_04092_),
    .X(_04093_));
 sg13g2_o21ai_1 _11766_ (.B1(_04093_),
    .Y(_04094_),
    .A1(\i_latch_mem.genblk1[0].l_ram.data_out[1] ),
    .A2(_02236_));
 sg13g2_nor2_1 _11767_ (.A(net3734),
    .B(net2391),
    .Y(_04095_));
 sg13g2_a21oi_1 _11768_ (.A1(net2391),
    .A2(_04094_),
    .Y(_00023_),
    .B1(_04095_));
 sg13g2_and2_1 _11769_ (.A(\i_latch_mem.genblk1[13].l_ram.data_out[2] ),
    .B(net2095),
    .X(_04096_));
 sg13g2_a22oi_1 _11770_ (.Y(_04097_),
    .B1(net2008),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[2] ),
    .A2(net2101),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11771_ (.Y(_04098_),
    .B1(net2092),
    .B2(\i_latch_mem.genblk1[21].l_ram.data_out[2] ),
    .A2(net2026),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11772_ (.Y(_04099_),
    .B1(net2090),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[2] ),
    .A2(net2093),
    .A1(\i_latch_mem.genblk1[20].l_ram.data_out[2] ));
 sg13g2_nand3_1 _11773_ (.B(_04098_),
    .C(_04099_),
    .A(_04097_),
    .Y(_04100_));
 sg13g2_a221oi_1 _11774_ (.B2(\i_latch_mem.genblk1[22].l_ram.data_out[2] ),
    .C1(_04100_),
    .B1(net2091),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[2] ),
    .Y(_04101_),
    .A2(net2096));
 sg13g2_a221oi_1 _11775_ (.B2(\i_latch_mem.genblk1[28].l_ram.data_out[2] ),
    .C1(_04096_),
    .B1(net2009),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[2] ),
    .Y(_04102_),
    .A2(_02158_));
 sg13g2_a22oi_1 _11776_ (.Y(_04103_),
    .B1(net2029),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[2] ),
    .A2(net2099),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11777_ (.Y(_04104_),
    .B1(net2097),
    .B2(\i_latch_mem.genblk1[6].l_ram.data_out[2] ),
    .A2(net2098),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[2] ));
 sg13g2_nand4_1 _11778_ (.B(_04102_),
    .C(_04103_),
    .A(_04101_),
    .Y(_04105_),
    .D(_04104_));
 sg13g2_a22oi_1 _11779_ (.Y(_04106_),
    .B1(net1992),
    .B2(\i_latch_mem.genblk1[3].l_ram.data_out[2] ),
    .A2(net1993),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11780_ (.Y(_04107_),
    .B1(net2030),
    .B2(\i_latch_mem.genblk1[11].l_ram.data_out[2] ),
    .A2(net2031),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11781_ (.Y(_04108_),
    .B1(net1963),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[2] ),
    .A2(net1977),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11782_ (.Y(_04109_),
    .B1(net2007),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[2] ),
    .A2(net1980),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[2] ));
 sg13g2_nand4_1 _11783_ (.B(_04107_),
    .C(_04108_),
    .A(_04106_),
    .Y(_04110_),
    .D(_04109_));
 sg13g2_a221oi_1 _11784_ (.B2(\i_latch_mem.genblk1[1].l_ram.data_out[2] ),
    .C1(net1989),
    .B1(net2022),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[2] ),
    .Y(_04111_),
    .A2(net2094));
 sg13g2_a22oi_1 _11785_ (.Y(_04112_),
    .B1(net2013),
    .B2(\i_latch_mem.genblk1[24].l_ram.data_out[2] ),
    .A2(net2023),
    .A1(\i_latch_mem.genblk1[17].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11786_ (.Y(_04113_),
    .B1(net2011),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[2] ),
    .A2(net2012),
    .A1(\i_latch_mem.genblk1[25].l_ram.data_out[2] ));
 sg13g2_a22oi_1 _11787_ (.Y(_04114_),
    .B1(net2010),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[2] ),
    .A2(net2032),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[2] ));
 sg13g2_nand4_1 _11788_ (.B(_04112_),
    .C(_04113_),
    .A(_04111_),
    .Y(_04115_),
    .D(_04114_));
 sg13g2_or3_1 _11789_ (.A(_04105_),
    .B(_04110_),
    .C(_04115_),
    .X(_04116_));
 sg13g2_o21ai_1 _11790_ (.B1(_04116_),
    .Y(_04117_),
    .A1(\i_latch_mem.genblk1[0].l_ram.data_out[2] ),
    .A2(_02236_));
 sg13g2_nor2_1 _11791_ (.A(net3806),
    .B(net2392),
    .Y(_04118_));
 sg13g2_a21oi_1 _11792_ (.A1(net2392),
    .A2(_04117_),
    .Y(_00034_),
    .B1(_04118_));
 sg13g2_nor2_1 _11793_ (.A(net3894),
    .B(net2391),
    .Y(_04119_));
 sg13g2_nand2_1 _11794_ (.Y(_04120_),
    .A(\i_latch_mem.genblk1[30].l_ram.data_out[3] ),
    .B(net2008));
 sg13g2_a22oi_1 _11795_ (.Y(_04121_),
    .B1(net2011),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[3] ),
    .A2(net1992),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11796_ (.Y(_04122_),
    .B1(net1977),
    .B2(\i_latch_mem.genblk1[18].l_ram.data_out[3] ),
    .A2(net2030),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11797_ (.Y(_04123_),
    .B1(_02360_),
    .B2(\i_latch_mem.genblk1[21].l_ram.data_out[3] ),
    .A2(net2026),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11798_ (.Y(_04124_),
    .B1(_02350_),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[3] ),
    .A2(_02213_),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11799_ (.Y(_04125_),
    .B1(_02298_),
    .B2(\i_latch_mem.genblk1[15].l_ram.data_out[3] ),
    .A2(_02148_),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11800_ (.Y(_04126_),
    .B1(net2090),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[3] ),
    .A2(net2097),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[3] ));
 sg13g2_nand4_1 _11801_ (.B(_04124_),
    .C(_04125_),
    .A(_04123_),
    .Y(_04127_),
    .D(_04126_));
 sg13g2_a22oi_1 _11802_ (.Y(_04128_),
    .B1(net2029),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[3] ),
    .A2(net2098),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11803_ (.Y(_04129_),
    .B1(net2095),
    .B2(\i_latch_mem.genblk1[13].l_ram.data_out[3] ),
    .A2(net2100),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11804_ (.Y(_04130_),
    .B1(net2009),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[3] ),
    .A2(net2091),
    .A1(\i_latch_mem.genblk1[22].l_ram.data_out[3] ));
 sg13g2_nand4_1 _11805_ (.B(_04128_),
    .C(_04129_),
    .A(_04120_),
    .Y(_04131_),
    .D(_04130_));
 sg13g2_nor2_1 _11806_ (.A(_04127_),
    .B(_04131_),
    .Y(_04132_));
 sg13g2_a22oi_1 _11807_ (.Y(_04133_),
    .B1(net2031),
    .B2(\i_latch_mem.genblk1[10].l_ram.data_out[3] ),
    .A2(_02182_),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11808_ (.Y(_04134_),
    .B1(net2010),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[3] ),
    .A2(net2032),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[3] ));
 sg13g2_a22oi_1 _11809_ (.Y(_04135_),
    .B1(net2022),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[3] ),
    .A2(net2023),
    .A1(\i_latch_mem.genblk1[17].l_ram.data_out[3] ));
 sg13g2_nand4_1 _11810_ (.B(_04133_),
    .C(_04134_),
    .A(_02236_),
    .Y(_04136_),
    .D(_04135_));
 sg13g2_a221oi_1 _11811_ (.B2(\i_latch_mem.genblk1[9].l_ram.data_out[3] ),
    .C1(_04136_),
    .B1(net2007),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[3] ),
    .Y(_04137_),
    .A2(net2013));
 sg13g2_a22oi_1 _11812_ (.Y(_04138_),
    .B1(net2012),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[3] ),
    .A2(net1980),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[3] ));
 sg13g2_nand3_1 _11813_ (.B(_04122_),
    .C(_04138_),
    .A(_04121_),
    .Y(_04139_));
 sg13g2_a221oi_1 _11814_ (.B2(\i_latch_mem.genblk1[2].l_ram.data_out[3] ),
    .C1(_04139_),
    .B1(net1963),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[3] ),
    .Y(_04140_),
    .A2(_02107_));
 sg13g2_nand3_1 _11815_ (.B(_04137_),
    .C(_04140_),
    .A(_04132_),
    .Y(_04141_));
 sg13g2_o21ai_1 _11816_ (.B1(_04141_),
    .Y(_04142_),
    .A1(\i_latch_mem.genblk1[0].l_ram.data_out[3] ),
    .A2(_02236_));
 sg13g2_a21oi_1 _11817_ (.A1(net2391),
    .A2(_04142_),
    .Y(_00037_),
    .B1(_04119_));
 sg13g2_a22oi_1 _11818_ (.Y(_04143_),
    .B1(net2091),
    .B2(\i_latch_mem.genblk1[22].l_ram.data_out[4] ),
    .A2(net2026),
    .A1(\i_latch_mem.genblk1[14].l_ram.data_out[4] ));
 sg13g2_nand2_1 _11819_ (.Y(_04144_),
    .A(\i_latch_mem.genblk1[13].l_ram.data_out[4] ),
    .B(net2095));
 sg13g2_a22oi_1 _11820_ (.Y(_04145_),
    .B1(net2010),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[4] ),
    .A2(net1980),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11821_ (.Y(_04146_),
    .B1(net2022),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[4] ),
    .A2(net1992),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11822_ (.Y(_04147_),
    .B1(net2023),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[4] ),
    .A2(net1993),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11823_ (.Y(_04148_),
    .B1(_02410_),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[4] ),
    .A2(net2012),
    .A1(\i_latch_mem.genblk1[25].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11824_ (.Y(_04149_),
    .B1(net2031),
    .B2(\i_latch_mem.genblk1[10].l_ram.data_out[4] ),
    .A2(net2032),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11825_ (.Y(_04150_),
    .B1(_02267_),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[4] ),
    .A2(net2100),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11826_ (.Y(_04151_),
    .B1(net2090),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[4] ),
    .A2(net2096),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11827_ (.Y(_04152_),
    .B1(net2094),
    .B2(\i_latch_mem.genblk1[15].l_ram.data_out[4] ),
    .A2(net2098),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[4] ));
 sg13g2_nand4_1 _11828_ (.B(_04150_),
    .C(_04151_),
    .A(_04143_),
    .Y(_04153_),
    .D(_04152_));
 sg13g2_a22oi_1 _11829_ (.Y(_04154_),
    .B1(net2009),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[4] ),
    .A2(net2092),
    .A1(\i_latch_mem.genblk1[21].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11830_ (.Y(_04155_),
    .B1(net2097),
    .B2(\i_latch_mem.genblk1[6].l_ram.data_out[4] ),
    .A2(net2099),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[4] ));
 sg13g2_a22oi_1 _11831_ (.Y(_04156_),
    .B1(net2008),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[4] ),
    .A2(net2101),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[4] ));
 sg13g2_nand4_1 _11832_ (.B(_04154_),
    .C(_04155_),
    .A(_04144_),
    .Y(_04157_),
    .D(_04156_));
 sg13g2_nor2_1 _11833_ (.A(_04153_),
    .B(_04157_),
    .Y(_04158_));
 sg13g2_a22oi_1 _11834_ (.Y(_04159_),
    .B1(net2013),
    .B2(\i_latch_mem.genblk1[24].l_ram.data_out[4] ),
    .A2(net2030),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[4] ));
 sg13g2_a221oi_1 _11835_ (.B2(\i_latch_mem.genblk1[9].l_ram.data_out[4] ),
    .C1(net1989),
    .B1(net2007),
    .A1(\i_latch_mem.genblk1[20].l_ram.data_out[4] ),
    .Y(_04160_),
    .A2(net2093));
 sg13g2_nand4_1 _11836_ (.B(_04149_),
    .C(_04159_),
    .A(_04148_),
    .Y(_04161_),
    .D(_04160_));
 sg13g2_a22oi_1 _11837_ (.Y(_04162_),
    .B1(net1963),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[4] ),
    .A2(net1977),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[4] ));
 sg13g2_nand4_1 _11838_ (.B(_04146_),
    .C(_04147_),
    .A(_04145_),
    .Y(_04163_),
    .D(_04162_));
 sg13g2_nor2_1 _11839_ (.A(_04161_),
    .B(_04163_),
    .Y(_04164_));
 sg13g2_a22oi_1 _11840_ (.Y(_04165_),
    .B1(_04158_),
    .B2(_04164_),
    .A2(net1989),
    .A1(_01745_));
 sg13g2_nand2_1 _11841_ (.Y(_04166_),
    .A(net2393),
    .B(_04165_));
 sg13g2_o21ai_1 _11842_ (.B1(_04166_),
    .Y(_00038_),
    .A1(_02062_),
    .A2(net2393));
 sg13g2_nand2_1 _11843_ (.Y(_04167_),
    .A(\i_latch_mem.genblk1[14].l_ram.data_out[5] ),
    .B(net2026));
 sg13g2_a22oi_1 _11844_ (.Y(_04168_),
    .B1(net2091),
    .B2(\i_latch_mem.genblk1[22].l_ram.data_out[5] ),
    .A2(net2100),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11845_ (.Y(_04169_),
    .B1(net2012),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[5] ),
    .A2(net1993),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11846_ (.Y(_04170_),
    .B1(net2011),
    .B2(\i_latch_mem.genblk1[26].l_ram.data_out[5] ),
    .A2(net1977),
    .A1(\i_latch_mem.genblk1[18].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11847_ (.Y(_04171_),
    .B1(net2023),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[5] ),
    .A2(net1980),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11848_ (.Y(_04172_),
    .B1(net2010),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[5] ),
    .A2(net2013),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11849_ (.Y(_04173_),
    .B1(net2029),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[5] ),
    .A2(net2096),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11850_ (.Y(_04174_),
    .B1(net2093),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[5] ),
    .A2(net2094),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11851_ (.Y(_04175_),
    .B1(net2008),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[5] ),
    .A2(net2101),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[5] ));
 sg13g2_nand4_1 _11852_ (.B(_04173_),
    .C(_04174_),
    .A(_04168_),
    .Y(_04176_),
    .D(_04175_));
 sg13g2_a22oi_1 _11853_ (.Y(_04177_),
    .B1(net2009),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[5] ),
    .A2(net2095),
    .A1(\i_latch_mem.genblk1[13].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11854_ (.Y(_04178_),
    .B1(net2090),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[5] ),
    .A2(net2092),
    .A1(\i_latch_mem.genblk1[21].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11855_ (.Y(_04179_),
    .B1(net2098),
    .B2(\i_latch_mem.genblk1[5].l_ram.data_out[5] ),
    .A2(net2099),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[5] ));
 sg13g2_nand4_1 _11856_ (.B(_04177_),
    .C(_04178_),
    .A(_04167_),
    .Y(_04180_),
    .D(_04179_));
 sg13g2_nor2_1 _11857_ (.A(_04176_),
    .B(_04180_),
    .Y(_04181_));
 sg13g2_a22oi_1 _11858_ (.Y(_04182_),
    .B1(net2030),
    .B2(\i_latch_mem.genblk1[11].l_ram.data_out[5] ),
    .A2(net2031),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[5] ));
 sg13g2_a221oi_1 _11859_ (.B2(\i_latch_mem.genblk1[9].l_ram.data_out[5] ),
    .C1(net1989),
    .B1(net2007),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[5] ),
    .Y(_04183_),
    .A2(net2097));
 sg13g2_nand4_1 _11860_ (.B(_04171_),
    .C(_04182_),
    .A(_04170_),
    .Y(_04184_),
    .D(_04183_));
 sg13g2_a22oi_1 _11861_ (.Y(_04185_),
    .B1(net1963),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[5] ),
    .A2(net2032),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[5] ));
 sg13g2_a22oi_1 _11862_ (.Y(_04186_),
    .B1(net2022),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[5] ),
    .A2(net1992),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[5] ));
 sg13g2_nand4_1 _11863_ (.B(_04172_),
    .C(_04185_),
    .A(_04169_),
    .Y(_04187_),
    .D(_04186_));
 sg13g2_nor2_1 _11864_ (.A(_04184_),
    .B(_04187_),
    .Y(_04188_));
 sg13g2_a22oi_1 _11865_ (.Y(_04189_),
    .B1(_04181_),
    .B2(_04188_),
    .A2(net1989),
    .A1(_01744_));
 sg13g2_nand2_1 _11866_ (.Y(_04190_),
    .A(net2391),
    .B(_04189_));
 sg13g2_o21ai_1 _11867_ (.B1(_04190_),
    .Y(_00039_),
    .A1(_02070_),
    .A2(net2391));
 sg13g2_nand2_1 _11868_ (.Y(_04191_),
    .A(\i_latch_mem.genblk1[7].l_ram.data_out[6] ),
    .B(net2096));
 sg13g2_a22oi_1 _11869_ (.Y(_04192_),
    .B1(net1963),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[6] ),
    .A2(net2022),
    .A1(\i_latch_mem.genblk1[1].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11870_ (.Y(_04193_),
    .B1(net2023),
    .B2(\i_latch_mem.genblk1[17].l_ram.data_out[6] ),
    .A2(net1993),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11871_ (.Y(_04194_),
    .B1(net2007),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[6] ),
    .A2(net2011),
    .A1(\i_latch_mem.genblk1[26].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11872_ (.Y(_04195_),
    .B1(_02400_),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[6] ),
    .A2(net2013),
    .A1(\i_latch_mem.genblk1[24].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11873_ (.Y(_04196_),
    .B1(net2029),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[6] ),
    .A2(net2097),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11874_ (.Y(_04197_),
    .B1(_02380_),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[6] ),
    .A2(net2101),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11875_ (.Y(_04198_),
    .B1(net2009),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[6] ),
    .A2(net2099),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11876_ (.Y(_04199_),
    .B1(net2008),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[6] ),
    .A2(net2100),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[6] ));
 sg13g2_nand4_1 _11877_ (.B(_04197_),
    .C(_04198_),
    .A(_04196_),
    .Y(_04200_),
    .D(_04199_));
 sg13g2_a22oi_1 _11878_ (.Y(_04201_),
    .B1(net2093),
    .B2(\i_latch_mem.genblk1[20].l_ram.data_out[6] ),
    .A2(_02277_),
    .A1(\i_latch_mem.genblk1[13].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11879_ (.Y(_04202_),
    .B1(net2091),
    .B2(\i_latch_mem.genblk1[22].l_ram.data_out[6] ),
    .A2(net2094),
    .A1(\i_latch_mem.genblk1[15].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11880_ (.Y(_04203_),
    .B1(net2026),
    .B2(\i_latch_mem.genblk1[14].l_ram.data_out[6] ),
    .A2(net2098),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[6] ));
 sg13g2_nand4_1 _11881_ (.B(_04201_),
    .C(_04202_),
    .A(_04191_),
    .Y(_04204_),
    .D(_04203_));
 sg13g2_nor2_1 _11882_ (.A(_04200_),
    .B(_04204_),
    .Y(_04205_));
 sg13g2_a22oi_1 _11883_ (.Y(_04206_),
    .B1(net1977),
    .B2(\i_latch_mem.genblk1[18].l_ram.data_out[6] ),
    .A2(net2031),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[6] ));
 sg13g2_a22oi_1 _11884_ (.Y(_04207_),
    .B1(_02420_),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[6] ),
    .A2(net2030),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[6] ));
 sg13g2_nand4_1 _11885_ (.B(_04193_),
    .C(_04206_),
    .A(_04192_),
    .Y(_04208_),
    .D(_04207_));
 sg13g2_a22oi_1 _11886_ (.Y(_04209_),
    .B1(net1980),
    .B2(\i_latch_mem.genblk1[16].l_ram.data_out[6] ),
    .A2(net1992),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[6] ));
 sg13g2_a221oi_1 _11887_ (.B2(\i_latch_mem.genblk1[21].l_ram.data_out[6] ),
    .C1(_02235_),
    .B1(net2092),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[6] ),
    .Y(_04210_),
    .A2(_02224_));
 sg13g2_nand4_1 _11888_ (.B(_04195_),
    .C(_04209_),
    .A(_04194_),
    .Y(_04211_),
    .D(_04210_));
 sg13g2_nor2_1 _11889_ (.A(_04208_),
    .B(_04211_),
    .Y(_04212_));
 sg13g2_a22oi_1 _11890_ (.Y(_04213_),
    .B1(_04205_),
    .B2(_04212_),
    .A2(net1989),
    .A1(_01743_));
 sg13g2_nand2_1 _11891_ (.Y(_04214_),
    .A(net2391),
    .B(_04213_));
 sg13g2_o21ai_1 _11892_ (.B1(_04214_),
    .Y(_00040_),
    .A1(_02076_),
    .A2(net2391));
 sg13g2_nor2_1 _11893_ (.A(net3787),
    .B(net2393),
    .Y(_04215_));
 sg13g2_and2_1 _11894_ (.A(\i_latch_mem.genblk1[22].l_ram.data_out[7] ),
    .B(net2091),
    .X(_04216_));
 sg13g2_a22oi_1 _11895_ (.Y(_04217_),
    .B1(_02340_),
    .B2(\i_latch_mem.genblk1[1].l_ram.data_out[7] ),
    .A2(_02168_),
    .A1(\i_latch_mem.genblk1[3].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11896_ (.Y(_04218_),
    .B1(net2009),
    .B2(\i_latch_mem.genblk1[28].l_ram.data_out[7] ),
    .A2(net2092),
    .A1(\i_latch_mem.genblk1[21].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11897_ (.Y(_04219_),
    .B1(net2094),
    .B2(\i_latch_mem.genblk1[15].l_ram.data_out[7] ),
    .A2(_02203_),
    .A1(\i_latch_mem.genblk1[6].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11898_ (.Y(_04220_),
    .B1(net2029),
    .B2(\i_latch_mem.genblk1[12].l_ram.data_out[7] ),
    .A2(net2099),
    .A1(\i_latch_mem.genblk1[4].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11899_ (.Y(_04221_),
    .B1(_02450_),
    .B2(\i_latch_mem.genblk1[30].l_ram.data_out[7] ),
    .A2(net2100),
    .A1(\i_latch_mem.genblk1[31].l_ram.data_out[7] ));
 sg13g2_nand3_1 _11900_ (.B(_04220_),
    .C(_04221_),
    .A(_04219_),
    .Y(_04222_));
 sg13g2_a221oi_1 _11901_ (.B2(\i_latch_mem.genblk1[14].l_ram.data_out[7] ),
    .C1(_04222_),
    .B1(net2026),
    .A1(\i_latch_mem.genblk1[7].l_ram.data_out[7] ),
    .Y(_04223_),
    .A2(net2096));
 sg13g2_a221oi_1 _11902_ (.B2(\i_latch_mem.genblk1[13].l_ram.data_out[7] ),
    .C1(_04216_),
    .B1(net2095),
    .A1(\i_latch_mem.genblk1[29].l_ram.data_out[7] ),
    .Y(_04224_),
    .A2(net2101));
 sg13g2_a22oi_1 _11903_ (.Y(_04225_),
    .B1(net2090),
    .B2(\i_latch_mem.genblk1[23].l_ram.data_out[7] ),
    .A2(net2098),
    .A1(\i_latch_mem.genblk1[5].l_ram.data_out[7] ));
 sg13g2_nand4_1 _11904_ (.B(_04223_),
    .C(_04224_),
    .A(_04218_),
    .Y(_04226_),
    .D(_04225_));
 sg13g2_a22oi_1 _11905_ (.Y(_04227_),
    .B1(net1977),
    .B2(\i_latch_mem.genblk1[18].l_ram.data_out[7] ),
    .A2(net1993),
    .A1(\i_latch_mem.genblk1[19].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11906_ (.Y(_04228_),
    .B1(_02460_),
    .B2(\i_latch_mem.genblk1[9].l_ram.data_out[7] ),
    .A2(net1980),
    .A1(\i_latch_mem.genblk1[16].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11907_ (.Y(_04229_),
    .B1(net2010),
    .B2(\i_latch_mem.genblk1[27].l_ram.data_out[7] ),
    .A2(net2011),
    .A1(\i_latch_mem.genblk1[26].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11908_ (.Y(_04230_),
    .B1(net2013),
    .B2(\i_latch_mem.genblk1[24].l_ram.data_out[7] ),
    .A2(_02319_),
    .A1(\i_latch_mem.genblk1[17].l_ram.data_out[7] ));
 sg13g2_nand4_1 _11909_ (.B(_04228_),
    .C(_04229_),
    .A(_04227_),
    .Y(_04231_),
    .D(_04230_));
 sg13g2_a221oi_1 _11910_ (.B2(\i_latch_mem.genblk1[20].l_ram.data_out[7] ),
    .C1(_02235_),
    .B1(net2093),
    .A1(\i_latch_mem.genblk1[11].l_ram.data_out[7] ),
    .Y(_04232_),
    .A2(_02256_));
 sg13g2_a22oi_1 _11911_ (.Y(_04233_),
    .B1(net1963),
    .B2(\i_latch_mem.genblk1[2].l_ram.data_out[7] ),
    .A2(net2031),
    .A1(\i_latch_mem.genblk1[10].l_ram.data_out[7] ));
 sg13g2_a22oi_1 _11912_ (.Y(_04234_),
    .B1(net2012),
    .B2(\i_latch_mem.genblk1[25].l_ram.data_out[7] ),
    .A2(net2032),
    .A1(\i_latch_mem.genblk1[8].l_ram.data_out[7] ));
 sg13g2_nand4_1 _11913_ (.B(_04232_),
    .C(_04233_),
    .A(_04217_),
    .Y(_04235_),
    .D(_04234_));
 sg13g2_or3_1 _11914_ (.A(_04226_),
    .B(_04231_),
    .C(_04235_),
    .X(_04236_));
 sg13g2_o21ai_1 _11915_ (.B1(_04236_),
    .Y(_04237_),
    .A1(\i_latch_mem.genblk1[0].l_ram.data_out[7] ),
    .A2(_02236_));
 sg13g2_a21oi_1 _11916_ (.A1(net2393),
    .A2(_04237_),
    .Y(_00041_),
    .B1(_04215_));
 sg13g2_nor2_1 _11917_ (.A(net3875),
    .B(net2402),
    .Y(_04238_));
 sg13g2_a21oi_1 _11918_ (.A1(net2402),
    .A2(_04071_),
    .Y(_00042_),
    .B1(_04238_));
 sg13g2_nor2_1 _11919_ (.A(net3761),
    .B(net2402),
    .Y(_04239_));
 sg13g2_a21oi_1 _11920_ (.A1(net2402),
    .A2(_04094_),
    .Y(_00043_),
    .B1(_04239_));
 sg13g2_nor2_1 _11921_ (.A(net3853),
    .B(net2402),
    .Y(_04240_));
 sg13g2_a21oi_1 _11922_ (.A1(net2405),
    .A2(_04117_),
    .Y(_00013_),
    .B1(_04240_));
 sg13g2_nor2_1 _11923_ (.A(net3930),
    .B(net2404),
    .Y(_04241_));
 sg13g2_a21oi_1 _11924_ (.A1(net2403),
    .A2(_04142_),
    .Y(_00014_),
    .B1(_04241_));
 sg13g2_mux2_1 _11925_ (.A0(net4422),
    .A1(_04165_),
    .S(net2403),
    .X(_00015_));
 sg13g2_mux2_1 _11926_ (.A0(net4095),
    .A1(_04189_),
    .S(net2402),
    .X(_00016_));
 sg13g2_mux2_1 _11927_ (.A0(net4063),
    .A1(_04213_),
    .S(net2402),
    .X(_00017_));
 sg13g2_nor2_1 _11928_ (.A(net3703),
    .B(net2404),
    .Y(_04242_));
 sg13g2_a21oi_1 _11929_ (.A1(net2404),
    .A2(_04237_),
    .Y(_00018_),
    .B1(_04242_));
 sg13g2_nor2_1 _11930_ (.A(net3914),
    .B(net2397),
    .Y(_04243_));
 sg13g2_a21oi_1 _11931_ (.A1(_02112_),
    .A2(_04071_),
    .Y(_00019_),
    .B1(_04243_));
 sg13g2_nor2_1 _11932_ (.A(net3757),
    .B(net2396),
    .Y(_04244_));
 sg13g2_a21oi_1 _11933_ (.A1(net2396),
    .A2(_04094_),
    .Y(_00020_),
    .B1(_04244_));
 sg13g2_nor2_1 _11934_ (.A(net3736),
    .B(net2396),
    .Y(_04245_));
 sg13g2_a21oi_1 _11935_ (.A1(net2396),
    .A2(_04117_),
    .Y(_00021_),
    .B1(_04245_));
 sg13g2_nor2_1 _11936_ (.A(net3690),
    .B(net2397),
    .Y(_04246_));
 sg13g2_a21oi_1 _11937_ (.A1(net2397),
    .A2(_04142_),
    .Y(_00022_),
    .B1(_04246_));
 sg13g2_mux2_1 _11938_ (.A0(net4144),
    .A1(_04165_),
    .S(net2397),
    .X(_00024_));
 sg13g2_mux2_1 _11939_ (.A0(net4060),
    .A1(_04189_),
    .S(net2396),
    .X(_00025_));
 sg13g2_mux2_1 _11940_ (.A0(net4121),
    .A1(_04213_),
    .S(net2396),
    .X(_00026_));
 sg13g2_nor2_1 _11941_ (.A(net3816),
    .B(net2396),
    .Y(_04247_));
 sg13g2_a21oi_1 _11942_ (.A1(net2396),
    .A2(_04237_),
    .Y(_00027_),
    .B1(_04247_));
 sg13g2_nand2_1 _11943_ (.Y(_04248_),
    .A(net3490),
    .B(net2399));
 sg13g2_o21ai_1 _11944_ (.B1(_04248_),
    .Y(_00028_),
    .A1(net2399),
    .A2(_04071_));
 sg13g2_nor2_1 _11945_ (.A(net3809),
    .B(net2400),
    .Y(_04249_));
 sg13g2_a21oi_1 _11946_ (.A1(net2400),
    .A2(_04094_),
    .Y(_00029_),
    .B1(_04249_));
 sg13g2_nor2_1 _11947_ (.A(net3834),
    .B(net2400),
    .Y(_04250_));
 sg13g2_a21oi_1 _11948_ (.A1(net2400),
    .A2(_04117_),
    .Y(_00030_),
    .B1(_04250_));
 sg13g2_nor2_1 _11949_ (.A(net3810),
    .B(net2400),
    .Y(_04251_));
 sg13g2_a21oi_1 _11950_ (.A1(net2400),
    .A2(_04142_),
    .Y(_00031_),
    .B1(_04251_));
 sg13g2_nor2_1 _11951_ (.A(net2399),
    .B(_04165_),
    .Y(_04252_));
 sg13g2_a21oi_1 _11952_ (.A1(_02067_),
    .A2(_02111_),
    .Y(_00032_),
    .B1(_04252_));
 sg13g2_nor2_1 _11953_ (.A(net2399),
    .B(_04189_),
    .Y(_04253_));
 sg13g2_a21oi_1 _11954_ (.A1(_02074_),
    .A2(net2399),
    .Y(_00033_),
    .B1(_04253_));
 sg13g2_nor2_1 _11955_ (.A(net2399),
    .B(_04213_),
    .Y(_04254_));
 sg13g2_a21oi_1 _11956_ (.A1(_02080_),
    .A2(net2399),
    .Y(_00035_),
    .B1(_04254_));
 sg13g2_nor2_1 _11957_ (.A(net3764),
    .B(net2400),
    .Y(_04255_));
 sg13g2_a21oi_1 _11958_ (.A1(net2400),
    .A2(_04237_),
    .Y(_00036_),
    .B1(_04255_));
 sg13g2_nor2b_1 _11959_ (.A(_02705_),
    .B_N(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .Y(_04256_));
 sg13g2_nor2_1 _11960_ (.A(net4816),
    .B(net4338),
    .Y(_04257_));
 sg13g2_o21ai_1 _11961_ (.B1(_04257_),
    .Y(_04258_),
    .A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(net2322));
 sg13g2_nor3_1 _11962_ (.A(_03138_),
    .B(_04256_),
    .C(_04258_),
    .Y(_04259_));
 sg13g2_a21oi_1 _11963_ (.A1(net5204),
    .A2(net2318),
    .Y(_04260_),
    .B1(_04259_));
 sg13g2_a21o_1 _11964_ (.A2(_04259_),
    .A1(_03996_),
    .B1(net5205),
    .X(_04261_));
 sg13g2_inv_1 _11965_ (.Y(_00361_),
    .A(_04261_));
 sg13g2_nor3_2 _11966_ (.A(net2325),
    .B(_03436_),
    .C(_03452_),
    .Y(_04262_));
 sg13g2_o21ai_1 _11967_ (.B1(net2632),
    .Y(_04263_),
    .A1(net4934),
    .A2(net2070));
 sg13g2_a21oi_1 _11968_ (.A1(_01779_),
    .A2(net2070),
    .Y(_00362_),
    .B1(_04263_));
 sg13g2_nor2_1 _11969_ (.A(net4834),
    .B(net2070),
    .Y(_04264_));
 sg13g2_and2_1 _11970_ (.A(net2452),
    .B(net2071),
    .X(_04265_));
 sg13g2_nor3_1 _11971_ (.A(net2417),
    .B(_04264_),
    .C(_04265_),
    .Y(_00363_));
 sg13g2_o21ai_1 _11972_ (.B1(net2624),
    .Y(_04266_),
    .A1(net4973),
    .A2(net2071));
 sg13g2_a21oi_1 _11973_ (.A1(_01777_),
    .A2(net2071),
    .Y(_00364_),
    .B1(_04266_));
 sg13g2_o21ai_1 _11974_ (.B1(net2628),
    .Y(_04267_),
    .A1(net4965),
    .A2(net2070));
 sg13g2_a21oi_1 _11975_ (.A1(net2453),
    .A2(net2070),
    .Y(_00365_),
    .B1(_04267_));
 sg13g2_o21ai_1 _11976_ (.B1(net2625),
    .Y(_04268_),
    .A1(net4895),
    .A2(net2071));
 sg13g2_a21oi_1 _11977_ (.A1(_01775_),
    .A2(net2071),
    .Y(_00366_),
    .B1(_04268_));
 sg13g2_o21ai_1 _11978_ (.B1(net2628),
    .Y(_04269_),
    .A1(net4918),
    .A2(net2070));
 sg13g2_a21oi_1 _11979_ (.A1(_01774_),
    .A2(net2070),
    .Y(_00367_),
    .B1(_04269_));
 sg13g2_o21ai_1 _11980_ (.B1(net2626),
    .Y(_04270_),
    .A1(net5049),
    .A2(net2071));
 sg13g2_a21oi_1 _11981_ (.A1(_01773_),
    .A2(net2071),
    .Y(_00368_),
    .B1(_04270_));
 sg13g2_o21ai_1 _11982_ (.B1(net2631),
    .Y(_04271_),
    .A1(net4826),
    .A2(net2070));
 sg13g2_a21oi_1 _11983_ (.A1(_01772_),
    .A2(_04262_),
    .Y(_00369_),
    .B1(_04271_));
 sg13g2_nor4_2 _11984_ (.A(\addr[4] ),
    .B(net2325),
    .C(_03431_),
    .Y(_04272_),
    .D(_03474_));
 sg13g2_o21ai_1 _11985_ (.B1(net2632),
    .Y(_04273_),
    .A1(net4608),
    .A2(net2115));
 sg13g2_a21oi_1 _11986_ (.A1(_01779_),
    .A2(net2115),
    .Y(_00370_),
    .B1(_04273_));
 sg13g2_nor2_1 _11987_ (.A(net3904),
    .B(net2115),
    .Y(_04274_));
 sg13g2_a21oi_1 _11988_ (.A1(_01778_),
    .A2(net2115),
    .Y(_04275_),
    .B1(net2417));
 sg13g2_nor2b_1 _11989_ (.A(_04274_),
    .B_N(_04275_),
    .Y(_00371_));
 sg13g2_o21ai_1 _11990_ (.B1(net2624),
    .Y(_04276_),
    .A1(net4450),
    .A2(net2114));
 sg13g2_a21oi_1 _11991_ (.A1(_01777_),
    .A2(net2114),
    .Y(_00372_),
    .B1(_04276_));
 sg13g2_o21ai_1 _11992_ (.B1(net2628),
    .Y(_04277_),
    .A1(net4636),
    .A2(net2115));
 sg13g2_a21oi_1 _11993_ (.A1(net2453),
    .A2(net2115),
    .Y(_00373_),
    .B1(_04277_));
 sg13g2_o21ai_1 _11994_ (.B1(net2625),
    .Y(_04278_),
    .A1(net4721),
    .A2(net2114));
 sg13g2_a21oi_1 _11995_ (.A1(_01775_),
    .A2(net2114),
    .Y(_00374_),
    .B1(_04278_));
 sg13g2_o21ai_1 _11996_ (.B1(net2626),
    .Y(_04279_),
    .A1(net4456),
    .A2(net2114));
 sg13g2_a21oi_1 _11997_ (.A1(_01774_),
    .A2(net2114),
    .Y(_00375_),
    .B1(_04279_));
 sg13g2_o21ai_1 _11998_ (.B1(net2626),
    .Y(_04280_),
    .A1(net4513),
    .A2(net2114));
 sg13g2_a21oi_1 _11999_ (.A1(_01773_),
    .A2(net2114),
    .Y(_00376_),
    .B1(_04280_));
 sg13g2_o21ai_1 _12000_ (.B1(net2631),
    .Y(_04281_),
    .A1(net4610),
    .A2(net2115));
 sg13g2_a21oi_1 _12001_ (.A1(_01772_),
    .A2(net2115),
    .Y(_00377_),
    .B1(_04281_));
 sg13g2_or3_1 _12002_ (.A(net5152),
    .B(\i_wdt.counter[1] ),
    .C(\i_wdt.counter[0] ),
    .X(_04282_));
 sg13g2_or3_1 _12003_ (.A(net5084),
    .B(\i_wdt.counter[3] ),
    .C(_04282_),
    .X(_04283_));
 sg13g2_nor3_1 _12004_ (.A(net5317),
    .B(net4717),
    .C(_04283_),
    .Y(_04284_));
 sg13g2_nor2b_1 _12005_ (.A(net4395),
    .B_N(_04284_),
    .Y(_04285_));
 sg13g2_nand2b_2 _12006_ (.Y(_04286_),
    .B(_04285_),
    .A_N(net5011));
 sg13g2_or3_1 _12007_ (.A(net5105),
    .B(\i_wdt.counter[9] ),
    .C(_04286_),
    .X(_04287_));
 sg13g2_or2_1 _12008_ (.X(_04288_),
    .B(_04287_),
    .A(net5136));
 sg13g2_nor4_1 _12009_ (.A(net5210),
    .B(net5102),
    .C(\i_wdt.counter[12] ),
    .D(_04288_),
    .Y(_04289_));
 sg13g2_nand2b_1 _12010_ (.Y(_04290_),
    .B(_04289_),
    .A_N(net5384));
 sg13g2_or2_1 _12011_ (.X(_04291_),
    .B(_04290_),
    .A(net5117));
 sg13g2_or3_1 _12012_ (.A(\i_wdt.counter[18] ),
    .B(\i_wdt.counter[17] ),
    .C(_04291_),
    .X(_04292_));
 sg13g2_nor4_1 _12013_ (.A(net5125),
    .B(net5123),
    .C(net4663),
    .D(net5006),
    .Y(_04293_));
 sg13g2_nor2_1 _12014_ (.A(net4869),
    .B(net4432),
    .Y(_04294_));
 sg13g2_nor3_1 _12015_ (.A(net4265),
    .B(net4236),
    .C(net4702),
    .Y(_04295_));
 sg13g2_nand3_1 _12016_ (.B(_04294_),
    .C(_04295_),
    .A(_04293_),
    .Y(_04296_));
 sg13g2_or3_1 _12017_ (.A(net5281),
    .B(_04292_),
    .C(_04296_),
    .X(_04297_));
 sg13g2_nor3_1 _12018_ (.A(net4391),
    .B(net4346),
    .C(net5215),
    .Y(_04298_));
 sg13g2_nor3_1 _12019_ (.A(net4346),
    .B(\i_wdt.counter[29] ),
    .C(_04297_),
    .Y(_04299_));
 sg13g2_nand2b_1 _12020_ (.Y(_04300_),
    .B(_04298_),
    .A_N(_04297_));
 sg13g2_nand2_1 _12021_ (.Y(_04301_),
    .A(net4129),
    .B(net5381));
 sg13g2_nor4_1 _12022_ (.A(net3412),
    .B(net3575),
    .C(net3704),
    .D(_04301_),
    .Y(_04302_));
 sg13g2_nand3_1 _12023_ (.B(_04300_),
    .C(net2302),
    .A(\i_wdt.enabled ),
    .Y(_04303_));
 sg13g2_inv_1 _12024_ (.Y(_04304_),
    .A(_04303_));
 sg13g2_nor4_1 _12025_ (.A(\data_to_write[19] ),
    .B(\data_to_write[18] ),
    .C(\data_to_write[17] ),
    .D(\data_to_write[16] ),
    .Y(_04305_));
 sg13g2_nor4_1 _12026_ (.A(\data_to_write[23] ),
    .B(\data_to_write[22] ),
    .C(\data_to_write[21] ),
    .D(\data_to_write[20] ),
    .Y(_04306_));
 sg13g2_nor4_1 _12027_ (.A(\data_to_write[27] ),
    .B(\data_to_write[26] ),
    .C(\data_to_write[25] ),
    .D(\data_to_write[24] ),
    .Y(_04307_));
 sg13g2_nand3_1 _12028_ (.B(_04306_),
    .C(_04307_),
    .A(_04305_),
    .Y(_04308_));
 sg13g2_nor2_2 _12029_ (.A(\data_to_write[11] ),
    .B(\data_to_write[10] ),
    .Y(_04309_));
 sg13g2_nor3_2 _12030_ (.A(\data_to_write[11] ),
    .B(\data_to_write[10] ),
    .C(net2549),
    .Y(_04310_));
 sg13g2_nand2_2 _12031_ (.Y(_04311_),
    .A(_01796_),
    .B(_04310_));
 sg13g2_nand2_1 _12032_ (.Y(_04312_),
    .A(net2452),
    .B(_01779_));
 sg13g2_nor4_1 _12033_ (.A(net2553),
    .B(net2554),
    .C(net2555),
    .D(\crc_peri_data[2] ),
    .Y(_04313_));
 sg13g2_nor3_1 _12034_ (.A(net2551),
    .B(net2552),
    .C(_04312_),
    .Y(_04314_));
 sg13g2_nor4_1 _12035_ (.A(\data_to_write[31] ),
    .B(\data_to_write[30] ),
    .C(\data_to_write[29] ),
    .D(\data_to_write[28] ),
    .Y(_04315_));
 sg13g2_nor4_1 _12036_ (.A(net2547),
    .B(\data_to_write[15] ),
    .C(\data_to_write[14] ),
    .D(\data_to_write[13] ),
    .Y(_04316_));
 sg13g2_nand4_1 _12037_ (.B(_04314_),
    .C(_04315_),
    .A(_04313_),
    .Y(_04317_),
    .D(_04316_));
 sg13g2_nor3_1 _12038_ (.A(_04308_),
    .B(_04311_),
    .C(_04317_),
    .Y(_04318_));
 sg13g2_nor3_2 _12039_ (.A(net2325),
    .B(_02475_),
    .C(_03430_),
    .Y(_04319_));
 sg13g2_nor2b_2 _12040_ (.A(_04318_),
    .B_N(_04319_),
    .Y(_04320_));
 sg13g2_inv_4 _12041_ (.A(net2068),
    .Y(_04321_));
 sg13g2_nor2_2 _12042_ (.A(_04303_),
    .B(net2066),
    .Y(_04322_));
 sg13g2_nand2_1 _12043_ (.Y(_04323_),
    .A(_04304_),
    .B(_04321_));
 sg13g2_nor3_1 _12044_ (.A(net4395),
    .B(net5084),
    .C(net5143),
    .Y(_04324_));
 sg13g2_nor4_1 _12045_ (.A(net5157),
    .B(\i_wdt.counter[12] ),
    .C(net5136),
    .D(net5011),
    .Y(_04325_));
 sg13g2_nand3_1 _12046_ (.B(_04324_),
    .C(_04325_),
    .A(_04298_),
    .Y(_04326_));
 sg13g2_and2_1 _12047_ (.A(net5291),
    .B(net2638),
    .X(_04327_));
 sg13g2_nor4_1 _12048_ (.A(net5027),
    .B(net4817),
    .C(net5105),
    .D(net5173),
    .Y(_04328_));
 sg13g2_nor4_1 _12049_ (.A(net4893),
    .B(net5117),
    .C(net5210),
    .D(net5102),
    .Y(_04329_));
 sg13g2_nor4_1 _12050_ (.A(\i_wdt.counter[6] ),
    .B(net4717),
    .C(net4628),
    .D(net5152),
    .Y(_04330_));
 sg13g2_nand4_1 _12051_ (.B(_04328_),
    .C(_04329_),
    .A(_04327_),
    .Y(_04331_),
    .D(_04330_));
 sg13g2_nor4_2 _12052_ (.A(_04296_),
    .B(net1885),
    .C(net5216),
    .Y(_00378_),
    .D(_04331_));
 sg13g2_xnor2_1 _12053_ (.Y(_04332_),
    .A(net4674),
    .B(net2303));
 sg13g2_nor2_1 _12054_ (.A(net2425),
    .B(_04332_),
    .Y(_00379_));
 sg13g2_a21oi_1 _12055_ (.A1(\session_ms_div[0] ),
    .A2(net2302),
    .Y(_04333_),
    .B1(net3746));
 sg13g2_nand3_1 _12056_ (.B(\session_ms_div[0] ),
    .C(net2302),
    .A(net3746),
    .Y(_04334_));
 sg13g2_inv_1 _12057_ (.Y(_04335_),
    .A(_04334_));
 sg13g2_nor3_1 _12058_ (.A(net2425),
    .B(net3747),
    .C(_04335_),
    .Y(_00380_));
 sg13g2_nand3_1 _12059_ (.B(net3746),
    .C(net4674),
    .A(net3416),
    .Y(_04336_));
 sg13g2_o21ai_1 _12060_ (.B1(net2672),
    .Y(_04337_),
    .A1(net3416),
    .A2(_04335_));
 sg13g2_a21oi_1 _12061_ (.A1(net3416),
    .A2(_04335_),
    .Y(_00381_),
    .B1(_04337_));
 sg13g2_nand2b_2 _12062_ (.Y(_04338_),
    .B(net2672),
    .A_N(net2303));
 sg13g2_nand2b_1 _12063_ (.Y(_04339_),
    .B(\session_ms_div[7] ),
    .A_N(\session_ms_div[4] ));
 sg13g2_nand4_1 _12064_ (.B(\session_ms_div[8] ),
    .C(\session_ms_div[6] ),
    .A(\session_ms_div[9] ),
    .Y(_04340_),
    .D(\session_ms_div[5] ));
 sg13g2_nor4_1 _12065_ (.A(\session_ms_div[3] ),
    .B(_04336_),
    .C(_04339_),
    .D(_04340_),
    .Y(_04341_));
 sg13g2_nor2_1 _12066_ (.A(net2426),
    .B(_04341_),
    .Y(_04342_));
 sg13g2_nor2_1 _12067_ (.A(_01987_),
    .B(_04336_),
    .Y(_04343_));
 sg13g2_xnor2_1 _12068_ (.Y(_04344_),
    .A(net4829),
    .B(_04336_));
 sg13g2_nand3_1 _12069_ (.B(_04342_),
    .C(_04344_),
    .A(net2303),
    .Y(_04345_));
 sg13g2_o21ai_1 _12070_ (.B1(_04345_),
    .Y(_00382_),
    .A1(_01987_),
    .A2(_04338_));
 sg13g2_a21oi_1 _12071_ (.A1(net2303),
    .A2(_04343_),
    .Y(_04346_),
    .B1(net3710));
 sg13g2_and3_1 _12072_ (.X(_04347_),
    .A(net3710),
    .B(net2303),
    .C(_04343_));
 sg13g2_nor3_1 _12073_ (.A(net2426),
    .B(net3711),
    .C(_04347_),
    .Y(_00383_));
 sg13g2_a21oi_1 _12074_ (.A1(_04342_),
    .A2(_04347_),
    .Y(_04348_),
    .B1(net3830));
 sg13g2_and2_1 _12075_ (.A(net3830),
    .B(_04347_),
    .X(_04349_));
 sg13g2_and2_1 _12076_ (.A(net2303),
    .B(_04341_),
    .X(_04350_));
 sg13g2_nand2b_1 _12077_ (.Y(_04351_),
    .B(net2672),
    .A_N(_04350_));
 sg13g2_nor3_1 _12078_ (.A(_04348_),
    .B(_04349_),
    .C(_04351_),
    .Y(_00384_));
 sg13g2_nor2_1 _12079_ (.A(net4520),
    .B(_04349_),
    .Y(_04352_));
 sg13g2_and2_1 _12080_ (.A(net4520),
    .B(_04349_),
    .X(_04353_));
 sg13g2_nor3_1 _12081_ (.A(_04351_),
    .B(_04352_),
    .C(_04353_),
    .Y(_00385_));
 sg13g2_nor2b_1 _12082_ (.A(_04350_),
    .B_N(net3514),
    .Y(_04354_));
 sg13g2_o21ai_1 _12083_ (.B1(net2672),
    .Y(_04355_),
    .A1(_04353_),
    .A2(_04354_));
 sg13g2_a21oi_1 _12084_ (.A1(net3514),
    .A2(_04353_),
    .Y(_00386_),
    .B1(_04355_));
 sg13g2_and3_1 _12085_ (.X(_04356_),
    .A(net3755),
    .B(net3514),
    .C(_04353_));
 sg13g2_a21oi_1 _12086_ (.A1(net3514),
    .A2(_04353_),
    .Y(_04357_),
    .B1(net3755));
 sg13g2_nor3_1 _12087_ (.A(_04351_),
    .B(_04356_),
    .C(net3756),
    .Y(_00387_));
 sg13g2_nor2b_1 _12088_ (.A(_04350_),
    .B_N(net3414),
    .Y(_04358_));
 sg13g2_o21ai_1 _12089_ (.B1(net2672),
    .Y(_04359_),
    .A1(_04356_),
    .A2(_04358_));
 sg13g2_a21oi_1 _12090_ (.A1(net3414),
    .A2(_04356_),
    .Y(_00388_),
    .B1(_04359_));
 sg13g2_xnor2_1 _12091_ (.Y(_04360_),
    .A(net3899),
    .B(_04350_));
 sg13g2_nor2_1 _12092_ (.A(net2429),
    .B(_04360_),
    .Y(_00389_));
 sg13g2_a21oi_1 _12093_ (.A1(net3899),
    .A2(_04350_),
    .Y(_04361_),
    .B1(net3789));
 sg13g2_nand3_1 _12094_ (.B(net3899),
    .C(_04350_),
    .A(net3789),
    .Y(_04362_));
 sg13g2_nand2_1 _12095_ (.Y(_04363_),
    .A(net2656),
    .B(_04362_));
 sg13g2_nor2_1 _12096_ (.A(_04361_),
    .B(_04363_),
    .Y(_00390_));
 sg13g2_and2_1 _12097_ (.A(_01927_),
    .B(_04362_),
    .X(_04364_));
 sg13g2_nor2_2 _12098_ (.A(_01927_),
    .B(_04362_),
    .Y(_04365_));
 sg13g2_nor3_1 _12099_ (.A(net2429),
    .B(_04364_),
    .C(_04365_),
    .Y(_00391_));
 sg13g2_xnor2_1 _12100_ (.Y(_04366_),
    .A(net4138),
    .B(_04365_));
 sg13g2_nor2_1 _12101_ (.A(net2429),
    .B(_04366_),
    .Y(_00392_));
 sg13g2_a21oi_1 _12102_ (.A1(\i_seal.session_ctr_in[3] ),
    .A2(_04365_),
    .Y(_04367_),
    .B1(net3779));
 sg13g2_nand3_1 _12103_ (.B(net4138),
    .C(_04365_),
    .A(net3779),
    .Y(_04368_));
 sg13g2_nand2_1 _12104_ (.Y(_04369_),
    .A(net2656),
    .B(_04368_));
 sg13g2_nor2_1 _12105_ (.A(net3780),
    .B(_04369_),
    .Y(_00393_));
 sg13g2_and2_1 _12106_ (.A(_01924_),
    .B(_04368_),
    .X(_04370_));
 sg13g2_nor2_1 _12107_ (.A(_01924_),
    .B(_04368_),
    .Y(_04371_));
 sg13g2_nor3_1 _12108_ (.A(net2429),
    .B(_04370_),
    .C(_04371_),
    .Y(_00394_));
 sg13g2_o21ai_1 _12109_ (.B1(_01923_),
    .Y(_04372_),
    .A1(_01924_),
    .A2(_04368_));
 sg13g2_nand2_1 _12110_ (.Y(_04373_),
    .A(net3928),
    .B(_04371_));
 sg13g2_and3_1 _12111_ (.X(_00395_),
    .A(net2655),
    .B(_04372_),
    .C(_04373_));
 sg13g2_o21ai_1 _12112_ (.B1(net2655),
    .Y(_04374_),
    .A1(_01922_),
    .A2(_04373_));
 sg13g2_a21oi_1 _12113_ (.A1(_01922_),
    .A2(_04373_),
    .Y(_00396_),
    .B1(_04374_));
 sg13g2_nor2b_2 _12114_ (.A(pps_prev),
    .B_N(net3413),
    .Y(_04375_));
 sg13g2_nor2_1 _12115_ (.A(net4692),
    .B(_04375_),
    .Y(_04376_));
 sg13g2_a21oi_1 _12116_ (.A1(net4692),
    .A2(_04375_),
    .Y(_04377_),
    .B1(net2418));
 sg13g2_nor2b_1 _12117_ (.A(net4693),
    .B_N(_04377_),
    .Y(_00397_));
 sg13g2_a21oi_1 _12118_ (.A1(\pps_count[0] ),
    .A2(_04375_),
    .Y(_04378_),
    .B1(net4041));
 sg13g2_and3_1 _12119_ (.X(_04379_),
    .A(net4041),
    .B(net4692),
    .C(_04375_));
 sg13g2_nor3_1 _12120_ (.A(net2418),
    .B(net4042),
    .C(_04379_),
    .Y(_00398_));
 sg13g2_and2_1 _12121_ (.A(net4882),
    .B(_04379_),
    .X(_04380_));
 sg13g2_o21ai_1 _12122_ (.B1(net2641),
    .Y(_04381_),
    .A1(net4882),
    .A2(_04379_));
 sg13g2_nor2_1 _12123_ (.A(_04380_),
    .B(net4883),
    .Y(_00399_));
 sg13g2_and2_1 _12124_ (.A(net4853),
    .B(_04380_),
    .X(_04382_));
 sg13g2_o21ai_1 _12125_ (.B1(net2642),
    .Y(_04383_),
    .A1(net4853),
    .A2(_04380_));
 sg13g2_nor2_1 _12126_ (.A(_04382_),
    .B(net4854),
    .Y(_00400_));
 sg13g2_and2_1 _12127_ (.A(net4856),
    .B(_04382_),
    .X(_04384_));
 sg13g2_o21ai_1 _12128_ (.B1(net2642),
    .Y(_04385_),
    .A1(net4856),
    .A2(_04382_));
 sg13g2_nor2_1 _12129_ (.A(_04384_),
    .B(net4857),
    .Y(_00401_));
 sg13g2_xnor2_1 _12130_ (.Y(_04386_),
    .A(net4789),
    .B(_04384_));
 sg13g2_nor2_1 _12131_ (.A(net2421),
    .B(net4790),
    .Y(_00402_));
 sg13g2_a21oi_1 _12132_ (.A1(\pps_count[5] ),
    .A2(_04384_),
    .Y(_04387_),
    .B1(net4009));
 sg13g2_and3_1 _12133_ (.X(_04388_),
    .A(net4009),
    .B(net4789),
    .C(_04384_));
 sg13g2_nor3_1 _12134_ (.A(net2421),
    .B(net4010),
    .C(_04388_),
    .Y(_00403_));
 sg13g2_and2_1 _12135_ (.A(net4926),
    .B(_04388_),
    .X(_04389_));
 sg13g2_o21ai_1 _12136_ (.B1(net2642),
    .Y(_04390_),
    .A1(net4926),
    .A2(_04388_));
 sg13g2_nor2_1 _12137_ (.A(_04389_),
    .B(_04390_),
    .Y(_00404_));
 sg13g2_and2_1 _12138_ (.A(net4888),
    .B(_04389_),
    .X(_04391_));
 sg13g2_o21ai_1 _12139_ (.B1(net2641),
    .Y(_04392_),
    .A1(net4888),
    .A2(_04389_));
 sg13g2_nor2_1 _12140_ (.A(_04391_),
    .B(net4889),
    .Y(_00405_));
 sg13g2_xnor2_1 _12141_ (.Y(_04393_),
    .A(net4727),
    .B(_04391_));
 sg13g2_nor2_1 _12142_ (.A(net2418),
    .B(net4728),
    .Y(_00406_));
 sg13g2_a21oi_1 _12143_ (.A1(\pps_count[9] ),
    .A2(_04391_),
    .Y(_04394_),
    .B1(net4023));
 sg13g2_and3_1 _12144_ (.X(_04395_),
    .A(net4023),
    .B(net4727),
    .C(_04391_));
 sg13g2_nor3_1 _12145_ (.A(net2419),
    .B(net4024),
    .C(_04395_),
    .Y(_00407_));
 sg13g2_and2_1 _12146_ (.A(net4919),
    .B(_04395_),
    .X(_04396_));
 sg13g2_o21ai_1 _12147_ (.B1(net2636),
    .Y(_04397_),
    .A1(net4919),
    .A2(_04395_));
 sg13g2_nor2_1 _12148_ (.A(_04396_),
    .B(_04397_),
    .Y(_00408_));
 sg13g2_o21ai_1 _12149_ (.B1(net2636),
    .Y(_04398_),
    .A1(net3570),
    .A2(_04396_));
 sg13g2_a21oi_1 _12150_ (.A1(net3570),
    .A2(_04396_),
    .Y(_00409_),
    .B1(_04398_));
 sg13g2_a21oi_1 _12151_ (.A1(net3570),
    .A2(_04396_),
    .Y(_04399_),
    .B1(net3857));
 sg13g2_and3_1 _12152_ (.X(_04400_),
    .A(net3857),
    .B(net3570),
    .C(_04396_));
 sg13g2_nor3_1 _12153_ (.A(net2418),
    .B(net3858),
    .C(_04400_),
    .Y(_00410_));
 sg13g2_nand2_1 _12154_ (.Y(_04401_),
    .A(net4917),
    .B(_04400_));
 sg13g2_o21ai_1 _12155_ (.B1(net2636),
    .Y(_04402_),
    .A1(net4917),
    .A2(_04400_));
 sg13g2_nor2b_1 _12156_ (.A(_04402_),
    .B_N(_04401_),
    .Y(_00411_));
 sg13g2_o21ai_1 _12157_ (.B1(net2635),
    .Y(_04403_),
    .A1(_01986_),
    .A2(_04401_));
 sg13g2_a21oi_1 _12158_ (.A1(_01986_),
    .A2(_04401_),
    .Y(_00412_),
    .B1(_04403_));
 sg13g2_and2_1 _12159_ (.A(net2639),
    .B(net2),
    .X(_00413_));
 sg13g2_and2_1 _12160_ (.A(net2635),
    .B(net4081),
    .X(_00414_));
 sg13g2_and2_1 _12161_ (.A(net2634),
    .B(net6),
    .X(_00415_));
 sg13g2_and2_1 _12162_ (.A(net2635),
    .B(net3411),
    .X(_00416_));
 sg13g2_nor4_1 _12163_ (.A(\timer_count[9] ),
    .B(\timer_count[8] ),
    .C(\timer_count[7] ),
    .D(\timer_count[4] ),
    .Y(_04404_));
 sg13g2_nor4_1 _12164_ (.A(net4333),
    .B(\timer_count[10] ),
    .C(\timer_count[6] ),
    .D(\timer_count[5] ),
    .Y(_04405_));
 sg13g2_nand2_1 _12165_ (.Y(_04406_),
    .A(_04404_),
    .B(_04405_));
 sg13g2_nor3_1 _12166_ (.A(\timer_count[3] ),
    .B(\timer_count[2] ),
    .C(\timer_count[1] ),
    .Y(_04407_));
 sg13g2_nand4_1 _12167_ (.B(_04404_),
    .C(_04405_),
    .A(_01985_),
    .Y(_04408_),
    .D(_04407_));
 sg13g2_nor4_1 _12168_ (.A(\timer_count[15] ),
    .B(\timer_count[14] ),
    .C(\timer_count[13] ),
    .D(net5387),
    .Y(_04409_));
 sg13g2_nor3_1 _12169_ (.A(net4755),
    .B(\timer_count[17] ),
    .C(\timer_count[16] ),
    .Y(_04410_));
 sg13g2_nor3_1 _12170_ (.A(\timer_count[21] ),
    .B(\timer_count[20] ),
    .C(\timer_count[19] ),
    .Y(_04411_));
 sg13g2_nand3_1 _12171_ (.B(_04410_),
    .C(_04411_),
    .A(_04409_),
    .Y(_04412_));
 sg13g2_inv_1 _12172_ (.Y(_04413_),
    .A(_04412_));
 sg13g2_nor4_1 _12173_ (.A(\timer_count[30] ),
    .B(\timer_count[29] ),
    .C(\timer_count[28] ),
    .D(\timer_count[27] ),
    .Y(_04414_));
 sg13g2_nor2_1 _12174_ (.A(\timer_count[26] ),
    .B(\timer_count[25] ),
    .Y(_04415_));
 sg13g2_nor4_1 _12175_ (.A(\timer_count[31] ),
    .B(\timer_count[24] ),
    .C(\timer_count[23] ),
    .D(\timer_count[22] ),
    .Y(_04416_));
 sg13g2_nand4_1 _12176_ (.B(_04414_),
    .C(_04415_),
    .A(_04413_),
    .Y(_04417_),
    .D(_04416_));
 sg13g2_o21ai_1 _12177_ (.B1(net2302),
    .Y(_04418_),
    .A1(_04408_),
    .A2(_04417_));
 sg13g2_nor2_1 _12178_ (.A(\timer_count[0] ),
    .B(net2113),
    .Y(_04419_));
 sg13g2_xnor2_1 _12179_ (.Y(_04420_),
    .A(_01985_),
    .B(net2113));
 sg13g2_nor3_1 _12180_ (.A(net2325),
    .B(_03430_),
    .C(_03431_),
    .Y(_04421_));
 sg13g2_nand2_2 _12181_ (.Y(_04422_),
    .A(net2326),
    .B(net2121));
 sg13g2_or3_1 _12182_ (.A(net2325),
    .B(_03431_),
    .C(_03476_),
    .X(_04423_));
 sg13g2_nand2_1 _12183_ (.Y(_04424_),
    .A(net2645),
    .B(_04423_));
 sg13g2_nand2_2 _12184_ (.Y(_04425_),
    .A(net2559),
    .B(net2638));
 sg13g2_a22oi_1 _12185_ (.Y(_00417_),
    .B1(net2058),
    .B2(_04425_),
    .A2(net2060),
    .A1(_04420_));
 sg13g2_nor3_1 _12186_ (.A(net5131),
    .B(net5388),
    .C(net2113),
    .Y(_04426_));
 sg13g2_xnor2_1 _12187_ (.Y(_04427_),
    .A(net5131),
    .B(_04419_));
 sg13g2_nand2_1 _12188_ (.Y(_04428_),
    .A(net2557),
    .B(net2639));
 sg13g2_a22oi_1 _12189_ (.Y(_00418_),
    .B1(_04428_),
    .B2(net2058),
    .A2(net5132),
    .A1(net2061));
 sg13g2_nand2_2 _12190_ (.Y(_04429_),
    .A(net5012),
    .B(net2638));
 sg13g2_nand2b_2 _12191_ (.Y(_04430_),
    .B(_04426_),
    .A_N(net5018));
 sg13g2_xnor2_1 _12192_ (.Y(_04431_),
    .A(net5018),
    .B(_04426_));
 sg13g2_a22oi_1 _12193_ (.Y(_00419_),
    .B1(net5019),
    .B2(net2060),
    .A2(_04429_),
    .A1(net2057));
 sg13g2_xor2_1 _12194_ (.B(_04430_),
    .A(net5251),
    .X(_04432_));
 sg13g2_nand2_2 _12195_ (.Y(_04433_),
    .A(net2555),
    .B(net2637));
 sg13g2_a22oi_1 _12196_ (.Y(_00420_),
    .B1(_04433_),
    .B2(net2058),
    .A2(net5252),
    .A1(net2060));
 sg13g2_nand2_2 _12197_ (.Y(_04434_),
    .A(net2554),
    .B(net2633));
 sg13g2_nor3_1 _12198_ (.A(net5330),
    .B(net5251),
    .C(_04430_),
    .Y(_04435_));
 sg13g2_o21ai_1 _12199_ (.B1(net5330),
    .Y(_04436_),
    .A1(net5251),
    .A2(_04430_));
 sg13g2_nor2b_1 _12200_ (.A(_04435_),
    .B_N(_04436_),
    .Y(_04437_));
 sg13g2_a22oi_1 _12201_ (.Y(_00421_),
    .B1(_04437_),
    .B2(net2060),
    .A2(_04434_),
    .A1(net2057));
 sg13g2_nand2_2 _12202_ (.Y(_04438_),
    .A(net2553),
    .B(net2633));
 sg13g2_nor2b_1 _12203_ (.A(net5063),
    .B_N(_04435_),
    .Y(_04439_));
 sg13g2_xnor2_1 _12204_ (.Y(_04440_),
    .A(net5063),
    .B(_04435_));
 sg13g2_a22oi_1 _12205_ (.Y(_00422_),
    .B1(net5064),
    .B2(net2060),
    .A2(_04438_),
    .A1(net2057));
 sg13g2_nand2_2 _12206_ (.Y(_04441_),
    .A(net2552),
    .B(net2633));
 sg13g2_nand2b_2 _12207_ (.Y(_04442_),
    .B(_04439_),
    .A_N(net5108));
 sg13g2_xnor2_1 _12208_ (.Y(_04443_),
    .A(net5108),
    .B(_04439_));
 sg13g2_a22oi_1 _12209_ (.Y(_00423_),
    .B1(net5109),
    .B2(net2060),
    .A2(_04441_),
    .A1(net2057));
 sg13g2_nand2_2 _12210_ (.Y(_04444_),
    .A(net2551),
    .B(net2633));
 sg13g2_xor2_1 _12211_ (.B(_04442_),
    .A(net5229),
    .X(_04445_));
 sg13g2_a22oi_1 _12212_ (.Y(_00424_),
    .B1(_04445_),
    .B2(net2060),
    .A2(_04444_),
    .A1(net2057));
 sg13g2_o21ai_1 _12213_ (.B1(net5218),
    .Y(_04446_),
    .A1(\timer_count[7] ),
    .A2(_04442_));
 sg13g2_nor3_1 _12214_ (.A(net5218),
    .B(\timer_count[7] ),
    .C(_04442_),
    .Y(_04447_));
 sg13g2_nand2_1 _12215_ (.Y(_04448_),
    .A(net2060),
    .B(_04446_));
 sg13g2_nor2_1 _12216_ (.A(net5219),
    .B(_04448_),
    .Y(_04449_));
 sg13g2_nand2_2 _12217_ (.Y(_04450_),
    .A(net2549),
    .B(net2637));
 sg13g2_a21oi_1 _12218_ (.A1(net2057),
    .A2(_04450_),
    .Y(_00425_),
    .B1(net5220));
 sg13g2_nor4_1 _12219_ (.A(net5353),
    .B(net5218),
    .C(net5229),
    .D(_04442_),
    .Y(_04451_));
 sg13g2_nor2b_1 _12220_ (.A(net5219),
    .B_N(net5353),
    .Y(_04452_));
 sg13g2_nor3_1 _12221_ (.A(net2112),
    .B(_04451_),
    .C(_04452_),
    .Y(_04453_));
 sg13g2_nand2_2 _12222_ (.Y(_04454_),
    .A(net2548),
    .B(net2637));
 sg13g2_a21oi_1 _12223_ (.A1(net2057),
    .A2(_04454_),
    .Y(_00426_),
    .B1(_04453_));
 sg13g2_nor2b_1 _12224_ (.A(\timer_count[10] ),
    .B_N(_04451_),
    .Y(_04455_));
 sg13g2_xnor2_1 _12225_ (.Y(_04456_),
    .A(net5129),
    .B(_04451_));
 sg13g2_nand2_1 _12226_ (.Y(_04457_),
    .A(net4958),
    .B(net2633));
 sg13g2_a22oi_1 _12227_ (.Y(_00427_),
    .B1(_04457_),
    .B2(net2057),
    .A2(net5130),
    .A1(_04423_));
 sg13g2_nand2b_1 _12228_ (.Y(_04458_),
    .B(net4333),
    .A_N(_04455_));
 sg13g2_nor2_1 _12229_ (.A(_04408_),
    .B(net2113),
    .Y(_04459_));
 sg13g2_nor2_1 _12230_ (.A(net2112),
    .B(_04459_),
    .Y(_04460_));
 sg13g2_a221oi_1 _12231_ (.B2(_04460_),
    .C1(net2415),
    .B1(net4334),
    .A1(_01794_),
    .Y(_00428_),
    .A2(net2112));
 sg13g2_nor3_1 _12232_ (.A(net5154),
    .B(_04408_),
    .C(net2113),
    .Y(_04461_));
 sg13g2_xnor2_1 _12233_ (.Y(_04462_),
    .A(net5154),
    .B(_04459_));
 sg13g2_nand2_1 _12234_ (.Y(_04463_),
    .A(net2547),
    .B(net2637));
 sg13g2_a22oi_1 _12235_ (.Y(_00429_),
    .B1(_04463_),
    .B2(net2058),
    .A2(_04462_),
    .A1(net2061));
 sg13g2_nand2_1 _12236_ (.Y(_04464_),
    .A(\data_to_write[13] ),
    .B(net2635));
 sg13g2_nand2b_1 _12237_ (.Y(_04465_),
    .B(_04461_),
    .A_N(net5036));
 sg13g2_xnor2_1 _12238_ (.Y(_04466_),
    .A(net5036),
    .B(_04461_));
 sg13g2_a22oi_1 _12239_ (.Y(_00430_),
    .B1(net5037),
    .B2(_04423_),
    .A2(_04464_),
    .A1(net2058));
 sg13g2_xor2_1 _12240_ (.B(_04465_),
    .A(net5178),
    .X(_04467_));
 sg13g2_nand2_1 _12241_ (.Y(_04468_),
    .A(net4962),
    .B(net2635));
 sg13g2_a22oi_1 _12242_ (.Y(_00431_),
    .B1(_04468_),
    .B2(net2058),
    .A2(_04467_),
    .A1(net2061));
 sg13g2_o21ai_1 _12243_ (.B1(net4385),
    .Y(_04469_),
    .A1(\timer_count[14] ),
    .A2(_04465_));
 sg13g2_and2_1 _12244_ (.A(_04409_),
    .B(_04459_),
    .X(_04470_));
 sg13g2_inv_1 _12245_ (.Y(_04471_),
    .A(_04470_));
 sg13g2_nor2_1 _12246_ (.A(net2112),
    .B(_04470_),
    .Y(_04472_));
 sg13g2_a221oi_1 _12247_ (.B2(_04472_),
    .C1(net2422),
    .B1(net4386),
    .A1(_01790_),
    .Y(_00432_),
    .A2(net2112));
 sg13g2_nand2b_2 _12248_ (.Y(_04473_),
    .B(_04470_),
    .A_N(net5072));
 sg13g2_a21oi_1 _12249_ (.A1(net5072),
    .A2(_04471_),
    .Y(_04474_),
    .B1(net2110));
 sg13g2_a221oi_1 _12250_ (.B2(_04474_),
    .C1(net2419),
    .B1(_04473_),
    .A1(_01842_),
    .Y(_00433_),
    .A2(net2110));
 sg13g2_xor2_1 _12251_ (.B(_04473_),
    .A(\timer_count[17] ),
    .X(_04475_));
 sg13g2_nand2_1 _12252_ (.Y(_04476_),
    .A(net4914),
    .B(net2636));
 sg13g2_nand3_1 _12253_ (.B(net2636),
    .C(net2112),
    .A(net4914),
    .Y(_04477_));
 sg13g2_o21ai_1 _12254_ (.B1(_04477_),
    .Y(_00434_),
    .A1(net2059),
    .A2(_04475_));
 sg13g2_o21ai_1 _12255_ (.B1(net4755),
    .Y(_04478_),
    .A1(\timer_count[17] ),
    .A2(_04473_));
 sg13g2_a21oi_1 _12256_ (.A1(_04410_),
    .A2(_04470_),
    .Y(_04479_),
    .B1(net2110));
 sg13g2_nor3_1 _12257_ (.A(net4755),
    .B(\timer_count[17] ),
    .C(_04473_),
    .Y(_04480_));
 sg13g2_a221oi_1 _12258_ (.B2(_04479_),
    .C1(net2419),
    .B1(net4756),
    .A1(_01838_),
    .Y(_00435_),
    .A2(net2110));
 sg13g2_nand2b_1 _12259_ (.Y(_04481_),
    .B(_04480_),
    .A_N(\timer_count[19] ));
 sg13g2_xnor2_1 _12260_ (.Y(_04482_),
    .A(\timer_count[19] ),
    .B(_04480_));
 sg13g2_nand3_1 _12261_ (.B(net2636),
    .C(net2110),
    .A(net4912),
    .Y(_04483_));
 sg13g2_o21ai_1 _12262_ (.B1(_04483_),
    .Y(_00436_),
    .A1(net2059),
    .A2(_04482_));
 sg13g2_o21ai_1 _12263_ (.B1(_04423_),
    .Y(_04484_),
    .A1(net4799),
    .A2(_04481_));
 sg13g2_a21oi_1 _12264_ (.A1(net4799),
    .A2(_04481_),
    .Y(_04485_),
    .B1(_04484_));
 sg13g2_o21ai_1 _12265_ (.B1(net2640),
    .Y(_04486_),
    .A1(\data_to_write[20] ),
    .A2(_04422_));
 sg13g2_nor2_1 _12266_ (.A(net4800),
    .B(_04486_),
    .Y(_00437_));
 sg13g2_or2_1 _12267_ (.X(_04487_),
    .B(_04412_),
    .A(_04408_));
 sg13g2_or2_1 _12268_ (.X(_04488_),
    .B(_04487_),
    .A(net2113));
 sg13g2_nand2_1 _12269_ (.Y(_04489_),
    .A(net2062),
    .B(_04488_));
 sg13g2_o21ai_1 _12270_ (.B1(_04489_),
    .Y(_04490_),
    .A1(net4933),
    .A2(net2062));
 sg13g2_or2_1 _12271_ (.X(_04491_),
    .B(net2111),
    .A(_04418_));
 sg13g2_o21ai_1 _12272_ (.B1(_04490_),
    .Y(_04492_),
    .A1(_01984_),
    .A2(_04484_));
 sg13g2_and2_1 _12273_ (.A(net2640),
    .B(_04492_),
    .X(_00438_));
 sg13g2_nand2_1 _12274_ (.Y(_04493_),
    .A(net4462),
    .B(_04488_));
 sg13g2_o21ai_1 _12275_ (.B1(net2062),
    .Y(_04494_),
    .A1(net4462),
    .A2(_04488_));
 sg13g2_inv_1 _12276_ (.Y(_04495_),
    .A(_04494_));
 sg13g2_a221oi_1 _12277_ (.B2(_04495_),
    .C1(net2420),
    .B1(_04493_),
    .A1(_01830_),
    .Y(_00439_),
    .A2(net2111));
 sg13g2_nor4_1 _12278_ (.A(net5134),
    .B(net4462),
    .C(_04487_),
    .D(_04491_),
    .Y(_04496_));
 sg13g2_a221oi_1 _12279_ (.B2(net5134),
    .C1(_04496_),
    .B1(_04495_),
    .A1(net4928),
    .Y(_04497_),
    .A2(net2111));
 sg13g2_nor2_1 _12280_ (.A(net2420),
    .B(_04497_),
    .Y(_00440_));
 sg13g2_nor4_1 _12281_ (.A(net5287),
    .B(net5134),
    .C(net4462),
    .D(_04487_),
    .Y(_04498_));
 sg13g2_nand2b_2 _12282_ (.Y(_04499_),
    .B(_04498_),
    .A_N(net2113));
 sg13g2_o21ai_1 _12283_ (.B1(net2640),
    .Y(_04500_),
    .A1(net4986),
    .A2(net2062));
 sg13g2_nor2_1 _12284_ (.A(net5287),
    .B(net2111),
    .Y(_04501_));
 sg13g2_or3_1 _12285_ (.A(_04496_),
    .B(_04500_),
    .C(_04501_),
    .X(_04502_));
 sg13g2_o21ai_1 _12286_ (.B1(_04502_),
    .Y(_00441_),
    .A1(net2059),
    .A2(_04499_));
 sg13g2_nor2_1 _12287_ (.A(\timer_count[25] ),
    .B(_04499_),
    .Y(_04503_));
 sg13g2_xor2_1 _12288_ (.B(_04499_),
    .A(net5186),
    .X(_04504_));
 sg13g2_nand2_1 _12289_ (.Y(_04505_),
    .A(net5071),
    .B(net2640));
 sg13g2_a22oi_1 _12290_ (.Y(_00442_),
    .B1(_04505_),
    .B2(net2059),
    .A2(net5187),
    .A1(net2062));
 sg13g2_xnor2_1 _12291_ (.Y(_04506_),
    .A(net4970),
    .B(_04503_));
 sg13g2_o21ai_1 _12292_ (.B1(net2641),
    .Y(_04507_),
    .A1(\data_to_write[26] ),
    .A2(net2062));
 sg13g2_a21oi_1 _12293_ (.A1(net2062),
    .A2(net4971),
    .Y(_00443_),
    .B1(_04507_));
 sg13g2_nand2_1 _12294_ (.Y(_04508_),
    .A(_04415_),
    .B(_04498_));
 sg13g2_or2_1 _12295_ (.X(_04509_),
    .B(_04508_),
    .A(net5174));
 sg13g2_and2_1 _12296_ (.A(_04418_),
    .B(_04423_),
    .X(_04510_));
 sg13g2_nand2_1 _12297_ (.Y(_04511_),
    .A(net5174),
    .B(_04508_));
 sg13g2_a21oi_1 _12298_ (.A1(_04509_),
    .A2(_04511_),
    .Y(_04512_),
    .B1(_04491_));
 sg13g2_a221oi_1 _12299_ (.B2(net5174),
    .C1(_04512_),
    .B1(_04510_),
    .A1(net5079),
    .Y(_04513_),
    .A2(net2111));
 sg13g2_nor2_1 _12300_ (.A(net2419),
    .B(_04513_),
    .Y(_00444_));
 sg13g2_xor2_1 _12301_ (.B(_04509_),
    .A(net5207),
    .X(_04514_));
 sg13g2_nor2_1 _12302_ (.A(_04491_),
    .B(_04514_),
    .Y(_04515_));
 sg13g2_a221oi_1 _12303_ (.B2(net5207),
    .C1(_04515_),
    .B1(_04510_),
    .A1(net4927),
    .Y(_04516_),
    .A2(net2110));
 sg13g2_nor2_1 _12304_ (.A(net2419),
    .B(_04516_),
    .Y(_00445_));
 sg13g2_nor3_1 _12305_ (.A(net5322),
    .B(net5207),
    .C(_04509_),
    .Y(_04517_));
 sg13g2_o21ai_1 _12306_ (.B1(net5322),
    .Y(_04518_),
    .A1(\timer_count[28] ),
    .A2(_04509_));
 sg13g2_nor2b_1 _12307_ (.A(_04517_),
    .B_N(_04518_),
    .Y(_04519_));
 sg13g2_a22oi_1 _12308_ (.Y(_04520_),
    .B1(_04510_),
    .B2(net5322),
    .A2(net2110),
    .A1(net5055));
 sg13g2_o21ai_1 _12309_ (.B1(_04520_),
    .Y(_04521_),
    .A1(_04491_),
    .A2(_04519_));
 sg13g2_and2_1 _12310_ (.A(net2640),
    .B(_04521_),
    .X(_00446_));
 sg13g2_nand3_1 _12311_ (.B(_04415_),
    .C(_04498_),
    .A(_04414_),
    .Y(_04522_));
 sg13g2_xnor2_1 _12312_ (.Y(_04523_),
    .A(net5329),
    .B(_04517_));
 sg13g2_a22oi_1 _12313_ (.Y(_04524_),
    .B1(_04510_),
    .B2(net5329),
    .A2(net2110),
    .A1(net5005));
 sg13g2_o21ai_1 _12314_ (.B1(_04524_),
    .Y(_04525_),
    .A1(_04491_),
    .A2(_04523_));
 sg13g2_and2_1 _12315_ (.A(net2640),
    .B(_04525_),
    .X(_00447_));
 sg13g2_xor2_1 _12316_ (.B(_04522_),
    .A(net5318),
    .X(_04526_));
 sg13g2_a22oi_1 _12317_ (.Y(_04527_),
    .B1(_04510_),
    .B2(net5318),
    .A2(net2111),
    .A1(net5020));
 sg13g2_o21ai_1 _12318_ (.B1(_04527_),
    .Y(_04528_),
    .A1(_04491_),
    .A2(_04526_));
 sg13g2_and2_1 _12319_ (.A(net2640),
    .B(net5319),
    .X(_00448_));
 sg13g2_nand2_1 _12320_ (.Y(_04529_),
    .A(\timer_count[0] ),
    .B(_04407_));
 sg13g2_nor4_1 _12321_ (.A(_04406_),
    .B(_04417_),
    .C(net2113),
    .D(_04529_),
    .Y(_04530_));
 sg13g2_nor2_1 _12322_ (.A(net4436),
    .B(_04530_),
    .Y(_04531_));
 sg13g2_nor2_1 _12323_ (.A(net2058),
    .B(net4437),
    .Y(_00449_));
 sg13g2_and2_1 _12324_ (.A(net2635),
    .B(net3413),
    .X(_00450_));
 sg13g2_nand3_1 _12325_ (.B(_01773_),
    .C(net2553),
    .A(net2551),
    .Y(_04532_));
 sg13g2_nand4_1 _12326_ (.B(net2556),
    .C(net2452),
    .A(net2453),
    .Y(_04533_),
    .D(net2559));
 sg13g2_nor4_1 _12327_ (.A(net2554),
    .B(_02473_),
    .C(_04532_),
    .D(_04533_),
    .Y(_04534_));
 sg13g2_a21oi_2 _12328_ (.B1(net4132),
    .Y(_04535_),
    .A2(_04534_),
    .A1(net2074));
 sg13g2_nand2_2 _12329_ (.Y(_04536_),
    .A(net1),
    .B(_04535_));
 sg13g2_nor3_1 _12330_ (.A(net3430),
    .B(_02754_),
    .C(_04536_),
    .Y(_00451_));
 sg13g2_nor3_1 _12331_ (.A(net4298),
    .B(net3430),
    .C(_02754_),
    .Y(_04537_));
 sg13g2_a21oi_1 _12332_ (.A1(net4298),
    .A2(net3430),
    .Y(_04538_),
    .B1(_04537_));
 sg13g2_nor2_1 _12333_ (.A(_04536_),
    .B(_04538_),
    .Y(_00452_));
 sg13g2_nor2b_1 _12334_ (.A(net4685),
    .B_N(_04537_),
    .Y(_04539_));
 sg13g2_xnor2_1 _12335_ (.Y(_04540_),
    .A(net4685),
    .B(_04537_));
 sg13g2_nor2_1 _12336_ (.A(_04536_),
    .B(_04540_),
    .Y(_00453_));
 sg13g2_nor2b_1 _12337_ (.A(\reset_hold_counter[3] ),
    .B_N(_04539_),
    .Y(_04541_));
 sg13g2_xnor2_1 _12338_ (.Y(_04542_),
    .A(net4739),
    .B(_04539_));
 sg13g2_nor2_1 _12339_ (.A(_04536_),
    .B(_04542_),
    .Y(_00454_));
 sg13g2_xnor2_1 _12340_ (.Y(_04543_),
    .A(net4322),
    .B(_04541_));
 sg13g2_nor2_1 _12341_ (.A(_04536_),
    .B(net4323),
    .Y(_00455_));
 sg13g2_nor4_2 _12342_ (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .C(_02810_),
    .Y(_04544_),
    .D(_03154_));
 sg13g2_nand2_2 _12343_ (.Y(_04545_),
    .A(net2320),
    .B(_04544_));
 sg13g2_inv_1 _12344_ (.Y(_04546_),
    .A(_04545_));
 sg13g2_and2_1 _12345_ (.A(net5261),
    .B(net2320),
    .X(_04547_));
 sg13g2_nor2_2 _12346_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(_04544_),
    .Y(_04548_));
 sg13g2_or2_1 _12347_ (.X(_04549_),
    .B(_04544_),
    .A(\i_tinyqv.cpu.i_core.is_interrupt ));
 sg13g2_nand2_2 _12348_ (.Y(_04550_),
    .A(net2320),
    .B(_04549_));
 sg13g2_nor2_2 _12349_ (.A(net2318),
    .B(_04548_),
    .Y(_04551_));
 sg13g2_nand2_1 _12350_ (.Y(_04552_),
    .A(net4637),
    .B(net4122));
 sg13g2_a21oi_1 _12351_ (.A1(net4357),
    .A2(net4828),
    .Y(_04553_),
    .B1(_04552_));
 sg13g2_nor3_1 _12352_ (.A(net4937),
    .B(_03385_),
    .C(_04545_),
    .Y(_04554_));
 sg13g2_a221oi_1 _12353_ (.B2(_04547_),
    .C1(_04554_),
    .B1(_04553_),
    .A1(net5137),
    .Y(_04555_),
    .A2(_04550_));
 sg13g2_nor4_1 _12354_ (.A(net4937),
    .B(_02689_),
    .C(_02719_),
    .D(_04545_),
    .Y(_04556_));
 sg13g2_nand3_1 _12355_ (.B(_02641_),
    .C(_04556_),
    .A(_02571_),
    .Y(_04557_));
 sg13g2_a21oi_1 _12356_ (.A1(net5138),
    .A2(_04557_),
    .Y(_00456_),
    .B1(net2450));
 sg13g2_a22oi_1 _12357_ (.Y(_04558_),
    .B1(net4122),
    .B2(net4637),
    .A2(\i_tinyqv.cpu.i_core.mie[0] ),
    .A1(net4357));
 sg13g2_nand2_1 _12358_ (.Y(_04559_),
    .A(net4177),
    .B(_03671_));
 sg13g2_nand3_1 _12359_ (.B(_03671_),
    .C(_04558_),
    .A(net4177),
    .Y(_04560_));
 sg13g2_o21ai_1 _12360_ (.B1(net2499),
    .Y(_04561_),
    .A1(net4670),
    .A2(_04551_));
 sg13g2_a21oi_1 _12361_ (.A1(_04547_),
    .A2(_04560_),
    .Y(_00457_),
    .B1(_04561_));
 sg13g2_nand2_1 _12362_ (.Y(_04562_),
    .A(net3774),
    .B(_04550_));
 sg13g2_a21oi_1 _12363_ (.A1(_04557_),
    .A2(_04562_),
    .Y(_00458_),
    .B1(net2450));
 sg13g2_a21oi_1 _12364_ (.A1(net4320),
    .A2(_04545_),
    .Y(_04563_),
    .B1(_04547_));
 sg13g2_nor2_1 _12365_ (.A(net2450),
    .B(net4321),
    .Y(_00459_));
 sg13g2_nand2_1 _12366_ (.Y(_04564_),
    .A(net3405),
    .B(_02753_));
 sg13g2_a21oi_1 _12367_ (.A1(_04535_),
    .A2(_04564_),
    .Y(_00460_),
    .B1(_02026_));
 sg13g2_nor2b_1 _12368_ (.A(net2612),
    .B_N(net2613),
    .Y(_04565_));
 sg13g2_and2_1 _12369_ (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(_04565_),
    .X(_04566_));
 sg13g2_and3_2 _12370_ (.X(_04567_),
    .A(net5111),
    .B(net2611),
    .C(net2299));
 sg13g2_nand3_1 _12371_ (.B(net2611),
    .C(net2299),
    .A(\i_tinyqv.cpu.instr_fetch_running ),
    .Y(_04568_));
 sg13g2_xnor2_1 _12372_ (.Y(_04569_),
    .A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .B(\i_tinyqv.cpu.i_core.cmp_out ));
 sg13g2_nor3_2 _12373_ (.A(_02810_),
    .B(_03154_),
    .C(_03374_),
    .Y(_04570_));
 sg13g2_nand4_1 _12374_ (.B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .C(_02809_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .Y(_04571_),
    .D(_03153_));
 sg13g2_nor3_1 _12375_ (.A(_02803_),
    .B(_04549_),
    .C(net2298),
    .Y(_04572_));
 sg13g2_o21ai_1 _12376_ (.B1(_04572_),
    .Y(_04573_),
    .A1(net2360),
    .A2(_04569_));
 sg13g2_and2_1 _12377_ (.A(net2317),
    .B(_04573_),
    .X(_04574_));
 sg13g2_nor2_1 _12378_ (.A(net2510),
    .B(net2315),
    .Y(_04575_));
 sg13g2_a21o_1 _12379_ (.A2(_02823_),
    .A1(_02814_),
    .B1(_04575_),
    .X(_04576_));
 sg13g2_a21oi_2 _12380_ (.B1(_01959_),
    .Y(_04577_),
    .A2(_04559_),
    .A1(_04558_));
 sg13g2_and2_1 _12381_ (.A(_02813_),
    .B(_04577_),
    .X(_04578_));
 sg13g2_nor2_1 _12382_ (.A(net2509),
    .B(\i_tinyqv.cpu.pc[1] ),
    .Y(_04579_));
 sg13g2_a21oi_1 _12383_ (.A1(net2509),
    .A2(_03630_),
    .Y(_04580_),
    .B1(_04579_));
 sg13g2_a21o_2 _12384_ (.A2(_03630_),
    .A1(net2509),
    .B1(_04579_),
    .X(_04581_));
 sg13g2_nor2_1 _12385_ (.A(net2509),
    .B(\i_tinyqv.cpu.pc[2] ),
    .Y(_04582_));
 sg13g2_a21o_2 _12386_ (.A2(_03760_),
    .A1(net2509),
    .B1(_04582_),
    .X(_04583_));
 sg13g2_a21oi_2 _12387_ (.B1(_04582_),
    .Y(_04584_),
    .A2(_03760_),
    .A1(net2512));
 sg13g2_mux4_1 _12388_ (.S0(net2288),
    .A0(\i_tinyqv.cpu.instr_data[1][1] ),
    .A1(\i_tinyqv.cpu.instr_data[0][1] ),
    .A2(\i_tinyqv.cpu.instr_data[3][1] ),
    .A3(\i_tinyqv.cpu.instr_data[2][1] ),
    .S1(net2238),
    .X(_04585_));
 sg13g2_mux4_1 _12389_ (.S0(net2291),
    .A0(\i_tinyqv.cpu.instr_data[0][0] ),
    .A1(\i_tinyqv.cpu.instr_data[1][0] ),
    .A2(\i_tinyqv.cpu.instr_data[2][0] ),
    .A3(\i_tinyqv.cpu.instr_data[3][0] ),
    .S1(net2238),
    .X(_04586_));
 sg13g2_and2_1 _12390_ (.A(net2173),
    .B(_04586_),
    .X(_04587_));
 sg13g2_nand2_2 _12391_ (.Y(_04588_),
    .A(net2173),
    .B(_04586_));
 sg13g2_nand2_1 _12392_ (.Y(_04589_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_04583_));
 sg13g2_xnor2_1 _12393_ (.Y(_04590_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_04583_));
 sg13g2_nor2_1 _12394_ (.A(_02002_),
    .B(net2291),
    .Y(_04591_));
 sg13g2_o21ai_1 _12395_ (.B1(_04588_),
    .Y(_04592_),
    .A1(_04590_),
    .A2(_04591_));
 sg13g2_nand2_1 _12396_ (.Y(_04593_),
    .A(_02002_),
    .B(net2291));
 sg13g2_nand2_1 _12397_ (.Y(_04594_),
    .A(net2512),
    .B(_03348_));
 sg13g2_xnor2_1 _12398_ (.Y(_04595_),
    .A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B(_04594_));
 sg13g2_o21ai_1 _12399_ (.B1(_04595_),
    .Y(_04596_),
    .A1(\i_tinyqv.cpu.instr_write_offset[2] ),
    .A2(_04583_));
 sg13g2_nor2_1 _12400_ (.A(_04593_),
    .B(_04595_),
    .Y(_04597_));
 sg13g2_a22oi_1 _12401_ (.Y(_04598_),
    .B1(_04597_),
    .B2(_04589_),
    .A2(_04593_),
    .A1(_04590_));
 sg13g2_nand3_1 _12402_ (.B(_04596_),
    .C(_04598_),
    .A(_04592_),
    .Y(_04599_));
 sg13g2_nand2_1 _12403_ (.Y(_04600_),
    .A(net2441),
    .B(_04599_));
 sg13g2_or2_1 _12404_ (.X(_04601_),
    .B(_04600_),
    .A(_04578_));
 sg13g2_a221oi_1 _12405_ (.B2(_02813_),
    .C1(_04600_),
    .B1(_04577_),
    .A1(net2317),
    .Y(_04602_),
    .A2(_04573_));
 sg13g2_nand2_2 _12406_ (.Y(_04603_),
    .A(_02814_),
    .B(_02824_));
 sg13g2_a21oi_1 _12407_ (.A1(_02814_),
    .A2(_02824_),
    .Y(_04604_),
    .B1(net2444));
 sg13g2_and3_2 _12408_ (.X(_04605_),
    .A(_04576_),
    .B(_04602_),
    .C(_04604_));
 sg13g2_mux4_1 _12409_ (.S0(net2288),
    .A0(\i_tinyqv.cpu.instr_data[1][14] ),
    .A1(\i_tinyqv.cpu.instr_data[0][14] ),
    .A2(\i_tinyqv.cpu.instr_data[3][14] ),
    .A3(\i_tinyqv.cpu.instr_data[2][14] ),
    .S1(net2239),
    .X(_04606_));
 sg13g2_inv_2 _12410_ (.Y(_04607_),
    .A(net2169));
 sg13g2_mux4_1 _12411_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][13] ),
    .A1(\i_tinyqv.cpu.instr_data[0][13] ),
    .A2(\i_tinyqv.cpu.instr_data[3][13] ),
    .A3(\i_tinyqv.cpu.instr_data[2][13] ),
    .S1(net2239),
    .X(_04608_));
 sg13g2_nor2_2 _12412_ (.A(net2169),
    .B(net2167),
    .Y(_04609_));
 sg13g2_or2_1 _12413_ (.X(_04610_),
    .B(net2167),
    .A(net2169));
 sg13g2_mux4_1 _12414_ (.S0(net2288),
    .A0(\i_tinyqv.cpu.instr_data[1][15] ),
    .A1(\i_tinyqv.cpu.instr_data[0][15] ),
    .A2(\i_tinyqv.cpu.instr_data[3][15] ),
    .A3(\i_tinyqv.cpu.instr_data[2][15] ),
    .S1(net2239),
    .X(_04611_));
 sg13g2_inv_2 _12415_ (.Y(_04612_),
    .A(_04611_));
 sg13g2_nor2_2 _12416_ (.A(_04586_),
    .B(_04612_),
    .Y(_04613_));
 sg13g2_and2_1 _12417_ (.A(net2171),
    .B(_04613_),
    .X(_04614_));
 sg13g2_nand2_2 _12418_ (.Y(_04615_),
    .A(net2171),
    .B(_04613_));
 sg13g2_nor2_2 _12419_ (.A(_04610_),
    .B(_04615_),
    .Y(_04616_));
 sg13g2_nand2_1 _12420_ (.Y(_04617_),
    .A(_04609_),
    .B(_04614_));
 sg13g2_mux4_1 _12421_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][5] ),
    .A1(\i_tinyqv.cpu.instr_data[0][5] ),
    .A2(\i_tinyqv.cpu.instr_data[3][5] ),
    .A3(\i_tinyqv.cpu.instr_data[2][5] ),
    .S1(net2235),
    .X(_04618_));
 sg13g2_inv_2 _12422_ (.Y(_04619_),
    .A(net2166));
 sg13g2_mux4_1 _12423_ (.S0(net2289),
    .A0(\i_tinyqv.cpu.instr_data[0][3] ),
    .A1(\i_tinyqv.cpu.instr_data[1][3] ),
    .A2(\i_tinyqv.cpu.instr_data[2][3] ),
    .A3(\i_tinyqv.cpu.instr_data[3][3] ),
    .S1(net2238),
    .X(_04620_));
 sg13g2_mux4_1 _12424_ (.S0(net2289),
    .A0(\i_tinyqv.cpu.instr_data[0][2] ),
    .A1(\i_tinyqv.cpu.instr_data[1][2] ),
    .A2(\i_tinyqv.cpu.instr_data[2][2] ),
    .A3(\i_tinyqv.cpu.instr_data[3][2] ),
    .S1(net2238),
    .X(_04621_));
 sg13g2_nor2_1 _12425_ (.A(net2165),
    .B(net2164),
    .Y(_04622_));
 sg13g2_mux4_1 _12426_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][4] ),
    .A1(\i_tinyqv.cpu.instr_data[0][4] ),
    .A2(\i_tinyqv.cpu.instr_data[3][4] ),
    .A3(\i_tinyqv.cpu.instr_data[2][4] ),
    .S1(net2236),
    .X(_04623_));
 sg13g2_nor3_1 _12427_ (.A(net2165),
    .B(net2164),
    .C(net2163),
    .Y(_04624_));
 sg13g2_inv_1 _12428_ (.Y(_04625_),
    .A(_04624_));
 sg13g2_mux4_1 _12429_ (.S0(net2288),
    .A0(\i_tinyqv.cpu.instr_data[1][6] ),
    .A1(\i_tinyqv.cpu.instr_data[0][6] ),
    .A2(\i_tinyqv.cpu.instr_data[3][6] ),
    .A3(\i_tinyqv.cpu.instr_data[2][6] ),
    .S1(net2236),
    .X(_04626_));
 sg13g2_inv_4 _12430_ (.A(net2161),
    .Y(_04627_));
 sg13g2_nor2_1 _12431_ (.A(_04625_),
    .B(net2161),
    .Y(_04628_));
 sg13g2_nand2_1 _12432_ (.Y(_04629_),
    .A(_04619_),
    .B(_04627_));
 sg13g2_nor2_2 _12433_ (.A(_04625_),
    .B(_04629_),
    .Y(_04630_));
 sg13g2_nand2_2 _12434_ (.Y(_04631_),
    .A(_04616_),
    .B(_04630_));
 sg13g2_mux4_1 _12435_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][10] ),
    .A1(\i_tinyqv.cpu.instr_data[0][10] ),
    .A2(\i_tinyqv.cpu.instr_data[3][10] ),
    .A3(\i_tinyqv.cpu.instr_data[2][10] ),
    .S1(net2237),
    .X(_04632_));
 sg13g2_mux4_1 _12436_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][9] ),
    .A1(\i_tinyqv.cpu.instr_data[0][9] ),
    .A2(\i_tinyqv.cpu.instr_data[3][9] ),
    .A3(\i_tinyqv.cpu.instr_data[2][9] ),
    .S1(net2237),
    .X(_04633_));
 sg13g2_or2_1 _12437_ (.X(_04634_),
    .B(_04633_),
    .A(net2159));
 sg13g2_mux4_1 _12438_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][8] ),
    .A1(\i_tinyqv.cpu.instr_data[0][8] ),
    .A2(\i_tinyqv.cpu.instr_data[3][8] ),
    .A3(\i_tinyqv.cpu.instr_data[2][8] ),
    .S1(net2236),
    .X(_04635_));
 sg13g2_inv_1 _12439_ (.Y(_04636_),
    .A(_04635_));
 sg13g2_nand2b_1 _12440_ (.Y(_04637_),
    .B(_04636_),
    .A_N(_04634_));
 sg13g2_nand2_1 _12441_ (.Y(_04638_),
    .A(\i_tinyqv.cpu.instr_data[0][12] ),
    .B(_04583_));
 sg13g2_a21oi_1 _12442_ (.A1(\i_tinyqv.cpu.instr_data[2][12] ),
    .A2(net2238),
    .Y(_04639_),
    .B1(net2289));
 sg13g2_a21o_1 _12443_ (.A2(net2238),
    .A1(\i_tinyqv.cpu.instr_data[3][12] ),
    .B1(net2288),
    .X(_04640_));
 sg13g2_a21oi_1 _12444_ (.A1(\i_tinyqv.cpu.instr_data[1][12] ),
    .A2(_04583_),
    .Y(_04641_),
    .B1(_04640_));
 sg13g2_a21o_2 _12445_ (.A2(_04639_),
    .A1(_04638_),
    .B1(_04641_),
    .X(_04642_));
 sg13g2_a21oi_2 _12446_ (.B1(_04641_),
    .Y(_04643_),
    .A2(_04639_),
    .A1(_04638_));
 sg13g2_mux4_1 _12447_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][7] ),
    .A1(\i_tinyqv.cpu.instr_data[0][7] ),
    .A2(\i_tinyqv.cpu.instr_data[3][7] ),
    .A3(\i_tinyqv.cpu.instr_data[2][7] ),
    .S1(net2235),
    .X(_04644_));
 sg13g2_inv_1 _12448_ (.Y(_04645_),
    .A(_04644_));
 sg13g2_nor4_2 _12449_ (.A(_04631_),
    .B(_04637_),
    .C(net2055),
    .Y(_04646_),
    .D(_04645_));
 sg13g2_and4_1 _12450_ (.A(_04576_),
    .B(_04602_),
    .C(_04604_),
    .D(_04646_),
    .X(_04647_));
 sg13g2_nand2_2 _12451_ (.Y(_04648_),
    .A(_04605_),
    .B(_04646_));
 sg13g2_nor2_2 _12452_ (.A(net1883),
    .B(net1870),
    .Y(_04649_));
 sg13g2_or2_1 _12453_ (.X(_04650_),
    .B(net1868),
    .A(net1879));
 sg13g2_nand2_2 _12454_ (.Y(_04651_),
    .A(net2496),
    .B(_04649_));
 sg13g2_nor2_1 _12455_ (.A(_04568_),
    .B(_04651_),
    .Y(_04652_));
 sg13g2_nor3_1 _12456_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_04568_),
    .C(_04651_),
    .Y(_04653_));
 sg13g2_and2_1 _12457_ (.A(\i_tinyqv.cpu.instr_write_offset[1] ),
    .B(_04653_),
    .X(_04654_));
 sg13g2_mux2_1 _12458_ (.A0(net4562),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net1812),
    .X(_00461_));
 sg13g2_nor2_1 _12459_ (.A(net4269),
    .B(net1812),
    .Y(_04655_));
 sg13g2_a21oi_1 _12460_ (.A1(_02037_),
    .A2(net1812),
    .Y(_00462_),
    .B1(_04655_));
 sg13g2_mux2_1 _12461_ (.A0(net4434),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(net1813),
    .X(_00463_));
 sg13g2_mux2_1 _12462_ (.A0(net4464),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(net1811),
    .X(_00464_));
 sg13g2_mux2_1 _12463_ (.A0(net4614),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net1813),
    .X(_00465_));
 sg13g2_mux2_1 _12464_ (.A0(net4418),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(net1811),
    .X(_00466_));
 sg13g2_nor2_1 _12465_ (.A(net4163),
    .B(net1811),
    .Y(_04656_));
 sg13g2_a21oi_1 _12466_ (.A1(net2410),
    .A2(net1811),
    .Y(_00467_),
    .B1(_04656_));
 sg13g2_mux2_1 _12467_ (.A0(net4594),
    .A1(net2602),
    .S(net1811),
    .X(_00468_));
 sg13g2_mux2_1 _12468_ (.A0(net4484),
    .A1(net2600),
    .S(net1811),
    .X(_00469_));
 sg13g2_mux2_1 _12469_ (.A0(net4592),
    .A1(net2598),
    .S(net1811),
    .X(_00470_));
 sg13g2_mux2_1 _12470_ (.A0(net4521),
    .A1(net2596),
    .S(net1812),
    .X(_00471_));
 sg13g2_mux2_1 _12471_ (.A0(net4475),
    .A1(net2594),
    .S(net1811),
    .X(_00472_));
 sg13g2_mux2_1 _12472_ (.A0(net4516),
    .A1(net2592),
    .S(net1812),
    .X(_00473_));
 sg13g2_mux2_1 _12473_ (.A0(net4482),
    .A1(net2590),
    .S(net1813),
    .X(_00474_));
 sg13g2_nor2_1 _12474_ (.A(net3412),
    .B(_04338_),
    .Y(_00475_));
 sg13g2_o21ai_1 _12475_ (.B1(net2672),
    .Y(_04657_),
    .A1(net3412),
    .A2(net3575));
 sg13g2_a21oi_1 _12476_ (.A1(net3412),
    .A2(net3575),
    .Y(_00476_),
    .B1(_04657_));
 sg13g2_and3_1 _12477_ (.X(_04658_),
    .A(net3412),
    .B(net3575),
    .C(net3704));
 sg13g2_a21oi_1 _12478_ (.A1(net3412),
    .A2(net3575),
    .Y(_04659_),
    .B1(net3704));
 sg13g2_nor3_1 _12479_ (.A(_04338_),
    .B(_04658_),
    .C(_04659_),
    .Y(_00477_));
 sg13g2_and2_1 _12480_ (.A(net4129),
    .B(_04658_),
    .X(_04660_));
 sg13g2_nor2_1 _12481_ (.A(net4129),
    .B(_04658_),
    .Y(_04661_));
 sg13g2_nor3_1 _12482_ (.A(_04338_),
    .B(_04660_),
    .C(_04661_),
    .Y(_00478_));
 sg13g2_a21oi_1 _12483_ (.A1(net4845),
    .A2(_04660_),
    .Y(_04662_),
    .B1(_04338_));
 sg13g2_o21ai_1 _12484_ (.B1(_04662_),
    .Y(_04663_),
    .A1(net4845),
    .A2(_04660_));
 sg13g2_inv_1 _12485_ (.Y(_00479_),
    .A(_04663_));
 sg13g2_and2_1 _12486_ (.A(_02089_),
    .B(net2390),
    .X(_04664_));
 sg13g2_a21oi_2 _12487_ (.B1(net2388),
    .Y(_04665_),
    .A2(\i_tinyqv.cpu.data_read_n[0] ),
    .A1(\i_tinyqv.cpu.data_read_n[1] ));
 sg13g2_or2_1 _12488_ (.X(_04666_),
    .B(_04665_),
    .A(_04664_));
 sg13g2_nor2_1 _12489_ (.A(net2612),
    .B(net2613),
    .Y(_04667_));
 sg13g2_nand2_1 _12490_ (.Y(_04668_),
    .A(_04666_),
    .B(_04667_));
 sg13g2_o21ai_1 _12491_ (.B1(\i_tinyqv.mem.data_stall ),
    .Y(_04669_),
    .A1(_03132_),
    .A2(_04668_));
 sg13g2_xnor2_1 _12492_ (.Y(_04670_),
    .A(net2613),
    .B(_02758_));
 sg13g2_xor2_1 _12493_ (.B(net2613),
    .A(net2612),
    .X(_04671_));
 sg13g2_o21ai_1 _12494_ (.B1(\i_tinyqv.mem.q_ctrl.data_req ),
    .Y(_04672_),
    .A1(_02757_),
    .A2(_04671_));
 sg13g2_a21oi_1 _12495_ (.A1(_02757_),
    .A2(_04671_),
    .Y(_04673_),
    .B1(_04672_));
 sg13g2_a22oi_1 _12496_ (.Y(_04674_),
    .B1(_04670_),
    .B2(_04673_),
    .A2(_02763_),
    .A1(\i_tinyqv.mem.q_ctrl.data_ready ));
 sg13g2_a21oi_1 _12497_ (.A1(_04669_),
    .A2(_04674_),
    .Y(_00480_),
    .B1(_02018_));
 sg13g2_o21ai_1 _12498_ (.B1(_03116_),
    .Y(_04675_),
    .A1(_03113_),
    .A2(_03118_));
 sg13g2_nand2_1 _12499_ (.Y(_04676_),
    .A(net2576),
    .B(net2126));
 sg13g2_nand2_2 _12500_ (.Y(_04677_),
    .A(net2577),
    .B(net2135));
 sg13g2_or2_1 _12501_ (.X(_04678_),
    .B(_04677_),
    .A(_03114_));
 sg13g2_xor2_1 _12502_ (.B(_04677_),
    .A(_03114_),
    .X(_04679_));
 sg13g2_nand2b_1 _12503_ (.Y(_04680_),
    .B(_04679_),
    .A_N(_04676_));
 sg13g2_xnor2_1 _12504_ (.Y(_04681_),
    .A(_04676_),
    .B(_04679_));
 sg13g2_nand2_1 _12505_ (.Y(_04682_),
    .A(_04675_),
    .B(_04681_));
 sg13g2_xnor2_1 _12506_ (.Y(_04683_),
    .A(_04675_),
    .B(_04681_));
 sg13g2_o21ai_1 _12507_ (.B1(_03120_),
    .Y(_04684_),
    .A1(_03111_),
    .A2(_03121_));
 sg13g2_nand2b_1 _12508_ (.Y(_04685_),
    .B(_04684_),
    .A_N(_04683_));
 sg13g2_xor2_1 _12509_ (.B(_04684_),
    .A(_04683_),
    .X(_04686_));
 sg13g2_o21ai_1 _12510_ (.B1(_03123_),
    .Y(_04687_),
    .A1(_02060_),
    .A2(_03124_));
 sg13g2_nand2b_1 _12511_ (.Y(_04688_),
    .B(_04687_),
    .A_N(_04686_));
 sg13g2_xnor2_1 _12512_ (.Y(_04689_),
    .A(_04686_),
    .B(_04687_));
 sg13g2_o21ai_1 _12513_ (.B1(_04689_),
    .Y(_04690_),
    .A1(_03127_),
    .A2(_03129_));
 sg13g2_or3_1 _12514_ (.A(_03127_),
    .B(_03129_),
    .C(_04689_),
    .X(_04691_));
 sg13g2_and2_1 _12515_ (.A(_04690_),
    .B(_04691_),
    .X(_00481_));
 sg13g2_nand2_1 _12516_ (.Y(_04692_),
    .A(_04688_),
    .B(_04690_));
 sg13g2_nand2_1 _12517_ (.Y(_04693_),
    .A(net2576),
    .B(net2129));
 sg13g2_nor2_1 _12518_ (.A(_04677_),
    .B(_04693_),
    .Y(_04694_));
 sg13g2_a22oi_1 _12519_ (.Y(_04695_),
    .B1(net2129),
    .B2(net2577),
    .A2(net2135),
    .A1(net2576));
 sg13g2_or2_1 _12520_ (.X(_04696_),
    .B(_04695_),
    .A(_04694_));
 sg13g2_a21oi_1 _12521_ (.A1(_04678_),
    .A2(_04680_),
    .Y(_04697_),
    .B1(_04696_));
 sg13g2_nand3_1 _12522_ (.B(_04680_),
    .C(_04696_),
    .A(_04678_),
    .Y(_04698_));
 sg13g2_nand2b_1 _12523_ (.Y(_04699_),
    .B(_04698_),
    .A_N(_04697_));
 sg13g2_nor2_1 _12524_ (.A(_04685_),
    .B(_04699_),
    .Y(_04700_));
 sg13g2_nor2_1 _12525_ (.A(_04682_),
    .B(_04699_),
    .Y(_04701_));
 sg13g2_and2_1 _12526_ (.A(_04682_),
    .B(_04699_),
    .X(_04702_));
 sg13g2_o21ai_1 _12527_ (.B1(_04685_),
    .Y(_04703_),
    .A1(_04701_),
    .A2(_04702_));
 sg13g2_nand2b_1 _12528_ (.Y(_04704_),
    .B(_04703_),
    .A_N(_04700_));
 sg13g2_xnor2_1 _12529_ (.Y(_00482_),
    .A(_04692_),
    .B(_04704_));
 sg13g2_nand2b_1 _12530_ (.Y(_04705_),
    .B(_04677_),
    .A_N(_04693_));
 sg13g2_nor2_1 _12531_ (.A(_04697_),
    .B(_04701_),
    .Y(_04706_));
 sg13g2_xor2_1 _12532_ (.B(_04706_),
    .A(_04705_),
    .X(_04707_));
 sg13g2_a21o_1 _12533_ (.A2(_04703_),
    .A1(_04692_),
    .B1(_04700_),
    .X(_04708_));
 sg13g2_xor2_1 _12534_ (.B(_04708_),
    .A(_04707_),
    .X(_00483_));
 sg13g2_a21oi_1 _12535_ (.A1(_04677_),
    .A2(_04706_),
    .Y(_04709_),
    .B1(_04693_));
 sg13g2_a21o_1 _12536_ (.A2(_04708_),
    .A1(_04707_),
    .B1(_04709_),
    .X(_00484_));
 sg13g2_nor2_1 _12537_ (.A(net5292),
    .B(net4873),
    .Y(_04710_));
 sg13g2_nor2b_2 _12538_ (.A(net2169),
    .B_N(net2167),
    .Y(_04711_));
 sg13g2_nand2_1 _12539_ (.Y(_04712_),
    .A(_04607_),
    .B(net2167));
 sg13g2_nor2b_2 _12540_ (.A(net2171),
    .B_N(_04586_),
    .Y(_04713_));
 sg13g2_and2_1 _12541_ (.A(_04711_),
    .B(_04713_),
    .X(_04714_));
 sg13g2_nand2_2 _12542_ (.Y(_04715_),
    .A(_04711_),
    .B(_04713_));
 sg13g2_nand2_1 _12543_ (.Y(_04716_),
    .A(net2166),
    .B(net2161));
 sg13g2_nor2_1 _12544_ (.A(net2163),
    .B(_04716_),
    .Y(_04717_));
 sg13g2_and2_1 _12545_ (.A(_04621_),
    .B(_04717_),
    .X(_04718_));
 sg13g2_nand2_2 _12546_ (.Y(_04719_),
    .A(net2165),
    .B(_04718_));
 sg13g2_o21ai_1 _12547_ (.B1(_04715_),
    .Y(_04720_),
    .A1(net2105),
    .A2(_04719_));
 sg13g2_and4_1 _12548_ (.A(_04576_),
    .B(_04602_),
    .C(_04604_),
    .D(_04720_),
    .X(_04721_));
 sg13g2_nand2_1 _12549_ (.Y(_04722_),
    .A(_04605_),
    .B(_04720_));
 sg13g2_a21o_1 _12550_ (.A2(net1882),
    .A1(net2441),
    .B1(net5111),
    .X(_04723_));
 sg13g2_a221oi_1 _12551_ (.B2(_04720_),
    .C1(net1869),
    .B1(_04605_),
    .A1(net2441),
    .Y(_04724_),
    .A2(net1881));
 sg13g2_nor3_1 _12552_ (.A(net1870),
    .B(_04721_),
    .C(_04723_),
    .Y(_04725_));
 sg13g2_nor4_2 _12553_ (.A(net1870),
    .B(_04664_),
    .C(_04721_),
    .Y(_04726_),
    .D(_04723_));
 sg13g2_nor2_1 _12554_ (.A(net2606),
    .B(net2608),
    .Y(_04727_));
 sg13g2_nor3_2 _12555_ (.A(net2604),
    .B(net2606),
    .C(net2607),
    .Y(_04728_));
 sg13g2_nand2b_2 _12556_ (.Y(_04729_),
    .B(_04727_),
    .A_N(net2604));
 sg13g2_nor2_1 _12557_ (.A(net4033),
    .B(_04729_),
    .Y(_04730_));
 sg13g2_nor3_2 _12558_ (.A(net4033),
    .B(_04665_),
    .C(_04729_),
    .Y(_04731_));
 sg13g2_a21oi_1 _12559_ (.A1(_04726_),
    .A2(_04731_),
    .Y(_04732_),
    .B1(net2611));
 sg13g2_a21o_2 _12560_ (.A2(_04731_),
    .A1(_04726_),
    .B1(\i_tinyqv.mem.instr_active ),
    .X(_04733_));
 sg13g2_nand2b_1 _12561_ (.Y(_04734_),
    .B(net1855),
    .A_N(_04565_));
 sg13g2_a21oi_1 _12562_ (.A1(_02762_),
    .A2(net1859),
    .Y(_04735_),
    .B1(_02760_));
 sg13g2_a21oi_1 _12563_ (.A1(_04734_),
    .A2(_04735_),
    .Y(_04736_),
    .B1(_04710_));
 sg13g2_o21ai_1 _12564_ (.B1(_04730_),
    .Y(_04737_),
    .A1(_04665_),
    .A2(_04726_));
 sg13g2_nand2_1 _12565_ (.Y(_04738_),
    .A(_04664_),
    .B(_04731_));
 sg13g2_and2_1 _12566_ (.A(_04737_),
    .B(_04738_),
    .X(_04739_));
 sg13g2_nand2_1 _12567_ (.Y(_04740_),
    .A(_04737_),
    .B(_04738_));
 sg13g2_nand2_1 _12568_ (.Y(_04741_),
    .A(net2630),
    .B(net1835));
 sg13g2_o21ai_1 _12569_ (.B1(net2613),
    .Y(_04742_),
    .A1(net5292),
    .A2(net4873));
 sg13g2_o21ai_1 _12570_ (.B1(_04742_),
    .Y(_04743_),
    .A1(net2613),
    .A2(_04736_));
 sg13g2_nor2_1 _12571_ (.A(_04741_),
    .B(_04743_),
    .Y(_00485_));
 sg13g2_a22oi_1 _12572_ (.Y(_04744_),
    .B1(_04736_),
    .B2(_04671_),
    .A2(_04710_),
    .A1(net2612));
 sg13g2_nor2_1 _12573_ (.A(_04741_),
    .B(_04744_),
    .Y(_00486_));
 sg13g2_nand2_2 _12574_ (.Y(_04745_),
    .A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .B(_04667_));
 sg13g2_nor2_1 _12575_ (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .B(_04745_),
    .Y(_04746_));
 sg13g2_a21oi_1 _12576_ (.A1(_02035_),
    .A2(_04745_),
    .Y(_00487_),
    .B1(_04746_));
 sg13g2_nor2_1 _12577_ (.A(net2602),
    .B(net2286),
    .Y(_04747_));
 sg13g2_a21oi_1 _12578_ (.A1(_02036_),
    .A2(net2286),
    .Y(_00488_),
    .B1(_04747_));
 sg13g2_mux2_1 _12579_ (.A0(net2600),
    .A1(net5074),
    .S(net2286),
    .X(_00489_));
 sg13g2_nor2_1 _12580_ (.A(net2598),
    .B(net2286),
    .Y(_04748_));
 sg13g2_a21oi_1 _12581_ (.A1(_02037_),
    .A2(net2286),
    .Y(_00490_),
    .B1(_04748_));
 sg13g2_mux2_1 _12582_ (.A0(net2596),
    .A1(net5008),
    .S(net2286),
    .X(_00491_));
 sg13g2_mux2_1 _12583_ (.A0(net2594),
    .A1(net5097),
    .S(net2286),
    .X(_00492_));
 sg13g2_mux2_1 _12584_ (.A0(net2592),
    .A1(net5016),
    .S(net2286),
    .X(_00493_));
 sg13g2_mux2_1 _12585_ (.A0(net2590),
    .A1(net5254),
    .S(_04745_),
    .X(_00494_));
 sg13g2_nand2_1 _12586_ (.Y(_04749_),
    .A(\i_tinyqv.cpu.instr_data_in[8] ),
    .B(net2299));
 sg13g2_o21ai_1 _12587_ (.B1(_04749_),
    .Y(_00495_),
    .A1(_02063_),
    .A2(net2299));
 sg13g2_nand2_1 _12588_ (.Y(_04750_),
    .A(net2602),
    .B(net2299));
 sg13g2_o21ai_1 _12589_ (.B1(_04750_),
    .Y(_00496_),
    .A1(_02071_),
    .A2(net2299));
 sg13g2_nand2_1 _12590_ (.Y(_04751_),
    .A(net2601),
    .B(net2300));
 sg13g2_o21ai_1 _12591_ (.B1(_04751_),
    .Y(_00497_),
    .A1(_02077_),
    .A2(net2300));
 sg13g2_nand2_1 _12592_ (.Y(_04752_),
    .A(net2599),
    .B(net2299));
 sg13g2_o21ai_1 _12593_ (.B1(_04752_),
    .Y(_00498_),
    .A1(_02082_),
    .A2(net2299));
 sg13g2_nand2_1 _12594_ (.Y(_04753_),
    .A(net2597),
    .B(net2301));
 sg13g2_o21ai_1 _12595_ (.B1(_04753_),
    .Y(_00499_),
    .A1(_02064_),
    .A2(net2300));
 sg13g2_nand2_1 _12596_ (.Y(_04754_),
    .A(net2595),
    .B(net2301));
 sg13g2_o21ai_1 _12597_ (.B1(_04754_),
    .Y(_00500_),
    .A1(_02072_),
    .A2(net2300));
 sg13g2_nand2_1 _12598_ (.Y(_04755_),
    .A(net2593),
    .B(net2301));
 sg13g2_o21ai_1 _12599_ (.B1(_04755_),
    .Y(_00501_),
    .A1(_02078_),
    .A2(net2301));
 sg13g2_nand2_1 _12600_ (.Y(_04756_),
    .A(net2591),
    .B(net2300));
 sg13g2_o21ai_1 _12601_ (.B1(_04756_),
    .Y(_00502_),
    .A1(_02083_),
    .A2(net2300));
 sg13g2_nor3_2 _12602_ (.A(_01983_),
    .B(net2614),
    .C(_02003_),
    .Y(_04757_));
 sg13g2_nor2_1 _12603_ (.A(net3793),
    .B(net2285),
    .Y(_04758_));
 sg13g2_a21oi_1 _12604_ (.A1(net2410),
    .A2(net2285),
    .Y(_00503_),
    .B1(net3794));
 sg13g2_mux2_1 _12605_ (.A0(net4175),
    .A1(net2603),
    .S(net2285),
    .X(_00504_));
 sg13g2_mux2_1 _12606_ (.A0(net4263),
    .A1(net2601),
    .S(net2285),
    .X(_00505_));
 sg13g2_mux2_1 _12607_ (.A0(net4239),
    .A1(net2599),
    .S(net2285),
    .X(_00506_));
 sg13g2_mux2_1 _12608_ (.A0(net4096),
    .A1(net2597),
    .S(net2285),
    .X(_00507_));
 sg13g2_mux2_1 _12609_ (.A0(net4167),
    .A1(net2595),
    .S(net2285),
    .X(_00508_));
 sg13g2_mux2_1 _12610_ (.A0(net4195),
    .A1(net2593),
    .S(net2285),
    .X(_00509_));
 sg13g2_mux2_1 _12611_ (.A0(net4372),
    .A1(net2591),
    .S(_04757_),
    .X(_00510_));
 sg13g2_nand3_1 _12612_ (.B(net2614),
    .C(\i_tinyqv.mem.q_ctrl.data_ready ),
    .A(net2612),
    .Y(_04759_));
 sg13g2_nand2_1 _12613_ (.Y(_04760_),
    .A(net3486),
    .B(net2337));
 sg13g2_o21ai_1 _12614_ (.B1(_04760_),
    .Y(_00511_),
    .A1(net2410),
    .A2(net2337));
 sg13g2_mux2_1 _12615_ (.A0(net2603),
    .A1(net4158),
    .S(net2337),
    .X(_00512_));
 sg13g2_mux2_1 _12616_ (.A0(net2601),
    .A1(net4145),
    .S(net2337),
    .X(_00513_));
 sg13g2_mux2_1 _12617_ (.A0(net2599),
    .A1(net4100),
    .S(net2337),
    .X(_00514_));
 sg13g2_mux2_1 _12618_ (.A0(net2597),
    .A1(net4088),
    .S(net2337),
    .X(_00515_));
 sg13g2_mux2_1 _12619_ (.A0(net2595),
    .A1(net4153),
    .S(net2337),
    .X(_00516_));
 sg13g2_mux2_1 _12620_ (.A0(net2593),
    .A1(net4130),
    .S(_04759_),
    .X(_00517_));
 sg13g2_nor2_1 _12621_ (.A(net2591),
    .B(_04759_),
    .Y(_04761_));
 sg13g2_a21oi_1 _12622_ (.A1(_02085_),
    .A2(net2337),
    .Y(_00518_),
    .B1(_04761_));
 sg13g2_and3_1 _12623_ (.X(_00519_),
    .A(net2630),
    .B(_04726_),
    .C(net4034));
 sg13g2_nand3_1 _12624_ (.B(_02823_),
    .C(_03348_),
    .A(_02814_),
    .Y(_04762_));
 sg13g2_and3_2 _12625_ (.X(_04763_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(\i_tinyqv.cpu.instr_write_offset[1] ),
    .C(_04567_));
 sg13g2_xor2_1 _12626_ (.B(_04763_),
    .A(net5375),
    .X(_04764_));
 sg13g2_xnor2_1 _12627_ (.Y(_04765_),
    .A(_04762_),
    .B(_04764_));
 sg13g2_a21oi_1 _12628_ (.A1(net5355),
    .A2(_04567_),
    .Y(_04766_),
    .B1(net5369));
 sg13g2_or2_1 _12629_ (.X(_04767_),
    .B(_04766_),
    .A(_04763_));
 sg13g2_xnor2_1 _12630_ (.Y(_04768_),
    .A(net5355),
    .B(_04567_));
 sg13g2_xor2_1 _12631_ (.B(_04768_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .X(_04769_));
 sg13g2_xor2_1 _12632_ (.B(_04767_),
    .A(\i_tinyqv.cpu.pc[2] ),
    .X(_04770_));
 sg13g2_and3_2 _12633_ (.X(_04771_),
    .A(_04765_),
    .B(_04769_),
    .C(_04770_));
 sg13g2_nand4_1 _12634_ (.B(_02003_),
    .C(_04565_),
    .A(net2611),
    .Y(_04772_),
    .D(_04771_));
 sg13g2_nand2_1 _12635_ (.Y(_04773_),
    .A(net5269),
    .B(_04772_));
 sg13g2_o21ai_1 _12636_ (.B1(_04666_),
    .Y(_04774_),
    .A1(net2300),
    .A2(_04771_));
 sg13g2_nand2_1 _12637_ (.Y(_04775_),
    .A(net2611),
    .B(_04774_));
 sg13g2_a21oi_1 _12638_ (.A1(_04725_),
    .A2(_04773_),
    .Y(_04776_),
    .B1(_04775_));
 sg13g2_nor2_1 _12639_ (.A(net3652),
    .B(_04710_),
    .Y(_04777_));
 sg13g2_a21oi_1 _12640_ (.A1(_02763_),
    .A2(_04777_),
    .Y(_04778_),
    .B1(net2611));
 sg13g2_nor3_1 _12641_ (.A(_04730_),
    .B(_04776_),
    .C(_04778_),
    .Y(_04779_));
 sg13g2_a22oi_1 _12642_ (.Y(_04780_),
    .B1(_04731_),
    .B2(_04726_),
    .A2(_04729_),
    .A1(net4859));
 sg13g2_nor3_1 _12643_ (.A(net2431),
    .B(_04779_),
    .C(net4860),
    .Y(_00520_));
 sg13g2_nand2_1 _12644_ (.Y(_04781_),
    .A(net2624),
    .B(net4019));
 sg13g2_o21ai_1 _12645_ (.B1(_04781_),
    .Y(_00521_),
    .A1(net2624),
    .A2(_02042_));
 sg13g2_nor2_1 _12646_ (.A(net2623),
    .B(net11),
    .Y(_04782_));
 sg13g2_a21oi_1 _12647_ (.A1(net2623),
    .A2(_02039_),
    .Y(_00522_),
    .B1(_04782_));
 sg13g2_o21ai_1 _12648_ (.B1(_04779_),
    .Y(_04783_),
    .A1(net2439),
    .A2(net4625));
 sg13g2_nand3b_1 _12649_ (.B(_04783_),
    .C(net2630),
    .Y(_04784_),
    .A_N(net5033));
 sg13g2_nor2_1 _12650_ (.A(_04728_),
    .B(net1794),
    .Y(_04785_));
 sg13g2_nand2b_2 _12651_ (.Y(_04786_),
    .B(_04772_),
    .A_N(\i_tinyqv.mem.data_stall ));
 sg13g2_nor2_1 _12652_ (.A(net4910),
    .B(_04786_),
    .Y(_04787_));
 sg13g2_inv_1 _12653_ (.Y(_04788_),
    .A(_04787_));
 sg13g2_nand2_2 _12654_ (.Y(_04789_),
    .A(net2605),
    .B(net5327));
 sg13g2_nor2_2 _12655_ (.A(net2607),
    .B(_04789_),
    .Y(_04790_));
 sg13g2_or2_1 _12656_ (.X(_04791_),
    .B(_04789_),
    .A(net2607));
 sg13g2_nor3_2 _12657_ (.A(net4281),
    .B(net4380),
    .C(net4960),
    .Y(_04792_));
 sg13g2_or3_1 _12658_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .B(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .C(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .X(_04793_));
 sg13g2_nand2_1 _12659_ (.Y(_04794_),
    .A(_04791_),
    .B(_04792_));
 sg13g2_nand3_1 _12660_ (.B(net2606),
    .C(net2607),
    .A(net2605),
    .Y(_04795_));
 sg13g2_nand2_2 _12661_ (.Y(_04796_),
    .A(net2605),
    .B(net2607));
 sg13g2_a21oi_1 _12662_ (.A1(net2609),
    .A2(_04795_),
    .Y(_04797_),
    .B1(_04796_));
 sg13g2_nor2_1 _12663_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .Y(_04798_));
 sg13g2_nand2_1 _12664_ (.Y(_04799_),
    .A(_04797_),
    .B(_04798_));
 sg13g2_o21ai_1 _12665_ (.B1(_04799_),
    .Y(_04800_),
    .A1(_01982_),
    .A2(_04797_));
 sg13g2_nor2b_2 _12666_ (.A(_04794_),
    .B_N(_04800_),
    .Y(_04801_));
 sg13g2_and2_1 _12667_ (.A(net2605),
    .B(_04727_),
    .X(_04802_));
 sg13g2_o21ai_1 _12668_ (.B1(_04796_),
    .Y(_04803_),
    .A1(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .A2(_04802_));
 sg13g2_a21oi_1 _12669_ (.A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .A2(_04802_),
    .Y(_04804_),
    .B1(_04803_));
 sg13g2_a221oi_1 _12670_ (.B2(_04804_),
    .C1(net5035),
    .B1(_04801_),
    .A1(_04787_),
    .Y(_04805_),
    .A2(_04790_));
 sg13g2_nor2_1 _12671_ (.A(net2609),
    .B(_04791_),
    .Y(_04806_));
 sg13g2_and2_1 _12672_ (.A(_04787_),
    .B(_04806_),
    .X(_04807_));
 sg13g2_nor2_1 _12673_ (.A(_04786_),
    .B(_04796_),
    .Y(_04808_));
 sg13g2_nor2_1 _12674_ (.A(_04804_),
    .B(_04808_),
    .Y(_04809_));
 sg13g2_a22oi_1 _12675_ (.Y(_04810_),
    .B1(_04809_),
    .B2(_04801_),
    .A2(_04807_),
    .A1(net4019));
 sg13g2_nand2b_1 _12676_ (.Y(_04811_),
    .B(_04810_),
    .A_N(_04805_));
 sg13g2_mux2_1 _12677_ (.A0(net5035),
    .A1(_04811_),
    .S(_04785_),
    .X(_00523_));
 sg13g2_nor2b_1 _12678_ (.A(_04796_),
    .B_N(_04801_),
    .Y(_04812_));
 sg13g2_nand2_1 _12679_ (.Y(_04813_),
    .A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ));
 sg13g2_mux2_1 _12680_ (.A0(_04813_),
    .A1(_02039_),
    .S(_04786_),
    .X(_04814_));
 sg13g2_nor2b_1 _12681_ (.A(_04801_),
    .B_N(_04813_),
    .Y(_04815_));
 sg13g2_o21ai_1 _12682_ (.B1(_04796_),
    .Y(_04816_),
    .A1(_04802_),
    .A2(_04813_));
 sg13g2_a21oi_1 _12683_ (.A1(net4341),
    .A2(_04802_),
    .Y(_04817_),
    .B1(_04816_));
 sg13g2_a221oi_1 _12684_ (.B2(_04801_),
    .C1(_04815_),
    .B1(_04817_),
    .A1(_04812_),
    .Y(_04818_),
    .A2(_04814_));
 sg13g2_mux2_1 _12685_ (.A0(net4910),
    .A1(_04818_),
    .S(_04785_),
    .X(_00524_));
 sg13g2_nand2_1 _12686_ (.Y(_04819_),
    .A(net2609),
    .B(_04037_));
 sg13g2_nor4_1 _12687_ (.A(net1795),
    .B(_04794_),
    .C(_04800_),
    .D(_04819_),
    .Y(_00525_));
 sg13g2_nand2_2 _12688_ (.Y(_04820_),
    .A(_01982_),
    .B(_04791_));
 sg13g2_nand2_1 _12689_ (.Y(_04821_),
    .A(net4684),
    .B(net1858));
 sg13g2_nor2_1 _12690_ (.A(net4599),
    .B(_04821_),
    .Y(_04822_));
 sg13g2_or4_1 _12691_ (.A(_01808_),
    .B(\addr[23] ),
    .C(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .D(net1852),
    .X(_04823_));
 sg13g2_and3_1 _12692_ (.X(_04824_),
    .A(net4684),
    .B(net4599),
    .C(net1858));
 sg13g2_nand4_1 _12693_ (.B(\addr[23] ),
    .C(_02019_),
    .A(\addr[24] ),
    .Y(_04825_),
    .D(net1858));
 sg13g2_nand3_1 _12694_ (.B(_04823_),
    .C(_04825_),
    .A(net1831),
    .Y(_04826_));
 sg13g2_nand2_1 _12695_ (.Y(_04827_),
    .A(_04728_),
    .B(net1810));
 sg13g2_a221oi_1 _12696_ (.B2(_04827_),
    .C1(net1795),
    .B1(_04820_),
    .A1(_01982_),
    .Y(_00526_),
    .A2(_04728_));
 sg13g2_nor2_1 _12697_ (.A(_04728_),
    .B(_04800_),
    .Y(_04828_));
 sg13g2_a22oi_1 _12698_ (.Y(_04829_),
    .B1(_04828_),
    .B2(_04791_),
    .A2(net1810),
    .A1(_04728_));
 sg13g2_nand2_2 _12699_ (.Y(_04830_),
    .A(_04791_),
    .B(_04829_));
 sg13g2_a21oi_1 _12700_ (.A1(net4960),
    .A2(_04729_),
    .Y(_04831_),
    .B1(_04830_));
 sg13g2_a21oi_1 _12701_ (.A1(net4960),
    .A2(_04830_),
    .Y(_04832_),
    .B1(_04831_));
 sg13g2_nor2_1 _12702_ (.A(net1793),
    .B(_04832_),
    .Y(_00527_));
 sg13g2_a21oi_1 _12703_ (.A1(_04791_),
    .A2(_04829_),
    .Y(_04833_),
    .B1(net4380));
 sg13g2_nand2_1 _12704_ (.Y(_04834_),
    .A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .B(net2439));
 sg13g2_nand2b_1 _12705_ (.Y(_04835_),
    .B(_04834_),
    .A_N(net2608));
 sg13g2_nand2_1 _12706_ (.Y(_04836_),
    .A(_04038_),
    .B(_04835_));
 sg13g2_xor2_1 _12707_ (.B(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .A(net4380),
    .X(_04837_));
 sg13g2_a21oi_1 _12708_ (.A1(_04792_),
    .A2(_04836_),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_a21oi_1 _12709_ (.A1(_04729_),
    .A2(_04838_),
    .Y(_04839_),
    .B1(_04830_));
 sg13g2_nor3_1 _12710_ (.A(net1793),
    .B(_04833_),
    .C(_04839_),
    .Y(_00528_));
 sg13g2_a21oi_1 _12711_ (.A1(_04791_),
    .A2(_04829_),
    .Y(_04840_),
    .B1(net4281));
 sg13g2_nand3b_1 _12712_ (.B(_04034_),
    .C(_04792_),
    .Y(_04841_),
    .A_N(net2605));
 sg13g2_o21ai_1 _12713_ (.B1(net4281),
    .Y(_04842_),
    .A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_a21oi_1 _12714_ (.A1(_04841_),
    .A2(_04842_),
    .Y(_04843_),
    .B1(_04728_));
 sg13g2_a21oi_1 _12715_ (.A1(\addr[24] ),
    .A2(net1858),
    .Y(_04844_),
    .B1(_04729_));
 sg13g2_nor3_1 _12716_ (.A(_04830_),
    .B(_04843_),
    .C(_04844_),
    .Y(_04845_));
 sg13g2_nor3_1 _12717_ (.A(net1794),
    .B(_04840_),
    .C(_04845_),
    .Y(_00529_));
 sg13g2_nor2_1 _12718_ (.A(_04821_),
    .B(net1810),
    .Y(_04846_));
 sg13g2_nand2_1 _12719_ (.Y(_04847_),
    .A(_04737_),
    .B(_04846_));
 sg13g2_nand2_1 _12720_ (.Y(_04848_),
    .A(net2609),
    .B(_04826_));
 sg13g2_a21oi_1 _12721_ (.A1(_04847_),
    .A2(_04848_),
    .Y(_00530_),
    .B1(net1795));
 sg13g2_a22oi_1 _12722_ (.Y(_04849_),
    .B1(_04801_),
    .B2(_04808_),
    .A2(_04790_),
    .A1(_04787_));
 sg13g2_nor4_1 _12723_ (.A(net2609),
    .B(_04728_),
    .C(net1795),
    .D(net5328),
    .Y(_00531_));
 sg13g2_nand4_1 _12724_ (.B(_04789_),
    .C(_04793_),
    .A(_04729_),
    .Y(_04850_),
    .D(_04800_));
 sg13g2_nand2_1 _12725_ (.Y(_04851_),
    .A(_04829_),
    .B(_04850_));
 sg13g2_a21oi_1 _12726_ (.A1(_04788_),
    .A2(_04790_),
    .Y(_04852_),
    .B1(_04851_));
 sg13g2_o21ai_1 _12727_ (.B1(_04792_),
    .Y(_04853_),
    .A1(net2608),
    .A2(_04038_));
 sg13g2_nor2_1 _12728_ (.A(_04808_),
    .B(_04853_),
    .Y(_04854_));
 sg13g2_inv_1 _12729_ (.Y(_04855_),
    .A(_04854_));
 sg13g2_a21oi_1 _12730_ (.A1(_04835_),
    .A2(_04854_),
    .Y(_04856_),
    .B1(_04844_));
 sg13g2_a22oi_1 _12731_ (.Y(_04857_),
    .B1(_04852_),
    .B2(_04856_),
    .A2(_04851_),
    .A1(net2608));
 sg13g2_nor2_1 _12732_ (.A(net1793),
    .B(_04857_),
    .Y(_00532_));
 sg13g2_nor3_1 _12733_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .B(net2607),
    .C(net2609),
    .Y(_04858_));
 sg13g2_nor2_1 _12734_ (.A(_04039_),
    .B(_04858_),
    .Y(_04859_));
 sg13g2_nor2_1 _12735_ (.A(_04793_),
    .B(_04859_),
    .Y(_04860_));
 sg13g2_a21oi_1 _12736_ (.A1(net4341),
    .A2(_04806_),
    .Y(_04861_),
    .B1(_04844_));
 sg13g2_o21ai_1 _12737_ (.B1(_04861_),
    .Y(_04862_),
    .A1(_04855_),
    .A2(_04859_));
 sg13g2_mux2_1 _12738_ (.A0(net2606),
    .A1(_04862_),
    .S(_04852_),
    .X(_04863_));
 sg13g2_nor2b_1 _12739_ (.A(net1793),
    .B_N(_04863_),
    .Y(_00533_));
 sg13g2_nor2_1 _12740_ (.A(_04727_),
    .B(_04860_),
    .Y(_04864_));
 sg13g2_a21oi_1 _12741_ (.A1(_04852_),
    .A2(_04864_),
    .Y(_04865_),
    .B1(net2604));
 sg13g2_nor2_1 _12742_ (.A(net1793),
    .B(_04865_),
    .Y(_00534_));
 sg13g2_a21oi_1 _12743_ (.A1(net3561),
    .A2(net1810),
    .Y(_04866_),
    .B1(net1793));
 sg13g2_o21ai_1 _12744_ (.B1(_04866_),
    .Y(_00535_),
    .A1(_04824_),
    .A2(net1810));
 sg13g2_a21oi_1 _12745_ (.A1(net3744),
    .A2(net1810),
    .Y(_04867_),
    .B1(net1793));
 sg13g2_o21ai_1 _12746_ (.B1(_04867_),
    .Y(_00536_),
    .A1(net4600),
    .A2(net1810));
 sg13g2_a21oi_1 _12747_ (.A1(net4984),
    .A2(net1810),
    .Y(_04868_),
    .B1(net1793));
 sg13g2_nand2b_1 _12748_ (.Y(_00537_),
    .B(_04868_),
    .A_N(_04846_));
 sg13g2_a21oi_1 _12749_ (.A1(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .A2(_04834_),
    .Y(_04869_),
    .B1(net2604));
 sg13g2_nor4_1 _12750_ (.A(net2608),
    .B(_01982_),
    .C(_04793_),
    .D(_04869_),
    .Y(_04870_));
 sg13g2_o21ai_1 _12751_ (.B1(_04841_),
    .Y(_04871_),
    .A1(_04728_),
    .A2(_04792_));
 sg13g2_and2_1 _12752_ (.A(_04800_),
    .B(_04871_),
    .X(_04872_));
 sg13g2_nor4_1 _12753_ (.A(_04812_),
    .B(_04830_),
    .C(_04870_),
    .D(_04872_),
    .Y(_04873_));
 sg13g2_nor2_1 _12754_ (.A(net3874),
    .B(_04873_),
    .Y(_04874_));
 sg13g2_a21oi_1 _12755_ (.A1(_04729_),
    .A2(_04873_),
    .Y(_04875_),
    .B1(net1794));
 sg13g2_nor2b_1 _12756_ (.A(_04874_),
    .B_N(_04875_),
    .Y(_00538_));
 sg13g2_o21ai_1 _12757_ (.B1(_03167_),
    .Y(_04876_),
    .A1(_03145_),
    .A2(_03151_));
 sg13g2_nand2_2 _12758_ (.Y(_04877_),
    .A(_02817_),
    .B(_03145_));
 sg13g2_nor2_1 _12759_ (.A(_03161_),
    .B(_04877_),
    .Y(_04878_));
 sg13g2_nand2_1 _12760_ (.Y(_04879_),
    .A(net2365),
    .B(_02794_));
 sg13g2_nor2_2 _12761_ (.A(_02554_),
    .B(_02793_),
    .Y(_04880_));
 sg13g2_a21oi_1 _12762_ (.A1(_02730_),
    .A2(_04877_),
    .Y(_04881_),
    .B1(_04878_));
 sg13g2_nor2_2 _12763_ (.A(_04549_),
    .B(net2234),
    .Y(_04882_));
 sg13g2_o21ai_1 _12764_ (.B1(_04882_),
    .Y(_04883_),
    .A1(_02703_),
    .A2(_04880_));
 sg13g2_a21oi_1 _12765_ (.A1(_04880_),
    .A2(_04881_),
    .Y(_04884_),
    .B1(_04883_));
 sg13g2_a21o_1 _12766_ (.A2(net2234),
    .A1(net4963),
    .B1(_04884_),
    .X(_00539_));
 sg13g2_a21oi_1 _12767_ (.A1(_02683_),
    .A2(_04877_),
    .Y(_04885_),
    .B1(_04879_));
 sg13g2_o21ai_1 _12768_ (.B1(_04885_),
    .Y(_04886_),
    .A1(_03569_),
    .A2(_04877_));
 sg13g2_o21ai_1 _12769_ (.B1(_04882_),
    .Y(_04887_),
    .A1(_02667_),
    .A2(_04880_));
 sg13g2_inv_1 _12770_ (.Y(_04888_),
    .A(_04887_));
 sg13g2_a22oi_1 _12771_ (.Y(_04889_),
    .B1(_04886_),
    .B2(_04888_),
    .A2(net2234),
    .A1(net5042));
 sg13g2_inv_1 _12772_ (.Y(_00540_),
    .A(_04889_));
 sg13g2_nand2_1 _12773_ (.Y(_04890_),
    .A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B(_04806_));
 sg13g2_nor2_2 _12774_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .B(_04890_),
    .Y(_04891_));
 sg13g2_nor2_1 _12775_ (.A(net3719),
    .B(_04891_),
    .Y(_04892_));
 sg13g2_a21oi_1 _12776_ (.A1(_02042_),
    .A2(_04891_),
    .Y(_00541_),
    .B1(net3720));
 sg13g2_mux2_1 _12777_ (.A0(net4179),
    .A1(net11),
    .S(_04891_),
    .X(_00542_));
 sg13g2_mux2_1 _12778_ (.A0(net4090),
    .A1(net12),
    .S(_04891_),
    .X(_00543_));
 sg13g2_mux2_1 _12779_ (.A0(net4125),
    .A1(net13),
    .S(_04891_),
    .X(_00544_));
 sg13g2_nand2_1 _12780_ (.Y(_04893_),
    .A(net2614),
    .B(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_xor2_1 _12781_ (.B(\i_tinyqv.mem.q_ctrl.data_req ),
    .A(net2614),
    .X(_04894_));
 sg13g2_xnor2_1 _12782_ (.Y(_04895_),
    .A(net2614),
    .B(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_xnor2_1 _12783_ (.Y(_04896_),
    .A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_04893_));
 sg13g2_xnor2_1 _12784_ (.Y(_04897_),
    .A(_01983_),
    .B(_04893_));
 sg13g2_nor2_2 _12785_ (.A(_04790_),
    .B(_04792_),
    .Y(_04898_));
 sg13g2_o21ai_1 _12786_ (.B1(net2609),
    .Y(_04899_),
    .A1(_04790_),
    .A2(_04792_));
 sg13g2_nand2_1 _12787_ (.Y(_04900_),
    .A(_04819_),
    .B(net2228));
 sg13g2_nor4_1 _12788_ (.A(net2610),
    .B(net4910),
    .C(net5035),
    .D(_04796_),
    .Y(_04901_));
 sg13g2_a21oi_2 _12789_ (.B1(_04901_),
    .Y(_04902_),
    .A2(_04900_),
    .A1(_04820_));
 sg13g2_a21o_2 _12790_ (.A2(_04900_),
    .A1(_04820_),
    .B1(_04901_),
    .X(_04903_));
 sg13g2_and2_1 _12791_ (.A(_04037_),
    .B(_04798_),
    .X(_04904_));
 sg13g2_mux4_1 _12792_ (.S0(net2336),
    .A0(net2559),
    .A1(net2549),
    .A2(\data_to_write[16] ),
    .A3(\data_to_write[24] ),
    .S1(net2284),
    .X(_04905_));
 sg13g2_a21oi_1 _12793_ (.A1(_02042_),
    .A2(_04898_),
    .Y(_04906_),
    .B1(net2439));
 sg13g2_o21ai_1 _12794_ (.B1(_04906_),
    .Y(_04907_),
    .A1(_04898_),
    .A2(_04905_));
 sg13g2_nor2_1 _12795_ (.A(net3719),
    .B(_04904_),
    .Y(_04908_));
 sg13g2_a21oi_1 _12796_ (.A1(_02042_),
    .A2(_04904_),
    .Y(_04909_),
    .B1(_04908_));
 sg13g2_a21oi_1 _12797_ (.A1(net2439),
    .A2(_04909_),
    .Y(_04910_),
    .B1(_04902_));
 sg13g2_a22oi_1 _12798_ (.Y(_00545_),
    .B1(_04907_),
    .B2(_04910_),
    .A2(_04902_),
    .A1(_02038_));
 sg13g2_nand2_1 _12799_ (.Y(_04911_),
    .A(net2557),
    .B(net2334));
 sg13g2_a21oi_1 _12800_ (.A1(\data_to_write[9] ),
    .A2(net2336),
    .Y(_04912_),
    .B1(net2284));
 sg13g2_nand2_1 _12801_ (.Y(_04913_),
    .A(\data_to_write[17] ),
    .B(net2334));
 sg13g2_a21oi_1 _12802_ (.A1(\data_to_write[25] ),
    .A2(net2336),
    .Y(_04914_),
    .B1(_04897_));
 sg13g2_a221oi_1 _12803_ (.B2(_04914_),
    .C1(_04898_),
    .B1(_04913_),
    .A1(_04911_),
    .Y(_04915_),
    .A2(_04912_));
 sg13g2_a21oi_1 _12804_ (.A1(net11),
    .A2(_04898_),
    .Y(_04916_),
    .B1(_01981_));
 sg13g2_nand2b_1 _12805_ (.Y(_04917_),
    .B(_04916_),
    .A_N(_04915_));
 sg13g2_nand2b_1 _12806_ (.Y(_04918_),
    .B(net4179),
    .A_N(_04904_));
 sg13g2_a21oi_1 _12807_ (.A1(net11),
    .A2(_04904_),
    .Y(_04919_),
    .B1(net2610));
 sg13g2_a21oi_1 _12808_ (.A1(_04918_),
    .A2(_04919_),
    .Y(_04920_),
    .B1(_04902_));
 sg13g2_a22oi_1 _12809_ (.Y(_04921_),
    .B1(_04917_),
    .B2(_04920_),
    .A2(_04902_),
    .A1(net2603));
 sg13g2_inv_1 _12810_ (.Y(_00546_),
    .A(_04921_));
 sg13g2_nand2_1 _12811_ (.Y(_04922_),
    .A(net2556),
    .B(net2334));
 sg13g2_a21oi_1 _12812_ (.A1(\data_to_write[10] ),
    .A2(net2336),
    .Y(_04923_),
    .B1(net2284));
 sg13g2_nand2_1 _12813_ (.Y(_04924_),
    .A(\data_to_write[18] ),
    .B(net2334));
 sg13g2_a21oi_1 _12814_ (.A1(\data_to_write[26] ),
    .A2(net2336),
    .Y(_04925_),
    .B1(_04897_));
 sg13g2_a221oi_1 _12815_ (.B2(_04925_),
    .C1(_04898_),
    .B1(_04924_),
    .A1(_04922_),
    .Y(_04926_),
    .A2(_04923_));
 sg13g2_a21oi_1 _12816_ (.A1(net12),
    .A2(_04898_),
    .Y(_04927_),
    .B1(_01981_));
 sg13g2_nand2b_1 _12817_ (.Y(_04928_),
    .B(_04927_),
    .A_N(_04926_));
 sg13g2_nand2b_1 _12818_ (.Y(_04929_),
    .B(net4090),
    .A_N(_04904_));
 sg13g2_a21oi_1 _12819_ (.A1(net12),
    .A2(_04904_),
    .Y(_04930_),
    .B1(net2610));
 sg13g2_a21oi_1 _12820_ (.A1(_04929_),
    .A2(_04930_),
    .Y(_04931_),
    .B1(_04902_));
 sg13g2_a22oi_1 _12821_ (.Y(_04932_),
    .B1(_04928_),
    .B2(_04931_),
    .A2(_04902_),
    .A1(net2601));
 sg13g2_inv_1 _12822_ (.Y(_00547_),
    .A(_04932_));
 sg13g2_nand2_1 _12823_ (.Y(_04933_),
    .A(net2599),
    .B(_04902_));
 sg13g2_a21oi_1 _12824_ (.A1(\data_to_write[27] ),
    .A2(net2335),
    .Y(_04934_),
    .B1(_04897_));
 sg13g2_o21ai_1 _12825_ (.B1(_04934_),
    .Y(_04935_),
    .A1(_01836_),
    .A2(net2335));
 sg13g2_nand2_1 _12826_ (.Y(_04936_),
    .A(\data_to_write[11] ),
    .B(net2336));
 sg13g2_a21oi_1 _12827_ (.A1(net2555),
    .A2(net2334),
    .Y(_04937_),
    .B1(net2284));
 sg13g2_a21oi_1 _12828_ (.A1(_04936_),
    .A2(_04937_),
    .Y(_04938_),
    .B1(_04898_));
 sg13g2_a221oi_1 _12829_ (.B2(_04938_),
    .C1(_01981_),
    .B1(_04935_),
    .A1(net13),
    .Y(_04939_),
    .A2(_04898_));
 sg13g2_mux2_1 _12830_ (.A0(net4125),
    .A1(net13),
    .S(_04904_),
    .X(_04940_));
 sg13g2_o21ai_1 _12831_ (.B1(net2054),
    .Y(_04941_),
    .A1(net2610),
    .A2(_04940_));
 sg13g2_o21ai_1 _12832_ (.B1(_04933_),
    .Y(_00548_),
    .A1(_04939_),
    .A2(_04941_));
 sg13g2_nor2_1 _12833_ (.A(net2597),
    .B(net2054),
    .Y(_04942_));
 sg13g2_nand2_1 _12834_ (.Y(_04943_),
    .A(\data_to_write[12] ),
    .B(net2335));
 sg13g2_a21oi_1 _12835_ (.A1(net2554),
    .A2(net2333),
    .Y(_04944_),
    .B1(net2284));
 sg13g2_nand2_1 _12836_ (.Y(_04945_),
    .A(net4994),
    .B(net2334));
 sg13g2_a21oi_1 _12837_ (.A1(\data_to_write[28] ),
    .A2(net2335),
    .Y(_04946_),
    .B1(_04897_));
 sg13g2_a221oi_1 _12838_ (.B2(_04946_),
    .C1(net2228),
    .B1(_04945_),
    .A1(_04943_),
    .Y(_04947_),
    .A2(_04944_));
 sg13g2_a21oi_1 _12839_ (.A1(net5266),
    .A2(net2228),
    .Y(_04948_),
    .B1(_04947_));
 sg13g2_a21oi_1 _12840_ (.A1(net2054),
    .A2(net5267),
    .Y(_00549_),
    .B1(_04942_));
 sg13g2_nor2_1 _12841_ (.A(net2595),
    .B(net2054),
    .Y(_04949_));
 sg13g2_nor2_1 _12842_ (.A(_01816_),
    .B(net2333),
    .Y(_04950_));
 sg13g2_a21oi_1 _12843_ (.A1(\data_to_write[21] ),
    .A2(net2333),
    .Y(_04951_),
    .B1(_04950_));
 sg13g2_nand2_1 _12844_ (.Y(_04952_),
    .A(net5053),
    .B(net2336));
 sg13g2_a21oi_1 _12845_ (.A1(net2553),
    .A2(net2333),
    .Y(_04953_),
    .B1(net2284));
 sg13g2_a221oi_1 _12846_ (.B2(_04953_),
    .C1(net2228),
    .B1(_04952_),
    .A1(net2284),
    .Y(_04954_),
    .A2(_04951_));
 sg13g2_a21oi_1 _12847_ (.A1(net2603),
    .A2(net2228),
    .Y(_04955_),
    .B1(_04954_));
 sg13g2_a21oi_1 _12848_ (.A1(net2054),
    .A2(_04955_),
    .Y(_00550_),
    .B1(_04949_));
 sg13g2_nor2_1 _12849_ (.A(net2593),
    .B(net2054),
    .Y(_04956_));
 sg13g2_nand2_1 _12850_ (.Y(_04957_),
    .A(net5005),
    .B(net2335));
 sg13g2_a21oi_1 _12851_ (.A1(\data_to_write[22] ),
    .A2(net2333),
    .Y(_04958_),
    .B1(_04897_));
 sg13g2_nand2_1 _12852_ (.Y(_04959_),
    .A(net4962),
    .B(net2335));
 sg13g2_a21oi_1 _12853_ (.A1(net2552),
    .A2(net2333),
    .Y(_04960_),
    .B1(_04896_));
 sg13g2_a221oi_1 _12854_ (.B2(_04960_),
    .C1(net2228),
    .B1(_04959_),
    .A1(_04957_),
    .Y(_04961_),
    .A2(_04958_));
 sg13g2_a21oi_1 _12855_ (.A1(net2601),
    .A2(net2228),
    .Y(_04962_),
    .B1(_04961_));
 sg13g2_a21oi_1 _12856_ (.A1(net2054),
    .A2(_04962_),
    .Y(_00551_),
    .B1(_04956_));
 sg13g2_nor2_1 _12857_ (.A(net2591),
    .B(net2054),
    .Y(_04963_));
 sg13g2_nand2_1 _12858_ (.Y(_04964_),
    .A(\data_to_write[31] ),
    .B(net2335));
 sg13g2_a21oi_1 _12859_ (.A1(\data_to_write[23] ),
    .A2(net2333),
    .Y(_04965_),
    .B1(_04897_));
 sg13g2_nand2_1 _12860_ (.Y(_04966_),
    .A(\data_to_write[15] ),
    .B(net2335));
 sg13g2_a21oi_1 _12861_ (.A1(net2551),
    .A2(net2333),
    .Y(_04967_),
    .B1(net2284));
 sg13g2_a221oi_1 _12862_ (.B2(_04967_),
    .C1(net2228),
    .B1(_04966_),
    .A1(_04964_),
    .Y(_04968_),
    .A2(_04965_));
 sg13g2_a21oi_1 _12863_ (.A1(net2599),
    .A2(_04899_),
    .Y(_04969_),
    .B1(_04968_));
 sg13g2_a21oi_1 _12864_ (.A1(_04903_),
    .A2(_04969_),
    .Y(_00552_),
    .B1(_04963_));
 sg13g2_nand2b_1 _12865_ (.Y(_00553_),
    .B(net2620),
    .A_N(net3561));
 sg13g2_nand2b_1 _12866_ (.Y(_00554_),
    .B(net2620),
    .A_N(net3744));
 sg13g2_and2_1 _12867_ (.A(net2630),
    .B(_04779_),
    .X(_00555_));
 sg13g2_nor2_1 _12868_ (.A(net2442),
    .B(net1812),
    .Y(_04970_));
 sg13g2_a22oi_1 _12869_ (.Y(_00556_),
    .B1(_04970_),
    .B2(_02005_),
    .A2(net1812),
    .A1(_02035_));
 sg13g2_a22oi_1 _12870_ (.Y(_00557_),
    .B1(_04970_),
    .B2(_02008_),
    .A2(net1812),
    .A1(_02036_));
 sg13g2_mux2_1 _12871_ (.A0(net12),
    .A1(net4707),
    .S(net2623),
    .X(_00558_));
 sg13g2_nor2_1 _12872_ (.A(net2587),
    .B(net2233),
    .Y(_04971_));
 sg13g2_a21oi_1 _12873_ (.A1(_02048_),
    .A2(net2233),
    .Y(_00559_),
    .B1(_04971_));
 sg13g2_nor2_1 _12874_ (.A(net4689),
    .B(net2233),
    .Y(_04972_));
 sg13g2_a21oi_1 _12875_ (.A1(_02047_),
    .A2(net2233),
    .Y(_00560_),
    .B1(_04972_));
 sg13g2_mux2_1 _12876_ (.A0(net4997),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .S(net2234),
    .X(_00561_));
 sg13g2_mux2_1 _12877_ (.A0(net4995),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .S(net2234),
    .X(_00562_));
 sg13g2_mux2_1 _12878_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .A1(net4791),
    .S(net2233),
    .X(_00563_));
 sg13g2_mux2_1 _12879_ (.A0(net2582),
    .A1(net2586),
    .S(net2229),
    .X(_00564_));
 sg13g2_mux2_1 _12880_ (.A0(net2581),
    .A1(net2585),
    .S(net2229),
    .X(_00565_));
 sg13g2_mux2_1 _12881_ (.A0(net2580),
    .A1(net2584),
    .S(net2229),
    .X(_00566_));
 sg13g2_mux2_1 _12882_ (.A0(net2579),
    .A1(net2583),
    .S(net2229),
    .X(_00567_));
 sg13g2_mux2_1 _12883_ (.A0(net2578),
    .A1(net2582),
    .S(net2229),
    .X(_00568_));
 sg13g2_mux2_1 _12884_ (.A0(net2577),
    .A1(net2581),
    .S(net2229),
    .X(_00569_));
 sg13g2_mux2_1 _12885_ (.A0(net2576),
    .A1(net2580),
    .S(net2229),
    .X(_00570_));
 sg13g2_mux2_1 _12886_ (.A0(net4808),
    .A1(net2579),
    .S(net2232),
    .X(_00571_));
 sg13g2_mux2_1 _12887_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(net4736),
    .S(net2230),
    .X(_00572_));
 sg13g2_mux2_1 _12888_ (.A0(net4851),
    .A1(net2577),
    .S(net2229),
    .X(_00573_));
 sg13g2_mux2_1 _12889_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(net4758),
    .S(net2230),
    .X(_00574_));
 sg13g2_mux2_1 _12890_ (.A0(net4795),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net2232),
    .X(_00575_));
 sg13g2_mux2_1 _12891_ (.A0(net4947),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(net2230),
    .X(_00576_));
 sg13g2_mux2_1 _12892_ (.A0(net4887),
    .A1(net4851),
    .S(net2231),
    .X(_00577_));
 sg13g2_mux2_1 _12893_ (.A0(net4929),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(net2230),
    .X(_00578_));
 sg13g2_mux2_1 _12894_ (.A0(net4798),
    .A1(net4795),
    .S(net2231),
    .X(_00579_));
 sg13g2_mux2_1 _12895_ (.A0(net4961),
    .A1(net4947),
    .S(net2230),
    .X(_00580_));
 sg13g2_mux2_1 _12896_ (.A0(net4942),
    .A1(net4887),
    .S(net2230),
    .X(_00581_));
 sg13g2_mux2_1 _12897_ (.A0(net4811),
    .A1(net4929),
    .S(net2230),
    .X(_00582_));
 sg13g2_mux2_1 _12898_ (.A0(net4963),
    .A1(net4798),
    .S(net2230),
    .X(_00583_));
 sg13g2_mux2_1 _12899_ (.A0(net5042),
    .A1(net4961),
    .S(net2233),
    .X(_00584_));
 sg13g2_mux2_1 _12900_ (.A0(net5004),
    .A1(net4942),
    .S(net2231),
    .X(_00585_));
 sg13g2_mux2_1 _12901_ (.A0(net5146),
    .A1(net4811),
    .S(net2233),
    .X(_00586_));
 sg13g2_a21oi_1 _12902_ (.A1(_03869_),
    .A2(_03871_),
    .Y(_04973_),
    .B1(_04877_));
 sg13g2_a21oi_1 _12903_ (.A1(_02652_),
    .A2(_04877_),
    .Y(_04974_),
    .B1(_04879_));
 sg13g2_nor2b_1 _12904_ (.A(_04973_),
    .B_N(_04974_),
    .Y(_04975_));
 sg13g2_o21ai_1 _12905_ (.B1(_04882_),
    .Y(_04976_),
    .A1(_02626_),
    .A2(_04880_));
 sg13g2_a22oi_1 _12906_ (.Y(_04977_),
    .B1(net2233),
    .B2(net5004),
    .A2(_04546_),
    .A1(net4945));
 sg13g2_o21ai_1 _12907_ (.B1(_04977_),
    .Y(_00587_),
    .A1(_04975_),
    .A2(_04976_));
 sg13g2_nor2b_1 _12908_ (.A(net2234),
    .B_N(_04547_),
    .Y(_04978_));
 sg13g2_a21oi_1 _12909_ (.A1(net5146),
    .A2(net2234),
    .Y(_04979_),
    .B1(_04978_));
 sg13g2_o21ai_1 _12910_ (.B1(_04880_),
    .Y(_04980_),
    .A1(_04005_),
    .A2(_04877_));
 sg13g2_a21oi_1 _12911_ (.A1(_02604_),
    .A2(_04877_),
    .Y(_04981_),
    .B1(_04980_));
 sg13g2_o21ai_1 _12912_ (.B1(_04882_),
    .Y(_04982_),
    .A1(_02537_),
    .A2(_04880_));
 sg13g2_o21ai_1 _12913_ (.B1(_04979_),
    .Y(_00588_),
    .A1(_04981_),
    .A2(_04982_));
 sg13g2_nand2b_1 _12914_ (.Y(_04983_),
    .B(net3398),
    .A_N(net1879));
 sg13g2_nand2_1 _12915_ (.Y(_04984_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_xnor2_1 _12916_ (.Y(_04985_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_nand2_1 _12917_ (.Y(_04986_),
    .A(net2363),
    .B(_04985_));
 sg13g2_nand2b_1 _12918_ (.Y(_04987_),
    .B(net2294),
    .A_N(net2586));
 sg13g2_o21ai_1 _12919_ (.B1(_04987_),
    .Y(_04988_),
    .A1(net4481),
    .A2(net2294));
 sg13g2_nand2_1 _12920_ (.Y(_04989_),
    .A(net2359),
    .B(_04988_));
 sg13g2_nand3_1 _12921_ (.B(_04986_),
    .C(_04989_),
    .A(net1879),
    .Y(_04990_));
 sg13g2_o21ai_1 _12922_ (.B1(_04990_),
    .Y(_04991_),
    .A1(_04648_),
    .A2(_04983_));
 sg13g2_nor2_1 _12923_ (.A(_03630_),
    .B(_04650_),
    .Y(_04992_));
 sg13g2_and2_1 _12924_ (.A(_02827_),
    .B(_04649_),
    .X(_04993_));
 sg13g2_nand2_1 _12925_ (.Y(_04994_),
    .A(_02827_),
    .B(_04649_));
 sg13g2_nor3_1 _12926_ (.A(_04991_),
    .B(_04992_),
    .C(net1849),
    .Y(_04995_));
 sg13g2_o21ai_1 _12927_ (.B1(net2496),
    .Y(_04996_),
    .A1(net5285),
    .A2(net1845));
 sg13g2_nor2_1 _12928_ (.A(_04995_),
    .B(_04996_),
    .Y(_00589_));
 sg13g2_nand2b_1 _12929_ (.Y(_04997_),
    .B(net3403),
    .A_N(net1882));
 sg13g2_and2_1 _12930_ (.A(net4275),
    .B(net2298),
    .X(_04998_));
 sg13g2_a21oi_2 _12931_ (.B1(_04998_),
    .Y(_04999_),
    .A2(net2295),
    .A1(net2585));
 sg13g2_nor2_1 _12932_ (.A(\i_tinyqv.cpu.pc[2] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .Y(_05000_));
 sg13g2_nand2_1 _12933_ (.Y(_05001_),
    .A(\i_tinyqv.cpu.pc[2] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sg13g2_nor2b_1 _12934_ (.A(_05000_),
    .B_N(_05001_),
    .Y(_05002_));
 sg13g2_xnor2_1 _12935_ (.Y(_05003_),
    .A(_04984_),
    .B(_05002_));
 sg13g2_nor2_1 _12936_ (.A(net2359),
    .B(_05003_),
    .Y(_05004_));
 sg13g2_a21oi_1 _12937_ (.A1(net2360),
    .A2(_04999_),
    .Y(_05005_),
    .B1(_05004_));
 sg13g2_nand2_1 _12938_ (.Y(_05006_),
    .A(net1883),
    .B(_05005_));
 sg13g2_o21ai_1 _12939_ (.B1(_05006_),
    .Y(_05007_),
    .A1(net1865),
    .A2(_04997_));
 sg13g2_nor2_1 _12940_ (.A(_03760_),
    .B(_04650_),
    .Y(_05008_));
 sg13g2_nor3_1 _12941_ (.A(net1849),
    .B(_05007_),
    .C(_05008_),
    .Y(_05009_));
 sg13g2_o21ai_1 _12942_ (.B1(net2496),
    .Y(_05010_),
    .A1(net5260),
    .A2(net1845));
 sg13g2_nor2_1 _12943_ (.A(_05009_),
    .B(_05010_),
    .Y(_00590_));
 sg13g2_nand2b_1 _12944_ (.Y(_05011_),
    .B(_04571_),
    .A_N(net2584));
 sg13g2_o21ai_1 _12945_ (.B1(_05011_),
    .Y(_05012_),
    .A1(net4512),
    .A2(net2295));
 sg13g2_and2_1 _12946_ (.A(net2574),
    .B(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .X(_05013_));
 sg13g2_xor2_1 _12947_ (.B(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .A(net2574),
    .X(_05014_));
 sg13g2_o21ai_1 _12948_ (.B1(_05001_),
    .Y(_05015_),
    .A1(_04984_),
    .A2(_05000_));
 sg13g2_xor2_1 _12949_ (.B(_05015_),
    .A(_05014_),
    .X(_05016_));
 sg13g2_nor2_1 _12950_ (.A(net2360),
    .B(_05016_),
    .Y(_05017_));
 sg13g2_a21oi_1 _12951_ (.A1(net2360),
    .A2(_05012_),
    .Y(_05018_),
    .B1(_05017_));
 sg13g2_a21oi_1 _12952_ (.A1(net1882),
    .A2(_05018_),
    .Y(_05019_),
    .B1(net1850));
 sg13g2_nand2_1 _12953_ (.Y(_05020_),
    .A(_03885_),
    .B(net1865));
 sg13g2_o21ai_1 _12954_ (.B1(_05020_),
    .Y(_05021_),
    .A1(net3399),
    .A2(net1866));
 sg13g2_o21ai_1 _12955_ (.B1(_05019_),
    .Y(_05022_),
    .A1(net1882),
    .A2(_05021_));
 sg13g2_o21ai_1 _12956_ (.B1(_05022_),
    .Y(_05023_),
    .A1(net2575),
    .A2(net1847));
 sg13g2_nor2_1 _12957_ (.A(net2445),
    .B(_05023_),
    .Y(_00596_));
 sg13g2_nand2_1 _12958_ (.Y(_05024_),
    .A(_03365_),
    .B(net1865));
 sg13g2_a21oi_1 _12959_ (.A1(net3387),
    .A2(net1869),
    .Y(_05025_),
    .B1(net1880));
 sg13g2_nand2b_1 _12960_ (.Y(_05026_),
    .B(net2294),
    .A_N(net2583));
 sg13g2_o21ai_1 _12961_ (.B1(_05026_),
    .Y(_05027_),
    .A1(net3682),
    .A2(net2294));
 sg13g2_nand2_1 _12962_ (.Y(_05028_),
    .A(net2573),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_xnor2_1 _12963_ (.Y(_05029_),
    .A(net2573),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_a21oi_1 _12964_ (.A1(_05014_),
    .A2(_05015_),
    .Y(_05030_),
    .B1(_05013_));
 sg13g2_xnor2_1 _12965_ (.Y(_05031_),
    .A(_05029_),
    .B(_05030_));
 sg13g2_mux2_1 _12966_ (.A0(_05027_),
    .A1(_05031_),
    .S(net2364),
    .X(_05032_));
 sg13g2_a221oi_1 _12967_ (.B2(net1882),
    .C1(net1850),
    .B1(_05032_),
    .A1(_05024_),
    .Y(_05033_),
    .A2(_05025_));
 sg13g2_a21o_1 _12968_ (.A2(net1850),
    .A1(net2573),
    .B1(_05033_),
    .X(_05034_));
 sg13g2_and2_1 _12969_ (.A(net2501),
    .B(_05034_),
    .X(_00597_));
 sg13g2_and2_1 _12970_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .X(_05035_));
 sg13g2_xor2_1 _12971_ (.B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(_05036_));
 sg13g2_o21ai_1 _12972_ (.B1(_05028_),
    .Y(_05037_),
    .A1(_05029_),
    .A2(_05030_));
 sg13g2_xnor2_1 _12973_ (.Y(_05038_),
    .A(_05036_),
    .B(_05037_));
 sg13g2_mux2_1 _12974_ (.A0(net2582),
    .A1(\i_tinyqv.cpu.i_core.mepc[5] ),
    .S(net2297),
    .X(_05039_));
 sg13g2_o21ai_1 _12975_ (.B1(net1883),
    .Y(_05040_),
    .A1(net2364),
    .A2(_05039_));
 sg13g2_a21oi_1 _12976_ (.A1(net2364),
    .A2(_05038_),
    .Y(_05041_),
    .B1(_05040_));
 sg13g2_nor2_1 _12977_ (.A(net1851),
    .B(_05041_),
    .Y(_05042_));
 sg13g2_nand2_1 _12978_ (.Y(_05043_),
    .A(_03629_),
    .B(net1866));
 sg13g2_o21ai_1 _12979_ (.B1(_05043_),
    .Y(_05044_),
    .A1(net3391),
    .A2(net1865));
 sg13g2_o21ai_1 _12980_ (.B1(_05042_),
    .Y(_05045_),
    .A1(net1882),
    .A2(_05044_));
 sg13g2_o21ai_1 _12981_ (.B1(_05045_),
    .Y(_05046_),
    .A1(net5262),
    .A2(net1847));
 sg13g2_nor2_1 _12982_ (.A(net2445),
    .B(_05046_),
    .Y(_00598_));
 sg13g2_nor2_1 _12983_ (.A(_03758_),
    .B(net1870),
    .Y(_05047_));
 sg13g2_a221oi_1 _12984_ (.B2(net3392),
    .C1(_05047_),
    .B1(net1869),
    .A1(net2317),
    .Y(_05048_),
    .A2(_04573_));
 sg13g2_nand2b_1 _12985_ (.Y(_05049_),
    .B(net2294),
    .A_N(net2581));
 sg13g2_o21ai_1 _12986_ (.B1(_05049_),
    .Y(_05050_),
    .A1(net4510),
    .A2(net2294));
 sg13g2_nand2_1 _12987_ (.Y(_05051_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_xnor2_1 _12988_ (.Y(_05052_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_a21oi_1 _12989_ (.A1(_05036_),
    .A2(_05037_),
    .Y(_05053_),
    .B1(_05035_));
 sg13g2_xnor2_1 _12990_ (.Y(_05054_),
    .A(_05052_),
    .B(_05053_));
 sg13g2_mux2_1 _12991_ (.A0(_05050_),
    .A1(_05054_),
    .S(net2364),
    .X(_05055_));
 sg13g2_a221oi_1 _12992_ (.B2(net1882),
    .C1(_05048_),
    .B1(_05055_),
    .A1(_02827_),
    .Y(_05056_),
    .A2(_04649_));
 sg13g2_a21oi_1 _12993_ (.A1(net5001),
    .A2(net1851),
    .Y(_05057_),
    .B1(_05056_));
 sg13g2_nor2_1 _12994_ (.A(net2445),
    .B(_05057_),
    .Y(_00599_));
 sg13g2_nor2_1 _12995_ (.A(_03883_),
    .B(net1869),
    .Y(_05058_));
 sg13g2_and2_1 _12996_ (.A(net2572),
    .B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(_05059_));
 sg13g2_xor2_1 _12997_ (.B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .A(net2572),
    .X(_05060_));
 sg13g2_o21ai_1 _12998_ (.B1(_05051_),
    .Y(_05061_),
    .A1(_05052_),
    .A2(_05053_));
 sg13g2_xnor2_1 _12999_ (.Y(_05062_),
    .A(_05060_),
    .B(_05061_));
 sg13g2_and2_1 _13000_ (.A(\i_tinyqv.cpu.i_core.mepc[7] ),
    .B(net2297),
    .X(_05063_));
 sg13g2_a21oi_2 _13001_ (.B1(_05063_),
    .Y(_05064_),
    .A2(net2295),
    .A1(net2580));
 sg13g2_and2_1 _13002_ (.A(_02563_),
    .B(_05064_),
    .X(_05065_));
 sg13g2_a21oi_1 _13003_ (.A1(net2364),
    .A2(_05062_),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_a21oi_1 _13004_ (.A1(net3382),
    .A2(net1870),
    .Y(_05067_),
    .B1(_05058_));
 sg13g2_a21oi_1 _13005_ (.A1(net1881),
    .A2(_05066_),
    .Y(_05068_),
    .B1(net1850));
 sg13g2_o21ai_1 _13006_ (.B1(_05068_),
    .Y(_05069_),
    .A1(net1880),
    .A2(_05067_));
 sg13g2_o21ai_1 _13007_ (.B1(_05069_),
    .Y(_05070_),
    .A1(net2572),
    .A2(net1847));
 sg13g2_nor2_1 _13008_ (.A(net2444),
    .B(_05070_),
    .Y(_00600_));
 sg13g2_nand2_1 _13009_ (.Y(_05071_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_xnor2_1 _13010_ (.Y(_05072_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_a21oi_1 _13011_ (.A1(_05060_),
    .A2(_05061_),
    .Y(_05073_),
    .B1(_05059_));
 sg13g2_xor2_1 _13012_ (.B(_05073_),
    .A(_05072_),
    .X(_05074_));
 sg13g2_nor2_1 _13013_ (.A(net2360),
    .B(_05074_),
    .Y(_05075_));
 sg13g2_and2_1 _13014_ (.A(\i_tinyqv.cpu.i_core.mepc[8] ),
    .B(_04570_),
    .X(_05076_));
 sg13g2_a21oi_2 _13015_ (.B1(_05076_),
    .Y(_05077_),
    .A2(_04571_),
    .A1(net2579));
 sg13g2_a21oi_1 _13016_ (.A1(net2360),
    .A2(_05077_),
    .Y(_05078_),
    .B1(_05075_));
 sg13g2_a21oi_1 _13017_ (.A1(net1881),
    .A2(_05078_),
    .Y(_05079_),
    .B1(net1850));
 sg13g2_or2_1 _13018_ (.X(_05080_),
    .B(net1869),
    .A(_03367_));
 sg13g2_o21ai_1 _13019_ (.B1(_05080_),
    .Y(_05081_),
    .A1(net3388),
    .A2(net1866));
 sg13g2_o21ai_1 _13020_ (.B1(_05079_),
    .Y(_05082_),
    .A1(net1881),
    .A2(_05081_));
 sg13g2_o21ai_1 _13021_ (.B1(_05082_),
    .Y(_05083_),
    .A1(net5199),
    .A2(net1847));
 sg13g2_nor2_1 _13022_ (.A(net2444),
    .B(_05083_),
    .Y(_00601_));
 sg13g2_a21oi_1 _13023_ (.A1(_03632_),
    .A2(net1866),
    .Y(_05084_),
    .B1(net1880));
 sg13g2_o21ai_1 _13024_ (.B1(_05084_),
    .Y(_05085_),
    .A1(net3395),
    .A2(net1866));
 sg13g2_nand2b_1 _13025_ (.Y(_05086_),
    .B(net2293),
    .A_N(net2578));
 sg13g2_o21ai_1 _13026_ (.B1(_05086_),
    .Y(_05087_),
    .A1(\i_tinyqv.cpu.i_core.mepc[9] ),
    .A2(net2294));
 sg13g2_o21ai_1 _13027_ (.B1(_05071_),
    .Y(_05088_),
    .A1(_05072_),
    .A2(_05073_));
 sg13g2_and2_1 _13028_ (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .X(_05089_));
 sg13g2_xor2_1 _13029_ (.B(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .A(\i_tinyqv.cpu.instr_data_start[9] ),
    .X(_05090_));
 sg13g2_xor2_1 _13030_ (.B(_05090_),
    .A(_05088_),
    .X(_05091_));
 sg13g2_nand2_1 _13031_ (.Y(_05092_),
    .A(net2363),
    .B(_05091_));
 sg13g2_o21ai_1 _13032_ (.B1(_05092_),
    .Y(_05093_),
    .A1(net2363),
    .A2(_05087_));
 sg13g2_a21oi_1 _13033_ (.A1(net1880),
    .A2(_05093_),
    .Y(_05094_),
    .B1(net1850));
 sg13g2_a221oi_1 _13034_ (.B2(_05094_),
    .C1(net2443),
    .B1(_05085_),
    .A1(_01975_),
    .Y(_00602_),
    .A2(net1850));
 sg13g2_a21oi_1 _13035_ (.A1(_03756_),
    .A2(net1865),
    .Y(_05095_),
    .B1(net1883));
 sg13g2_o21ai_1 _13036_ (.B1(_05095_),
    .Y(_05096_),
    .A1(net3389),
    .A2(net1865));
 sg13g2_nand2b_1 _13037_ (.Y(_05097_),
    .B(net2293),
    .A_N(net2577));
 sg13g2_o21ai_1 _13038_ (.B1(_05097_),
    .Y(_05098_),
    .A1(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A2(net2294));
 sg13g2_a21oi_1 _13039_ (.A1(_05088_),
    .A2(_05090_),
    .Y(_05099_),
    .B1(_05089_));
 sg13g2_nor2_1 _13040_ (.A(net2570),
    .B(net2531),
    .Y(_05100_));
 sg13g2_xor2_1 _13041_ (.B(net2531),
    .A(net2570),
    .X(_05101_));
 sg13g2_xnor2_1 _13042_ (.Y(_05102_),
    .A(_05099_),
    .B(_05101_));
 sg13g2_nand2_1 _13043_ (.Y(_05103_),
    .A(net2363),
    .B(_05102_));
 sg13g2_o21ai_1 _13044_ (.B1(_05103_),
    .Y(_05104_),
    .A1(net2363),
    .A2(_05098_));
 sg13g2_a21oi_1 _13045_ (.A1(net1879),
    .A2(_05104_),
    .Y(_05105_),
    .B1(net1850));
 sg13g2_o21ai_1 _13046_ (.B1(net2497),
    .Y(_05106_),
    .A1(net2570),
    .A2(net1847));
 sg13g2_a21oi_1 _13047_ (.A1(_05096_),
    .A2(_05105_),
    .Y(_00603_),
    .B1(_05106_));
 sg13g2_nand2_1 _13048_ (.Y(_05107_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sg13g2_xnor2_1 _13049_ (.Y(_05108_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[11] ));
 sg13g2_a221oi_1 _13050_ (.B2(_05090_),
    .C1(_05089_),
    .B1(_05088_),
    .A1(net2570),
    .Y(_05109_),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[10] ));
 sg13g2_o21ai_1 _13051_ (.B1(_05108_),
    .Y(_05110_),
    .A1(_05100_),
    .A2(_05109_));
 sg13g2_or3_1 _13052_ (.A(_05100_),
    .B(_05108_),
    .C(_05109_),
    .X(_05111_));
 sg13g2_and2_1 _13053_ (.A(_05110_),
    .B(_05111_),
    .X(_05112_));
 sg13g2_nor2_1 _13054_ (.A(net2359),
    .B(_05112_),
    .Y(_05113_));
 sg13g2_and2_1 _13055_ (.A(\i_tinyqv.cpu.i_core.mepc[11] ),
    .B(net2296),
    .X(_05114_));
 sg13g2_a21oi_2 _13056_ (.B1(_05114_),
    .Y(_05115_),
    .A2(net2293),
    .A1(net2576));
 sg13g2_a21oi_1 _13057_ (.A1(net2359),
    .A2(_05115_),
    .Y(_05116_),
    .B1(_05113_));
 sg13g2_a21oi_1 _13058_ (.A1(net1878),
    .A2(_05116_),
    .Y(_05117_),
    .B1(net1848));
 sg13g2_nand2_1 _13059_ (.Y(_05118_),
    .A(_03888_),
    .B(net1864));
 sg13g2_o21ai_1 _13060_ (.B1(_05118_),
    .Y(_05119_),
    .A1(net3390),
    .A2(net1864));
 sg13g2_o21ai_1 _13061_ (.B1(_05117_),
    .Y(_05120_),
    .A1(net1878),
    .A2(_05119_));
 sg13g2_o21ai_1 _13062_ (.B1(_05120_),
    .Y(_05121_),
    .A1(net5244),
    .A2(net1846));
 sg13g2_nor2_1 _13063_ (.A(net2443),
    .B(_05121_),
    .Y(_00604_));
 sg13g2_mux2_1 _13064_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[12] ),
    .S(net2297),
    .X(_05122_));
 sg13g2_nand2_1 _13065_ (.Y(_05123_),
    .A(_05107_),
    .B(_05111_));
 sg13g2_nor2_1 _13066_ (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(\i_tinyqv.cpu.imm[12] ),
    .Y(_05124_));
 sg13g2_and2_1 _13067_ (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(\i_tinyqv.cpu.imm[12] ),
    .X(_05125_));
 sg13g2_nor2_1 _13068_ (.A(_05124_),
    .B(_05125_),
    .Y(_05126_));
 sg13g2_xnor2_1 _13069_ (.Y(_05127_),
    .A(_05123_),
    .B(_05126_));
 sg13g2_nor2_1 _13070_ (.A(net2360),
    .B(_05127_),
    .Y(_05128_));
 sg13g2_a21oi_1 _13071_ (.A1(net2359),
    .A2(_05122_),
    .Y(_05129_),
    .B1(_05128_));
 sg13g2_mux2_1 _13072_ (.A0(_03369_),
    .A1(net3377),
    .S(net1868),
    .X(_05130_));
 sg13g2_nand2_1 _13073_ (.Y(_05131_),
    .A(net1878),
    .B(_05129_));
 sg13g2_o21ai_1 _13074_ (.B1(_05131_),
    .Y(_05132_),
    .A1(net1878),
    .A2(_05130_));
 sg13g2_o21ai_1 _13075_ (.B1(net2496),
    .Y(_05133_),
    .A1(net5225),
    .A2(net1846));
 sg13g2_a21oi_1 _13076_ (.A1(net1846),
    .A2(_05132_),
    .Y(_00605_),
    .B1(_05133_));
 sg13g2_a21oi_1 _13077_ (.A1(_03628_),
    .A2(net1864),
    .Y(_05134_),
    .B1(net1880));
 sg13g2_o21ai_1 _13078_ (.B1(_05134_),
    .Y(_05135_),
    .A1(net3386),
    .A2(net1864));
 sg13g2_nand2_1 _13079_ (.Y(_05136_),
    .A(net2569),
    .B(\i_tinyqv.cpu.imm[13] ));
 sg13g2_xor2_1 _13080_ (.B(\i_tinyqv.cpu.imm[13] ),
    .A(net2569),
    .X(_05137_));
 sg13g2_a21oi_1 _13081_ (.A1(_05107_),
    .A2(_05111_),
    .Y(_05138_),
    .B1(_05124_));
 sg13g2_nor3_1 _13082_ (.A(_05125_),
    .B(_05137_),
    .C(_05138_),
    .Y(_05139_));
 sg13g2_o21ai_1 _13083_ (.B1(_05137_),
    .Y(_05140_),
    .A1(_05125_),
    .A2(_05138_));
 sg13g2_nand2b_1 _13084_ (.Y(_05141_),
    .B(_05140_),
    .A_N(_05139_));
 sg13g2_and2_1 _13085_ (.A(\i_tinyqv.cpu.i_core.mepc[13] ),
    .B(net2296),
    .X(_05142_));
 sg13g2_a21oi_2 _13086_ (.B1(_05142_),
    .Y(_05143_),
    .A2(net2293),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sg13g2_and2_1 _13087_ (.A(net2358),
    .B(_05143_),
    .X(_05144_));
 sg13g2_a21oi_1 _13088_ (.A1(net2361),
    .A2(_05141_),
    .Y(_05145_),
    .B1(_05144_));
 sg13g2_a21oi_1 _13089_ (.A1(net1876),
    .A2(_05145_),
    .Y(_05146_),
    .B1(net1848));
 sg13g2_o21ai_1 _13090_ (.B1(net2494),
    .Y(_05147_),
    .A1(net2569),
    .A2(net1845));
 sg13g2_a21oi_1 _13091_ (.A1(_05135_),
    .A2(_05146_),
    .Y(_00606_),
    .B1(_05147_));
 sg13g2_nor2_1 _13092_ (.A(net2568),
    .B(\i_tinyqv.cpu.imm[14] ),
    .Y(_05148_));
 sg13g2_and2_1 _13093_ (.A(net2568),
    .B(\i_tinyqv.cpu.imm[14] ),
    .X(_05149_));
 sg13g2_or2_1 _13094_ (.X(_05150_),
    .B(_05149_),
    .A(_05148_));
 sg13g2_nand2_1 _13095_ (.Y(_05151_),
    .A(_05136_),
    .B(_05140_));
 sg13g2_xnor2_1 _13096_ (.Y(_05152_),
    .A(_05150_),
    .B(_05151_));
 sg13g2_nand2_1 _13097_ (.Y(_05153_),
    .A(net2362),
    .B(_05152_));
 sg13g2_nand2b_1 _13098_ (.Y(_05154_),
    .B(net2292),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[18] ));
 sg13g2_o21ai_1 _13099_ (.B1(_05154_),
    .Y(_05155_),
    .A1(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A2(net2292));
 sg13g2_o21ai_1 _13100_ (.B1(_05153_),
    .Y(_05156_),
    .A1(net2362),
    .A2(_05155_));
 sg13g2_a21oi_1 _13101_ (.A1(net1879),
    .A2(_05156_),
    .Y(_05157_),
    .B1(net1849));
 sg13g2_a21oi_1 _13102_ (.A1(_03755_),
    .A2(net1865),
    .Y(_05158_),
    .B1(net1880));
 sg13g2_o21ai_1 _13103_ (.B1(_05158_),
    .Y(_05159_),
    .A1(net3385),
    .A2(net1865));
 sg13g2_a221oi_1 _13104_ (.B2(_05159_),
    .C1(net2443),
    .B1(_05157_),
    .A1(_01973_),
    .Y(_00607_),
    .A2(net1849));
 sg13g2_nand2_1 _13105_ (.Y(_05160_),
    .A(\i_tinyqv.cpu.instr_data_start[15] ),
    .B(\i_tinyqv.cpu.imm[15] ));
 sg13g2_xor2_1 _13106_ (.B(\i_tinyqv.cpu.imm[15] ),
    .A(\i_tinyqv.cpu.instr_data_start[15] ),
    .X(_05161_));
 sg13g2_a21oi_1 _13107_ (.A1(_05136_),
    .A2(_05140_),
    .Y(_05162_),
    .B1(_05148_));
 sg13g2_nor2_1 _13108_ (.A(_05149_),
    .B(_05162_),
    .Y(_05163_));
 sg13g2_o21ai_1 _13109_ (.B1(_05161_),
    .Y(_05164_),
    .A1(_05149_),
    .A2(_05162_));
 sg13g2_xor2_1 _13110_ (.B(_05163_),
    .A(_05161_),
    .X(_05165_));
 sg13g2_mux2_1 _13111_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(\i_tinyqv.cpu.i_core.mepc[15] ),
    .S(net2296),
    .X(_05166_));
 sg13g2_o21ai_1 _13112_ (.B1(net1877),
    .Y(_05167_),
    .A1(net2359),
    .A2(_05165_));
 sg13g2_a21o_1 _13113_ (.A2(_05166_),
    .A1(net2358),
    .B1(_05167_),
    .X(_05168_));
 sg13g2_nand2_1 _13114_ (.Y(_05169_),
    .A(net3381),
    .B(net1868));
 sg13g2_o21ai_1 _13115_ (.B1(_05169_),
    .Y(_05170_),
    .A1(_03882_),
    .A2(net1867));
 sg13g2_o21ai_1 _13116_ (.B1(_05168_),
    .Y(_05171_),
    .A1(net1877),
    .A2(_05170_));
 sg13g2_o21ai_1 _13117_ (.B1(net2494),
    .Y(_05172_),
    .A1(net5249),
    .A2(net1844));
 sg13g2_a21oi_1 _13118_ (.A1(net1844),
    .A2(_05171_),
    .Y(_00608_),
    .B1(_05172_));
 sg13g2_nor2_1 _13119_ (.A(net2567),
    .B(\i_tinyqv.cpu.imm[16] ),
    .Y(_05173_));
 sg13g2_and2_1 _13120_ (.A(net2567),
    .B(\i_tinyqv.cpu.imm[16] ),
    .X(_05174_));
 sg13g2_nor2_1 _13121_ (.A(_05173_),
    .B(_05174_),
    .Y(_05175_));
 sg13g2_nand2_1 _13122_ (.Y(_05176_),
    .A(_05160_),
    .B(_05164_));
 sg13g2_xor2_1 _13123_ (.B(_05176_),
    .A(_05175_),
    .X(_05177_));
 sg13g2_nand2b_1 _13124_ (.Y(_05178_),
    .B(net2292),
    .A_N(\i_tinyqv.cpu.i_core.i_shift.a[20] ));
 sg13g2_o21ai_1 _13125_ (.B1(_05178_),
    .Y(_05179_),
    .A1(\i_tinyqv.cpu.i_core.mepc[16] ),
    .A2(net2292));
 sg13g2_mux2_1 _13126_ (.A0(_03363_),
    .A1(net3384),
    .S(net1867),
    .X(_05180_));
 sg13g2_o21ai_1 _13127_ (.B1(net1877),
    .Y(_05181_),
    .A1(net2361),
    .A2(_05179_));
 sg13g2_a21o_1 _13128_ (.A2(_05177_),
    .A1(net2361),
    .B1(_05181_),
    .X(_05182_));
 sg13g2_o21ai_1 _13129_ (.B1(_05182_),
    .Y(_05183_),
    .A1(net1876),
    .A2(_05180_));
 sg13g2_o21ai_1 _13130_ (.B1(net2494),
    .Y(_05184_),
    .A1(net2567),
    .A2(net1844));
 sg13g2_a21oi_1 _13131_ (.A1(net1844),
    .A2(_05183_),
    .Y(_00609_),
    .B1(_05184_));
 sg13g2_nand2_1 _13132_ (.Y(_05185_),
    .A(net2566),
    .B(\i_tinyqv.cpu.imm[17] ));
 sg13g2_xor2_1 _13133_ (.B(\i_tinyqv.cpu.imm[17] ),
    .A(net2566),
    .X(_05186_));
 sg13g2_a21oi_1 _13134_ (.A1(_05160_),
    .A2(_05164_),
    .Y(_05187_),
    .B1(_05173_));
 sg13g2_nor2_1 _13135_ (.A(_05174_),
    .B(_05187_),
    .Y(_05188_));
 sg13g2_o21ai_1 _13136_ (.B1(_05186_),
    .Y(_05189_),
    .A1(_05174_),
    .A2(_05187_));
 sg13g2_xnor2_1 _13137_ (.Y(_05190_),
    .A(_05186_),
    .B(_05188_));
 sg13g2_mux2_1 _13138_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(net4551),
    .S(net2296),
    .X(_05191_));
 sg13g2_nand2_1 _13139_ (.Y(_05192_),
    .A(net2358),
    .B(_05191_));
 sg13g2_nand2_1 _13140_ (.Y(_05193_),
    .A(net2362),
    .B(_05190_));
 sg13g2_nand3_1 _13141_ (.B(_05192_),
    .C(_05193_),
    .A(net1877),
    .Y(_05194_));
 sg13g2_nand2_1 _13142_ (.Y(_05195_),
    .A(net3374),
    .B(net1867));
 sg13g2_o21ai_1 _13143_ (.B1(_05195_),
    .Y(_05196_),
    .A1(_03635_),
    .A2(net1867));
 sg13g2_o21ai_1 _13144_ (.B1(_05194_),
    .Y(_05197_),
    .A1(net1877),
    .A2(_05196_));
 sg13g2_o21ai_1 _13145_ (.B1(net2497),
    .Y(_05198_),
    .A1(net2566),
    .A2(net1845));
 sg13g2_a21oi_1 _13146_ (.A1(net1845),
    .A2(_05197_),
    .Y(_00610_),
    .B1(_05198_));
 sg13g2_a21oi_1 _13147_ (.A1(_02046_),
    .A2(net1870),
    .Y(_05199_),
    .B1(net1880));
 sg13g2_o21ai_1 _13148_ (.B1(_05199_),
    .Y(_05200_),
    .A1(_03753_),
    .A2(net1869));
 sg13g2_nand2_1 _13149_ (.Y(_05201_),
    .A(_05185_),
    .B(_05189_));
 sg13g2_nor2_1 _13150_ (.A(_01971_),
    .B(_01998_),
    .Y(_05202_));
 sg13g2_xnor2_1 _13151_ (.Y(_05203_),
    .A(\i_tinyqv.cpu.instr_data_start[18] ),
    .B(\i_tinyqv.cpu.imm[18] ));
 sg13g2_xnor2_1 _13152_ (.Y(_05204_),
    .A(_05201_),
    .B(_05203_));
 sg13g2_nor2_1 _13153_ (.A(net2359),
    .B(_05204_),
    .Y(_05205_));
 sg13g2_and2_1 _13154_ (.A(\i_tinyqv.cpu.i_core.mepc[18] ),
    .B(net2296),
    .X(_05206_));
 sg13g2_a21oi_2 _13155_ (.B1(_05206_),
    .Y(_05207_),
    .A2(net2292),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ));
 sg13g2_a21oi_1 _13156_ (.A1(net2358),
    .A2(_05207_),
    .Y(_05208_),
    .B1(_05205_));
 sg13g2_a21oi_1 _13157_ (.A1(net1877),
    .A2(_05208_),
    .Y(_05209_),
    .B1(net1848));
 sg13g2_a221oi_1 _13158_ (.B2(_05209_),
    .C1(net2443),
    .B1(_05200_),
    .A1(_01971_),
    .Y(_00611_),
    .A2(net1848));
 sg13g2_nand2_1 _13159_ (.Y(_05210_),
    .A(net2565),
    .B(\i_tinyqv.cpu.imm[19] ));
 sg13g2_xor2_1 _13160_ (.B(\i_tinyqv.cpu.imm[19] ),
    .A(net2565),
    .X(_05211_));
 sg13g2_a22oi_1 _13161_ (.Y(_05212_),
    .B1(_05185_),
    .B2(_05189_),
    .A2(_01998_),
    .A1(_01971_));
 sg13g2_nor2_1 _13162_ (.A(_05202_),
    .B(_05212_),
    .Y(_05213_));
 sg13g2_o21ai_1 _13163_ (.B1(_05211_),
    .Y(_05214_),
    .A1(_05202_),
    .A2(_05212_));
 sg13g2_xor2_1 _13164_ (.B(_05213_),
    .A(_05211_),
    .X(_05215_));
 sg13g2_mux2_1 _13165_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(net4296),
    .S(net2296),
    .X(_05216_));
 sg13g2_o21ai_1 _13166_ (.B1(net1876),
    .Y(_05217_),
    .A1(net2361),
    .A2(_05216_));
 sg13g2_a21oi_1 _13167_ (.A1(net2361),
    .A2(_05215_),
    .Y(_05218_),
    .B1(_05217_));
 sg13g2_nor2_1 _13168_ (.A(_03890_),
    .B(net1867),
    .Y(_05219_));
 sg13g2_a21oi_1 _13169_ (.A1(net3379),
    .A2(net1867),
    .Y(_05220_),
    .B1(_05219_));
 sg13g2_o21ai_1 _13170_ (.B1(net1846),
    .Y(_05221_),
    .A1(net1876),
    .A2(_05220_));
 sg13g2_o21ai_1 _13171_ (.B1(net2494),
    .Y(_05222_),
    .A1(_05218_),
    .A2(_05221_));
 sg13g2_a21oi_1 _13172_ (.A1(_01970_),
    .A2(net1848),
    .Y(_00612_),
    .B1(_05222_));
 sg13g2_nor2_1 _13173_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(\i_tinyqv.cpu.imm[20] ),
    .Y(_05223_));
 sg13g2_and2_1 _13174_ (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .B(\i_tinyqv.cpu.imm[20] ),
    .X(_05224_));
 sg13g2_or2_1 _13175_ (.X(_05225_),
    .B(_05224_),
    .A(_05223_));
 sg13g2_nand2_1 _13176_ (.Y(_05226_),
    .A(_05210_),
    .B(_05214_));
 sg13g2_xnor2_1 _13177_ (.Y(_05227_),
    .A(_05225_),
    .B(_05226_));
 sg13g2_nor2_1 _13178_ (.A(net2358),
    .B(_05227_),
    .Y(_05228_));
 sg13g2_and2_1 _13179_ (.A(net4061),
    .B(net2297),
    .X(_05229_));
 sg13g2_a21oi_2 _13180_ (.B1(_05229_),
    .Y(_05230_),
    .A2(net2293),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ));
 sg13g2_a21oi_1 _13181_ (.A1(net2358),
    .A2(_05230_),
    .Y(_05231_),
    .B1(_05228_));
 sg13g2_nand2b_1 _13182_ (.Y(_05232_),
    .B(net1867),
    .A_N(net3401));
 sg13g2_a21oi_1 _13183_ (.A1(_03362_),
    .A2(net1864),
    .Y(_05233_),
    .B1(net1878));
 sg13g2_a221oi_1 _13184_ (.B2(_05233_),
    .C1(net1848),
    .B1(_05232_),
    .A1(net1878),
    .Y(_05234_),
    .A2(_05231_));
 sg13g2_o21ai_1 _13185_ (.B1(net2495),
    .Y(_05235_),
    .A1(net5284),
    .A2(net1846));
 sg13g2_nor2_1 _13186_ (.A(_05234_),
    .B(_05235_),
    .Y(_00613_));
 sg13g2_and2_1 _13187_ (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(\i_tinyqv.cpu.imm[21] ),
    .X(_05236_));
 sg13g2_xor2_1 _13188_ (.B(\i_tinyqv.cpu.imm[21] ),
    .A(\i_tinyqv.cpu.instr_data_start[21] ),
    .X(_05237_));
 sg13g2_a21oi_1 _13189_ (.A1(_05210_),
    .A2(_05214_),
    .Y(_05238_),
    .B1(_05223_));
 sg13g2_or2_1 _13190_ (.X(_05239_),
    .B(_05238_),
    .A(_05224_));
 sg13g2_xnor2_1 _13191_ (.Y(_05240_),
    .A(_05237_),
    .B(_05239_));
 sg13g2_nand2_1 _13192_ (.Y(_05241_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .B(net2292));
 sg13g2_o21ai_1 _13193_ (.B1(_05241_),
    .Y(_05242_),
    .A1(_02043_),
    .A2(net2293));
 sg13g2_o21ai_1 _13194_ (.B1(net1876),
    .Y(_05243_),
    .A1(net2361),
    .A2(_05242_));
 sg13g2_a21oi_1 _13195_ (.A1(net2361),
    .A2(_05240_),
    .Y(_05244_),
    .B1(_05243_));
 sg13g2_nand2_1 _13196_ (.Y(_05245_),
    .A(_03627_),
    .B(net1864));
 sg13g2_o21ai_1 _13197_ (.B1(_05245_),
    .Y(_05246_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .A2(net1864));
 sg13g2_o21ai_1 _13198_ (.B1(net1844),
    .Y(_05247_),
    .A1(net1876),
    .A2(_05246_));
 sg13g2_o21ai_1 _13199_ (.B1(net2494),
    .Y(_05248_),
    .A1(_05244_),
    .A2(_05247_));
 sg13g2_a21oi_1 _13200_ (.A1(_01969_),
    .A2(net1848),
    .Y(_00614_),
    .B1(_05248_));
 sg13g2_a21o_1 _13201_ (.A2(_05239_),
    .A1(_05237_),
    .B1(_05236_),
    .X(_05249_));
 sg13g2_nor2_1 _13202_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(\i_tinyqv.cpu.imm[22] ),
    .Y(_05250_));
 sg13g2_xnor2_1 _13203_ (.Y(_05251_),
    .A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(\i_tinyqv.cpu.imm[22] ));
 sg13g2_xnor2_1 _13204_ (.Y(_05252_),
    .A(_05249_),
    .B(_05251_));
 sg13g2_nand2_1 _13205_ (.Y(_05253_),
    .A(_02044_),
    .B(net2296));
 sg13g2_o21ai_1 _13206_ (.B1(_05253_),
    .Y(_05254_),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A2(net2296));
 sg13g2_o21ai_1 _13207_ (.B1(net1876),
    .Y(_05255_),
    .A1(net2361),
    .A2(_05254_));
 sg13g2_a21oi_1 _13208_ (.A1(net2362),
    .A2(_05252_),
    .Y(_05256_),
    .B1(_05255_));
 sg13g2_nor2_1 _13209_ (.A(_03751_),
    .B(net1869),
    .Y(_05257_));
 sg13g2_a221oi_1 _13210_ (.B2(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .C1(_05257_),
    .B1(net1869),
    .A1(net2317),
    .Y(_05258_),
    .A2(_04573_));
 sg13g2_o21ai_1 _13211_ (.B1(net1844),
    .Y(_05259_),
    .A1(_05256_),
    .A2(_05258_));
 sg13g2_o21ai_1 _13212_ (.B1(_05259_),
    .Y(_05260_),
    .A1(net5259),
    .A2(net1844));
 sg13g2_nor2_1 _13213_ (.A(net2443),
    .B(_05260_),
    .Y(_00615_));
 sg13g2_a21oi_1 _13214_ (.A1(\i_tinyqv.cpu.instr_data_start[22] ),
    .A2(\i_tinyqv.cpu.imm[22] ),
    .Y(_05261_),
    .B1(_05249_));
 sg13g2_or2_1 _13215_ (.X(_05262_),
    .B(_05261_),
    .A(_05250_));
 sg13g2_xor2_1 _13216_ (.B(net4835),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .X(_05263_));
 sg13g2_xnor2_1 _13217_ (.Y(_05264_),
    .A(_05262_),
    .B(_05263_));
 sg13g2_nor2_1 _13218_ (.A(_02045_),
    .B(net2292),
    .Y(_05265_));
 sg13g2_a21oi_2 _13219_ (.B1(_05265_),
    .Y(_05266_),
    .A2(net2292),
    .A1(net4811));
 sg13g2_and2_1 _13220_ (.A(net2358),
    .B(_05266_),
    .X(_05267_));
 sg13g2_nor2b_1 _13221_ (.A(_05267_),
    .B_N(net1876),
    .Y(_05268_));
 sg13g2_o21ai_1 _13222_ (.B1(_05268_),
    .Y(_05269_),
    .A1(net2358),
    .A2(_05264_));
 sg13g2_nand2b_1 _13223_ (.Y(_05270_),
    .B(net1867),
    .A_N(net3402));
 sg13g2_a21oi_1 _13224_ (.A1(_03881_),
    .A2(net1864),
    .Y(_05271_),
    .B1(net1878));
 sg13g2_a21oi_1 _13225_ (.A1(_05270_),
    .A2(_05271_),
    .Y(_05272_),
    .B1(net1848));
 sg13g2_o21ai_1 _13226_ (.B1(net2494),
    .Y(_05273_),
    .A1(net5192),
    .A2(net1844));
 sg13g2_a21oi_1 _13227_ (.A1(_05269_),
    .A2(_05272_),
    .Y(_00616_),
    .B1(_05273_));
 sg13g2_a21o_1 _13228_ (.A2(_02021_),
    .A1(net5111),
    .B1(net5269),
    .X(_05274_));
 sg13g2_a22oi_1 _13229_ (.Y(_05275_),
    .B1(_04724_),
    .B2(net5270),
    .A2(net1882),
    .A1(net2564));
 sg13g2_nor2_1 _13230_ (.A(net2444),
    .B(net5271),
    .Y(_00617_));
 sg13g2_nand2_2 _13231_ (.Y(_05276_),
    .A(net2500),
    .B(net2315));
 sg13g2_o21ai_1 _13232_ (.B1(_04722_),
    .Y(_00618_),
    .A1(net2441),
    .A2(_05276_));
 sg13g2_nor2_2 _13233_ (.A(net2318),
    .B(_02808_),
    .Y(_05277_));
 sg13g2_nand2_2 _13234_ (.Y(_05278_),
    .A(_02730_),
    .B(_03415_));
 sg13g2_inv_1 _13235_ (.Y(_05279_),
    .A(_05278_));
 sg13g2_o21ai_1 _13236_ (.B1(net2501),
    .Y(_05280_),
    .A1(net2559),
    .A2(_05277_));
 sg13g2_a21oi_1 _13237_ (.A1(_05277_),
    .A2(_05278_),
    .Y(_00619_),
    .B1(_05280_));
 sg13g2_nand2_2 _13238_ (.Y(_05281_),
    .A(_02683_),
    .B(_03415_));
 sg13g2_inv_1 _13239_ (.Y(_05282_),
    .A(_05281_));
 sg13g2_o21ai_1 _13240_ (.B1(net2501),
    .Y(_05283_),
    .A1(net2557),
    .A2(_05277_));
 sg13g2_a21oi_1 _13241_ (.A1(_05277_),
    .A2(_05281_),
    .Y(_00620_),
    .B1(_05283_));
 sg13g2_nand2_2 _13242_ (.Y(_05284_),
    .A(_02652_),
    .B(_03415_));
 sg13g2_inv_1 _13243_ (.Y(_05285_),
    .A(_05284_));
 sg13g2_o21ai_1 _13244_ (.B1(net2502),
    .Y(_05286_),
    .A1(net2556),
    .A2(_05277_));
 sg13g2_a21oi_1 _13245_ (.A1(_05277_),
    .A2(_05284_),
    .Y(_00621_),
    .B1(_05286_));
 sg13g2_and2_1 _13246_ (.A(_02604_),
    .B(_03415_),
    .X(_05287_));
 sg13g2_inv_2 _13247_ (.Y(_05288_),
    .A(_05287_));
 sg13g2_o21ai_1 _13248_ (.B1(net2502),
    .Y(_05289_),
    .A1(net2555),
    .A2(_05277_));
 sg13g2_a21oi_1 _13249_ (.A1(_05277_),
    .A2(_05288_),
    .Y(_00622_),
    .B1(_05289_));
 sg13g2_and3_2 _13250_ (.X(_05290_),
    .A(net2318),
    .B(net2357),
    .C(_03386_));
 sg13g2_nor2_1 _13251_ (.A(net2366),
    .B(_05278_),
    .Y(_05291_));
 sg13g2_nand2_2 _13252_ (.Y(_05292_),
    .A(net2322),
    .B(net2357));
 sg13g2_a22oi_1 _13253_ (.Y(_05293_),
    .B1(_05292_),
    .B2(net2554),
    .A2(_05291_),
    .A1(net2226));
 sg13g2_nor2_1 _13254_ (.A(net2447),
    .B(_05293_),
    .Y(_00623_));
 sg13g2_nor2_1 _13255_ (.A(net2366),
    .B(_05281_),
    .Y(_05294_));
 sg13g2_a22oi_1 _13256_ (.Y(_05295_),
    .B1(_05294_),
    .B2(net2227),
    .A2(_05292_),
    .A1(net2553));
 sg13g2_nor2_1 _13257_ (.A(net2447),
    .B(_05295_),
    .Y(_00624_));
 sg13g2_nor2_1 _13258_ (.A(net2366),
    .B(_05284_),
    .Y(_05296_));
 sg13g2_a22oi_1 _13259_ (.Y(_05297_),
    .B1(_05296_),
    .B2(net2227),
    .A2(_05292_),
    .A1(net2552));
 sg13g2_nor2_1 _13260_ (.A(net2447),
    .B(_05297_),
    .Y(_00625_));
 sg13g2_nor2_1 _13261_ (.A(net2366),
    .B(_05288_),
    .Y(_05298_));
 sg13g2_a22oi_1 _13262_ (.Y(_05299_),
    .B1(_05298_),
    .B2(net2226),
    .A2(_05292_),
    .A1(net2551));
 sg13g2_nor2_1 _13263_ (.A(net2447),
    .B(_05299_),
    .Y(_00626_));
 sg13g2_nor2_1 _13264_ (.A(net2380),
    .B(_05278_),
    .Y(_05300_));
 sg13g2_nand2_2 _13265_ (.Y(_05301_),
    .A(_02619_),
    .B(net2357));
 sg13g2_a22oi_1 _13266_ (.Y(_05302_),
    .B1(_05301_),
    .B2(net2549),
    .A2(_05300_),
    .A1(net2227));
 sg13g2_nor2_1 _13267_ (.A(net2449),
    .B(_05302_),
    .Y(_00627_));
 sg13g2_nor2_1 _13268_ (.A(net2379),
    .B(_05281_),
    .Y(_05303_));
 sg13g2_a22oi_1 _13269_ (.Y(_05304_),
    .B1(_05303_),
    .B2(net2227),
    .A2(_05301_),
    .A1(net2548));
 sg13g2_nor2_1 _13270_ (.A(net2447),
    .B(_05304_),
    .Y(_00628_));
 sg13g2_nor2_1 _13271_ (.A(net2379),
    .B(_05284_),
    .Y(_05305_));
 sg13g2_a22oi_1 _13272_ (.Y(_05306_),
    .B1(_05305_),
    .B2(net2226),
    .A2(_05301_),
    .A1(net4958));
 sg13g2_nor2_1 _13273_ (.A(net2449),
    .B(_05306_),
    .Y(_00629_));
 sg13g2_nor2_1 _13274_ (.A(net2380),
    .B(_05288_),
    .Y(_05307_));
 sg13g2_a22oi_1 _13275_ (.Y(_05308_),
    .B1(_05307_),
    .B2(net2226),
    .A2(_05301_),
    .A1(net5104));
 sg13g2_nor2_1 _13276_ (.A(net2447),
    .B(_05308_),
    .Y(_00630_));
 sg13g2_nor2_1 _13277_ (.A(net2370),
    .B(_05278_),
    .Y(_05309_));
 sg13g2_nand2_2 _13278_ (.Y(_05310_),
    .A(_02705_),
    .B(_02807_));
 sg13g2_a22oi_1 _13279_ (.Y(_05311_),
    .B1(_05310_),
    .B2(net2547),
    .A2(_05309_),
    .A1(net2226));
 sg13g2_nor2_1 _13280_ (.A(net2446),
    .B(_05311_),
    .Y(_00631_));
 sg13g2_nor2_1 _13281_ (.A(net2370),
    .B(_05281_),
    .Y(_05312_));
 sg13g2_a22oi_1 _13282_ (.Y(_05313_),
    .B1(_05312_),
    .B2(net2226),
    .A2(_05310_),
    .A1(net5053));
 sg13g2_nor2_1 _13283_ (.A(net2446),
    .B(_05313_),
    .Y(_00632_));
 sg13g2_nor2_1 _13284_ (.A(net2370),
    .B(_05284_),
    .Y(_05314_));
 sg13g2_a22oi_1 _13285_ (.Y(_05315_),
    .B1(_05314_),
    .B2(net2226),
    .A2(_05310_),
    .A1(net4962));
 sg13g2_nor2_1 _13286_ (.A(net2446),
    .B(_05315_),
    .Y(_00633_));
 sg13g2_nor2_1 _13287_ (.A(net2370),
    .B(_05288_),
    .Y(_05316_));
 sg13g2_a22oi_1 _13288_ (.Y(_05317_),
    .B1(_05316_),
    .B2(net2226),
    .A2(_05310_),
    .A1(net4979));
 sg13g2_nor2_1 _13289_ (.A(net2446),
    .B(_05317_),
    .Y(_00634_));
 sg13g2_nand2_2 _13290_ (.Y(_05318_),
    .A(net2324),
    .B(net2357));
 sg13g2_o21ai_1 _13291_ (.B1(net2502),
    .Y(_05319_),
    .A1(_05279_),
    .A2(_05318_));
 sg13g2_a21oi_1 _13292_ (.A1(_01842_),
    .A2(_05318_),
    .Y(_00635_),
    .B1(_05319_));
 sg13g2_o21ai_1 _13293_ (.B1(net2502),
    .Y(_05320_),
    .A1(_05282_),
    .A2(_05318_));
 sg13g2_a21oi_1 _13294_ (.A1(_01840_),
    .A2(_05318_),
    .Y(_00636_),
    .B1(_05320_));
 sg13g2_o21ai_1 _13295_ (.B1(net2502),
    .Y(_05321_),
    .A1(_05285_),
    .A2(_05318_));
 sg13g2_a21oi_1 _13296_ (.A1(_01838_),
    .A2(_05318_),
    .Y(_00637_),
    .B1(_05321_));
 sg13g2_o21ai_1 _13297_ (.B1(net2502),
    .Y(_05322_),
    .A1(_05287_),
    .A2(_05318_));
 sg13g2_a21oi_1 _13298_ (.A1(_01836_),
    .A2(_05318_),
    .Y(_00638_),
    .B1(_05322_));
 sg13g2_a21oi_1 _13299_ (.A1(net2319),
    .A2(_03386_),
    .Y(_05323_),
    .B1(_02808_));
 sg13g2_nand2_2 _13300_ (.Y(_05324_),
    .A(_02550_),
    .B(net2357));
 sg13g2_a22oi_1 _13301_ (.Y(_05325_),
    .B1(_05324_),
    .B2(net4994),
    .A2(net2224),
    .A1(_05291_));
 sg13g2_nor2_1 _13302_ (.A(net2448),
    .B(_05325_),
    .Y(_00639_));
 sg13g2_a22oi_1 _13303_ (.Y(_05326_),
    .B1(_05324_),
    .B2(net4933),
    .A2(net2224),
    .A1(_05294_));
 sg13g2_nor2_1 _13304_ (.A(net2447),
    .B(_05326_),
    .Y(_00640_));
 sg13g2_a22oi_1 _13305_ (.Y(_05327_),
    .B1(_05324_),
    .B2(net4905),
    .A2(net2225),
    .A1(_05296_));
 sg13g2_nor2_1 _13306_ (.A(net2448),
    .B(_05327_),
    .Y(_00641_));
 sg13g2_a22oi_1 _13307_ (.Y(_05328_),
    .B1(_05324_),
    .B2(net4928),
    .A2(net2225),
    .A1(_05298_));
 sg13g2_nor2_1 _13308_ (.A(net2448),
    .B(_05328_),
    .Y(_00642_));
 sg13g2_nand2b_2 _13309_ (.Y(_05329_),
    .B(net2357),
    .A_N(_02524_));
 sg13g2_a22oi_1 _13310_ (.Y(_05330_),
    .B1(_05329_),
    .B2(net4986),
    .A2(net2225),
    .A1(_05300_));
 sg13g2_nor2_1 _13311_ (.A(net2448),
    .B(_05330_),
    .Y(_00643_));
 sg13g2_a22oi_1 _13312_ (.Y(_05331_),
    .B1(_05329_),
    .B2(net5071),
    .A2(net2225),
    .A1(_05303_));
 sg13g2_nor2_1 _13313_ (.A(net2449),
    .B(_05331_),
    .Y(_00644_));
 sg13g2_a22oi_1 _13314_ (.Y(_05332_),
    .B1(_05329_),
    .B2(net5054),
    .A2(net2224),
    .A1(_05305_));
 sg13g2_nor2_1 _13315_ (.A(net2449),
    .B(_05332_),
    .Y(_00645_));
 sg13g2_a22oi_1 _13316_ (.Y(_05333_),
    .B1(_05329_),
    .B2(net5079),
    .A2(net2224),
    .A1(_05307_));
 sg13g2_nor2_1 _13317_ (.A(net2447),
    .B(_05333_),
    .Y(_00646_));
 sg13g2_nand2_2 _13318_ (.Y(_05334_),
    .A(_02769_),
    .B(net2357));
 sg13g2_a22oi_1 _13319_ (.Y(_05335_),
    .B1(_05334_),
    .B2(net4927),
    .A2(net2224),
    .A1(_05309_));
 sg13g2_nor2_1 _13320_ (.A(net2446),
    .B(_05335_),
    .Y(_00647_));
 sg13g2_a22oi_1 _13321_ (.Y(_05336_),
    .B1(_05334_),
    .B2(net5055),
    .A2(net2224),
    .A1(_05312_));
 sg13g2_nor2_1 _13322_ (.A(net2448),
    .B(_05336_),
    .Y(_00648_));
 sg13g2_a22oi_1 _13323_ (.Y(_05337_),
    .B1(_05334_),
    .B2(net5005),
    .A2(net2224),
    .A1(_05314_));
 sg13g2_nor2_1 _13324_ (.A(net2446),
    .B(_05337_),
    .Y(_00649_));
 sg13g2_a22oi_1 _13325_ (.Y(_05338_),
    .B1(_05334_),
    .B2(net5020),
    .A2(net2224),
    .A1(_05316_));
 sg13g2_nor2_1 _13326_ (.A(net2451),
    .B(_05338_),
    .Y(_00650_));
 sg13g2_or2_1 _13327_ (.X(_05339_),
    .B(_03134_),
    .A(_02821_));
 sg13g2_nor2_1 _13328_ (.A(net5142),
    .B(_05339_),
    .Y(_05340_));
 sg13g2_nor2_1 _13329_ (.A(net4966),
    .B(_02819_),
    .Y(_05341_));
 sg13g2_o21ai_1 _13330_ (.B1(net2501),
    .Y(_00651_),
    .A1(_05340_),
    .A2(_05341_));
 sg13g2_nor2_1 _13331_ (.A(net5122),
    .B(_05339_),
    .Y(_05342_));
 sg13g2_nor2_1 _13332_ (.A(net4816),
    .B(_02819_),
    .Y(_05343_));
 sg13g2_o21ai_1 _13333_ (.B1(net2501),
    .Y(_00652_),
    .A1(_05342_),
    .A2(_05343_));
 sg13g2_a21oi_1 _13334_ (.A1(net3860),
    .A2(_03134_),
    .Y(_05344_),
    .B1(_02828_));
 sg13g2_nand2b_1 _13335_ (.Y(_05345_),
    .B(net2240),
    .A_N(\i_tinyqv.cpu.i_core.mem_op[0] ));
 sg13g2_o21ai_1 _13336_ (.B1(_05345_),
    .Y(_05346_),
    .A1(net4920),
    .A2(net2241));
 sg13g2_nand2_1 _13337_ (.Y(_00653_),
    .A(_05344_),
    .B(net4921));
 sg13g2_nand2b_1 _13338_ (.Y(_05347_),
    .B(net2241),
    .A_N(net4816));
 sg13g2_o21ai_1 _13339_ (.B1(_05347_),
    .Y(_05348_),
    .A1(net4949),
    .A2(net2241));
 sg13g2_nand2_1 _13340_ (.Y(_00654_),
    .A(_05344_),
    .B(_05348_));
 sg13g2_a21oi_1 _13341_ (.A1(net5122),
    .A2(net5142),
    .Y(_05349_),
    .B1(_03134_));
 sg13g2_nor2_1 _13342_ (.A(net2315),
    .B(_05349_),
    .Y(_05350_));
 sg13g2_a22oi_1 _13343_ (.Y(_05351_),
    .B1(_02819_),
    .B2(_05350_),
    .A2(net2315),
    .A1(net5073));
 sg13g2_nand2_1 _13344_ (.Y(_00655_),
    .A(net2501),
    .B(_05351_));
 sg13g2_nor2_1 _13345_ (.A(net3860),
    .B(net2240),
    .Y(_05352_));
 sg13g2_nor2_1 _13346_ (.A(_02828_),
    .B(_05352_),
    .Y(_00656_));
 sg13g2_nor2_1 _13347_ (.A(net2543),
    .B(net2544),
    .Y(_05353_));
 sg13g2_nand2_2 _13348_ (.Y(_05354_),
    .A(net2545),
    .B(net2546));
 sg13g2_nor3_1 _13349_ (.A(net2543),
    .B(net2544),
    .C(_05354_),
    .Y(_05355_));
 sg13g2_and2_1 _13350_ (.A(\i_i2c_peri.cmd_pending ),
    .B(\i_i2c_peri.i_i2c.s_axis_cmd_ready_reg ),
    .X(_05356_));
 sg13g2_nand2_2 _13351_ (.Y(_05357_),
    .A(net4055),
    .B(net4783));
 sg13g2_xnor2_1 _13352_ (.Y(_05358_),
    .A(\i_i2c_peri.cmd_read_reg ),
    .B(\i_i2c_peri.cmd_write_m_reg ));
 sg13g2_or2_1 _13353_ (.X(_05359_),
    .B(_05358_),
    .A(_05357_));
 sg13g2_nor3_1 _13354_ (.A(net2543),
    .B(net2544),
    .C(net2545),
    .Y(_05360_));
 sg13g2_nand2_1 _13355_ (.Y(_05361_),
    .A(_01966_),
    .B(_05353_));
 sg13g2_nor3_1 _13356_ (.A(net2546),
    .B(_05359_),
    .C(_05361_),
    .Y(_05362_));
 sg13g2_nor2_2 _13357_ (.A(net2461),
    .B(net2462),
    .Y(_05363_));
 sg13g2_nor3_2 _13358_ (.A(net2461),
    .B(net2462),
    .C(net2464),
    .Y(_05364_));
 sg13g2_nand2b_2 _13359_ (.Y(_05365_),
    .B(_05363_),
    .A_N(net2464));
 sg13g2_nand2b_2 _13360_ (.Y(_05366_),
    .B(net2545),
    .A_N(net2546));
 sg13g2_nor2b_1 _13361_ (.A(net2543),
    .B_N(net2544),
    .Y(_05367_));
 sg13g2_nand2b_2 _13362_ (.Y(_05368_),
    .B(net4976),
    .A_N(\i_i2c_peri.i_i2c.state_reg[3] ));
 sg13g2_nand2_1 _13363_ (.Y(_05369_),
    .A(net2545),
    .B(_05367_));
 sg13g2_nor2_2 _13364_ (.A(_05366_),
    .B(_05368_),
    .Y(_05370_));
 sg13g2_nand3_1 _13365_ (.B(_01781_),
    .C(net5365),
    .A(net5093),
    .Y(_05371_));
 sg13g2_nor2_2 _13366_ (.A(_05354_),
    .B(_05368_),
    .Y(_05372_));
 sg13g2_a22oi_1 _13367_ (.Y(_05373_),
    .B1(_05371_),
    .B2(net2283),
    .A2(_05370_),
    .A1(_02016_));
 sg13g2_nand2_1 _13368_ (.Y(_05374_),
    .A(net2332),
    .B(_05373_));
 sg13g2_nor3_1 _13369_ (.A(net2545),
    .B(\i_i2c_peri.i_i2c.state_reg[0] ),
    .C(_05368_),
    .Y(_05375_));
 sg13g2_nand3b_1 _13370_ (.B(net3988),
    .C(_05356_),
    .Y(_05376_),
    .A_N(\i_i2c_peri.cmd_read_reg ));
 sg13g2_nor2_1 _13371_ (.A(net4903),
    .B(_05376_),
    .Y(_05377_));
 sg13g2_nand2_2 _13372_ (.Y(_05378_),
    .A(net5358),
    .B(_05360_));
 sg13g2_inv_1 _13373_ (.Y(_05379_),
    .A(_05378_));
 sg13g2_nor2_1 _13374_ (.A(net2507),
    .B(net2506),
    .Y(_05380_));
 sg13g2_nor3_2 _13375_ (.A(net2507),
    .B(net2506),
    .C(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .Y(_05381_));
 sg13g2_nor3_1 _13376_ (.A(net2506),
    .B(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .C(\i_i2c_peri.i_i2c.bit_count_reg[3] ),
    .Y(_05382_));
 sg13g2_and2_1 _13377_ (.A(_02023_),
    .B(_05381_),
    .X(_05383_));
 sg13g2_nand2_2 _13378_ (.Y(_05384_),
    .A(_02023_),
    .B(_05381_));
 sg13g2_nor2b_2 _13379_ (.A(net2544),
    .B_N(net2543),
    .Y(_05385_));
 sg13g2_nor2b_1 _13380_ (.A(net2546),
    .B_N(_05385_),
    .Y(_05386_));
 sg13g2_nand2b_2 _13381_ (.Y(_05387_),
    .B(_05385_),
    .A_N(net2546));
 sg13g2_nor2_1 _13382_ (.A(_01966_),
    .B(_05387_),
    .Y(_05388_));
 sg13g2_nand3_1 _13383_ (.B(_05383_),
    .C(net2222),
    .A(\i_i2c_peri.i_i2c.mode_stop_reg ),
    .Y(_05389_));
 sg13g2_and3_2 _13384_ (.X(_05390_),
    .A(_01966_),
    .B(net2546),
    .C(_05367_));
 sg13g2_and2_1 _13385_ (.A(_05384_),
    .B(_05390_),
    .X(_05391_));
 sg13g2_inv_1 _13386_ (.Y(_05392_),
    .A(_05391_));
 sg13g2_nor3_1 _13387_ (.A(net2545),
    .B(_05384_),
    .C(_05387_),
    .Y(_05393_));
 sg13g2_nor3_2 _13388_ (.A(net2543),
    .B(net2544),
    .C(_05366_),
    .Y(_05394_));
 sg13g2_inv_1 _13389_ (.Y(_05395_),
    .A(_05394_));
 sg13g2_nand2_1 _13390_ (.Y(_05396_),
    .A(_05377_),
    .B(_05394_));
 sg13g2_nor2b_1 _13391_ (.A(\i_i2c_peri.i_i2c.last_reg ),
    .B_N(\i_i2c_peri.i_i2c.mode_write_multiple_reg ),
    .Y(_05397_));
 sg13g2_nand2b_1 _13392_ (.Y(_05398_),
    .B(net5348),
    .A_N(_05397_));
 sg13g2_nand2_1 _13393_ (.Y(_05399_),
    .A(net2546),
    .B(_05385_));
 sg13g2_nor2_1 _13394_ (.A(net2545),
    .B(_05399_),
    .Y(_05400_));
 sg13g2_nand2_1 _13395_ (.Y(_05401_),
    .A(_05398_),
    .B(_05400_));
 sg13g2_nor2_1 _13396_ (.A(_05355_),
    .B(_05375_),
    .Y(_05402_));
 sg13g2_nor2_1 _13397_ (.A(_05362_),
    .B(_05391_),
    .Y(_05403_));
 sg13g2_nand4_1 _13398_ (.B(_05396_),
    .C(_05402_),
    .A(_05389_),
    .Y(_05404_),
    .D(_05403_));
 sg13g2_o21ai_1 _13399_ (.B1(_05401_),
    .Y(_05405_),
    .A1(_05377_),
    .A2(_05378_));
 sg13g2_nor4_1 _13400_ (.A(_05374_),
    .B(_05393_),
    .C(_05404_),
    .D(_05405_),
    .Y(_05406_));
 sg13g2_o21ai_1 _13401_ (.B1(net2619),
    .Y(_05407_),
    .A1(net2546),
    .A2(net2332));
 sg13g2_nor2_1 _13402_ (.A(_05406_),
    .B(_05407_),
    .Y(_00657_));
 sg13g2_nand2_1 _13403_ (.Y(_05408_),
    .A(_01785_),
    .B(\i_i2c_peri.i_i2c.addr_reg[3] ));
 sg13g2_xor2_1 _13404_ (.B(\i_i2c_peri.i_i2c.addr_reg[5] ),
    .A(\i_i2c_peri.cmd_addr_reg[5] ),
    .X(_05409_));
 sg13g2_xor2_1 _13405_ (.B(\i_i2c_peri.i_i2c.addr_reg[4] ),
    .A(\i_i2c_peri.cmd_addr_reg[4] ),
    .X(_05410_));
 sg13g2_xor2_1 _13406_ (.B(\i_i2c_peri.i_i2c.addr_reg[1] ),
    .A(\i_i2c_peri.cmd_addr_reg[1] ),
    .X(_05411_));
 sg13g2_nor2_1 _13407_ (.A(_01788_),
    .B(\i_i2c_peri.i_i2c.addr_reg[0] ),
    .Y(_05412_));
 sg13g2_a21oi_1 _13408_ (.A1(net4331),
    .A2(_02017_),
    .Y(_05413_),
    .B1(_05409_));
 sg13g2_o21ai_1 _13409_ (.B1(_05408_),
    .Y(_05414_),
    .A1(_01782_),
    .A2(\i_i2c_peri.i_i2c.addr_reg[6] ));
 sg13g2_a221oi_1 _13410_ (.B2(_01782_),
    .C1(_05414_),
    .B1(\i_i2c_peri.i_i2c.addr_reg[6] ),
    .A1(_01788_),
    .Y(_05415_),
    .A2(\i_i2c_peri.i_i2c.addr_reg[0] ));
 sg13g2_xnor2_1 _13411_ (.Y(_05416_),
    .A(\i_i2c_peri.cmd_addr_reg[2] ),
    .B(\i_i2c_peri.i_i2c.addr_reg[2] ));
 sg13g2_nor4_1 _13412_ (.A(\i_i2c_peri.cmd_start_reg ),
    .B(_05410_),
    .C(_05411_),
    .D(_05412_),
    .Y(_05417_));
 sg13g2_nand4_1 _13413_ (.B(_05415_),
    .C(_05416_),
    .A(_05413_),
    .Y(_05418_),
    .D(_05417_));
 sg13g2_nand2b_1 _13414_ (.Y(_05419_),
    .B(_05418_),
    .A_N(_05358_));
 sg13g2_nand2_1 _13415_ (.Y(_05420_),
    .A(net4977),
    .B(_05419_));
 sg13g2_o21ai_1 _13416_ (.B1(\i_i2c_peri.i_i2c.bus_active_reg ),
    .Y(_05421_),
    .A1(_05355_),
    .A2(_05362_));
 sg13g2_nor3_1 _13417_ (.A(_05365_),
    .B(_05370_),
    .C(net2222),
    .Y(_05422_));
 sg13g2_a22oi_1 _13418_ (.Y(_05423_),
    .B1(_05394_),
    .B2(_05357_),
    .A2(net2283),
    .A1(_05371_));
 sg13g2_nand2_1 _13419_ (.Y(_05424_),
    .A(_05383_),
    .B(_05390_));
 sg13g2_a22oi_1 _13420_ (.Y(_05425_),
    .B1(_05397_),
    .B2(_05400_),
    .A2(_05390_),
    .A1(_05383_));
 sg13g2_nand4_1 _13421_ (.B(_05422_),
    .C(_05423_),
    .A(_05421_),
    .Y(_05426_),
    .D(_05425_));
 sg13g2_nor3_1 _13422_ (.A(net4723),
    .B(_05378_),
    .C(_05418_),
    .Y(_05427_));
 sg13g2_nand2b_1 _13423_ (.Y(_05428_),
    .B(_05427_),
    .A_N(_05359_));
 sg13g2_nor2b_1 _13424_ (.A(_05426_),
    .B_N(_05428_),
    .Y(_05429_));
 sg13g2_a221oi_1 _13425_ (.B2(_05429_),
    .C1(net2413),
    .B1(_05420_),
    .A1(_01966_),
    .Y(_00658_),
    .A2(_05365_));
 sg13g2_nor2b_1 _13426_ (.A(_05375_),
    .B_N(\i_i2c_peri.i_i2c.bus_active_reg ),
    .Y(_05430_));
 sg13g2_or2_1 _13427_ (.X(_05431_),
    .B(_05430_),
    .A(_05402_));
 sg13g2_a221oi_1 _13428_ (.B2(_05361_),
    .C1(_05359_),
    .B1(_05402_),
    .A1(\i_i2c_peri.i_i2c.bus_active_reg ),
    .Y(_05432_),
    .A2(_05378_));
 sg13g2_inv_1 _13429_ (.Y(_05433_),
    .A(_05432_));
 sg13g2_o21ai_1 _13430_ (.B1(_05431_),
    .Y(_05434_),
    .A1(_05427_),
    .A2(_05433_));
 sg13g2_and2_1 _13431_ (.A(_05364_),
    .B(_05434_),
    .X(_05435_));
 sg13g2_a21o_1 _13432_ (.A2(_05400_),
    .A1(_05397_),
    .B1(_05390_),
    .X(_05436_));
 sg13g2_or3_1 _13433_ (.A(_05357_),
    .B(_05395_),
    .C(_05419_),
    .X(_05437_));
 sg13g2_o21ai_1 _13434_ (.B1(_05431_),
    .Y(_05438_),
    .A1(_05359_),
    .A2(_05378_));
 sg13g2_nor4_1 _13435_ (.A(_05374_),
    .B(_05435_),
    .C(_05436_),
    .D(_05438_),
    .Y(_05439_));
 sg13g2_o21ai_1 _13436_ (.B1(net2619),
    .Y(_05440_),
    .A1(net2544),
    .A2(net2332));
 sg13g2_a21oi_1 _13437_ (.A1(_05437_),
    .A2(_05439_),
    .Y(_00659_),
    .B1(_05440_));
 sg13g2_a21oi_1 _13438_ (.A1(_05359_),
    .A2(_05376_),
    .Y(_05441_),
    .B1(_05395_));
 sg13g2_a21oi_1 _13439_ (.A1(net4566),
    .A2(_05370_),
    .Y(_05442_),
    .B1(_05365_));
 sg13g2_nand2b_1 _13440_ (.Y(_05443_),
    .B(net2283),
    .A_N(_05371_));
 sg13g2_o21ai_1 _13441_ (.B1(_05386_),
    .Y(_05444_),
    .A1(_01966_),
    .A2(net5348));
 sg13g2_nand3_1 _13442_ (.B(_05443_),
    .C(_05444_),
    .A(_05442_),
    .Y(_05445_));
 sg13g2_a221oi_1 _13443_ (.B2(_05441_),
    .C1(_05445_),
    .B1(_05419_),
    .A1(_05384_),
    .Y(_05446_),
    .A2(net2222));
 sg13g2_o21ai_1 _13444_ (.B1(net2619),
    .Y(_05447_),
    .A1(net2543),
    .A2(net2332));
 sg13g2_nor2_1 _13445_ (.A(_05446_),
    .B(_05447_),
    .Y(_00660_));
 sg13g2_nor2_1 _13446_ (.A(net2446),
    .B(net2539),
    .Y(_00661_));
 sg13g2_nor3_1 _13447_ (.A(net2446),
    .B(net2378),
    .C(net2374),
    .Y(_00662_));
 sg13g2_a21oi_1 _13448_ (.A1(net2435),
    .A2(net2371),
    .Y(_00663_),
    .B1(_05276_));
 sg13g2_nor3_1 _13449_ (.A(net2449),
    .B(_03135_),
    .C(_03136_),
    .Y(_00664_));
 sg13g2_a221oi_1 _13450_ (.B2(net4951),
    .C1(net2449),
    .B1(net2242),
    .A1(net2437),
    .Y(_05448_),
    .A2(_02538_));
 sg13g2_o21ai_1 _13451_ (.B1(_05448_),
    .Y(_05449_),
    .A1(net4951),
    .A2(_03134_));
 sg13g2_inv_1 _13452_ (.Y(_00665_),
    .A(net4952));
 sg13g2_or2_1 _13453_ (.X(_05450_),
    .B(_04576_),
    .A(net1880));
 sg13g2_nand2_1 _13454_ (.Y(_05451_),
    .A(net1875),
    .B(_05450_));
 sg13g2_nor2b_2 _13455_ (.A(_04601_),
    .B_N(_05450_),
    .Y(_05452_));
 sg13g2_nor2_2 _13456_ (.A(_04601_),
    .B(_05451_),
    .Y(_05453_));
 sg13g2_nand2_1 _13457_ (.Y(_05454_),
    .A(net1875),
    .B(_05452_));
 sg13g2_nor2_2 _13458_ (.A(net2105),
    .B(net1840),
    .Y(_05455_));
 sg13g2_nor2_1 _13459_ (.A(_04586_),
    .B(_04611_),
    .Y(_05456_));
 sg13g2_and2_1 _13460_ (.A(net2171),
    .B(_05456_),
    .X(_05457_));
 sg13g2_nand2_1 _13461_ (.Y(_05458_),
    .A(net2171),
    .B(_05456_));
 sg13g2_nor2_1 _13462_ (.A(_04609_),
    .B(_05458_),
    .Y(_05459_));
 sg13g2_nor4_2 _13463_ (.A(net2171),
    .B(_04586_),
    .C(_04607_),
    .Y(_05460_),
    .D(net2167));
 sg13g2_a21oi_1 _13464_ (.A1(_04612_),
    .A2(_05460_),
    .Y(_05461_),
    .B1(_05459_));
 sg13g2_nor2_1 _13465_ (.A(net2171),
    .B(_04610_),
    .Y(_05462_));
 sg13g2_and2_1 _13466_ (.A(_04613_),
    .B(_05462_),
    .X(_05463_));
 sg13g2_mux4_1 _13467_ (.S0(net2287),
    .A0(\i_tinyqv.cpu.instr_data[1][11] ),
    .A1(\i_tinyqv.cpu.instr_data[0][11] ),
    .A2(\i_tinyqv.cpu.instr_data[3][11] ),
    .A3(\i_tinyqv.cpu.instr_data[2][11] ),
    .S1(net2235),
    .X(_05464_));
 sg13g2_inv_4 _13468_ (.A(_05464_),
    .Y(_05465_));
 sg13g2_a22oi_1 _13469_ (.Y(_05466_),
    .B1(_05463_),
    .B2(_05465_),
    .A2(_04630_),
    .A1(net2109));
 sg13g2_nand3_1 _13470_ (.B(_05461_),
    .C(_05466_),
    .A(net1842),
    .Y(_05467_));
 sg13g2_o21ai_1 _13471_ (.B1(_05467_),
    .Y(_05468_),
    .A1(net5326),
    .A2(net1842));
 sg13g2_nor2_1 _13472_ (.A(net2442),
    .B(_05468_),
    .Y(_00666_));
 sg13g2_and2_1 _13473_ (.A(_04612_),
    .B(_04713_),
    .X(_05469_));
 sg13g2_and2_1 _13474_ (.A(net2170),
    .B(net2168),
    .X(_05470_));
 sg13g2_nand2_2 _13475_ (.Y(_05471_),
    .A(_05469_),
    .B(_05470_));
 sg13g2_nor3_1 _13476_ (.A(_04634_),
    .B(_04636_),
    .C(_04644_),
    .Y(_05472_));
 sg13g2_nor2b_1 _13477_ (.A(_05471_),
    .B_N(_05472_),
    .Y(_05473_));
 sg13g2_nand3_1 _13478_ (.B(_05470_),
    .C(_05472_),
    .A(_05469_),
    .Y(_05474_));
 sg13g2_nor2b_1 _13479_ (.A(net2167),
    .B_N(_05469_),
    .Y(_05475_));
 sg13g2_a21oi_1 _13480_ (.A1(_04609_),
    .A2(_05456_),
    .Y(_05476_),
    .B1(_05475_));
 sg13g2_nor2_1 _13481_ (.A(_04610_),
    .B(_05458_),
    .Y(_05477_));
 sg13g2_nor2_1 _13482_ (.A(_05475_),
    .B(_05477_),
    .Y(_05478_));
 sg13g2_nand2_1 _13483_ (.Y(_05479_),
    .A(_05474_),
    .B(_05476_));
 sg13g2_and3_2 _13484_ (.X(_05480_),
    .A(_04609_),
    .B(_04611_),
    .C(_04713_));
 sg13g2_nand3_1 _13485_ (.B(_04611_),
    .C(_04713_),
    .A(_04609_),
    .Y(_05481_));
 sg13g2_and2_1 _13486_ (.A(net2159),
    .B(_05464_),
    .X(_05482_));
 sg13g2_and2_1 _13487_ (.A(net2056),
    .B(_05482_),
    .X(_05483_));
 sg13g2_nor2_1 _13488_ (.A(_05481_),
    .B(_05483_),
    .Y(_05484_));
 sg13g2_nand2_1 _13489_ (.Y(_05485_),
    .A(_04622_),
    .B(net2163));
 sg13g2_nor3_1 _13490_ (.A(net2103),
    .B(_04629_),
    .C(_05485_),
    .Y(_05486_));
 sg13g2_nor3_1 _13491_ (.A(_05479_),
    .B(_05484_),
    .C(_05486_),
    .Y(_05487_));
 sg13g2_o21ai_1 _13492_ (.B1(net2495),
    .Y(_05488_),
    .A1(net5029),
    .A2(net1842));
 sg13g2_a21oi_1 _13493_ (.A1(net1843),
    .A2(_05487_),
    .Y(_00667_),
    .B1(_05488_));
 sg13g2_nor2b_1 _13494_ (.A(net2165),
    .B_N(net2164),
    .Y(_05489_));
 sg13g2_nand2_1 _13495_ (.Y(_05490_),
    .A(net2163),
    .B(_05489_));
 sg13g2_nand3_1 _13496_ (.B(_04627_),
    .C(_05489_),
    .A(net2163),
    .Y(_05491_));
 sg13g2_inv_1 _13497_ (.Y(_05492_),
    .A(net2052));
 sg13g2_nor2_1 _13498_ (.A(net2166),
    .B(net2053),
    .Y(_05493_));
 sg13g2_a22oi_1 _13499_ (.Y(_05494_),
    .B1(_05455_),
    .B2(_05493_),
    .A2(net1840),
    .A1(net5119));
 sg13g2_nor2_1 _13500_ (.A(net2442),
    .B(_05494_),
    .Y(_00668_));
 sg13g2_nand2_1 _13501_ (.Y(_05495_),
    .A(_05463_),
    .B(_05464_));
 sg13g2_nand2_1 _13502_ (.Y(_05496_),
    .A(net2170),
    .B(_04613_));
 sg13g2_nand3_1 _13503_ (.B(_05495_),
    .C(_05496_),
    .A(net2103),
    .Y(_05497_));
 sg13g2_nand2_2 _13504_ (.Y(_05498_),
    .A(net2166),
    .B(_04624_));
 sg13g2_nor2_1 _13505_ (.A(net2161),
    .B(net2051),
    .Y(_05499_));
 sg13g2_o21ai_1 _13506_ (.B1(_05497_),
    .Y(_05500_),
    .A1(net2105),
    .A2(_05499_));
 sg13g2_o21ai_1 _13507_ (.B1(net2495),
    .Y(_05501_),
    .A1(net5112),
    .A2(net1842));
 sg13g2_a21oi_1 _13508_ (.A1(net1842),
    .A2(_05500_),
    .Y(_00669_),
    .B1(_05501_));
 sg13g2_nor3_1 _13509_ (.A(_04619_),
    .B(net2161),
    .C(_05485_),
    .Y(_05502_));
 sg13g2_nor3_1 _13510_ (.A(net2103),
    .B(net1840),
    .C(_05502_),
    .Y(_05503_));
 sg13g2_o21ai_1 _13511_ (.B1(net2103),
    .Y(_05504_),
    .A1(_04617_),
    .A2(_04630_));
 sg13g2_and2_1 _13512_ (.A(_05480_),
    .B(_05483_),
    .X(_05505_));
 sg13g2_nor2_2 _13513_ (.A(_04615_),
    .B(_04712_),
    .Y(_05506_));
 sg13g2_nor4_1 _13514_ (.A(net1840),
    .B(_05504_),
    .C(_05505_),
    .D(_05506_),
    .Y(_05507_));
 sg13g2_nor2_1 _13515_ (.A(net2442),
    .B(net1840),
    .Y(_05508_));
 sg13g2_o21ai_1 _13516_ (.B1(net2495),
    .Y(_05509_),
    .A1(net5185),
    .A2(net1842));
 sg13g2_nor3_1 _13517_ (.A(_05503_),
    .B(_05507_),
    .C(_05509_),
    .Y(_00670_));
 sg13g2_nor2_2 _13518_ (.A(_05471_),
    .B(_05472_),
    .Y(_05510_));
 sg13g2_nor2_2 _13519_ (.A(net2107),
    .B(net2052),
    .Y(_05511_));
 sg13g2_a21oi_1 _13520_ (.A1(_04618_),
    .A2(_05511_),
    .Y(_05512_),
    .B1(_05510_));
 sg13g2_o21ai_1 _13521_ (.B1(net2495),
    .Y(_05513_),
    .A1(net4985),
    .A2(net1843));
 sg13g2_a21oi_1 _13522_ (.A1(net1842),
    .A2(_05512_),
    .Y(_00671_),
    .B1(_05513_));
 sg13g2_nor2_2 _13523_ (.A(_04627_),
    .B(net2051),
    .Y(_05514_));
 sg13g2_nand3_1 _13524_ (.B(_04624_),
    .C(net2161),
    .A(net2166),
    .Y(_05515_));
 sg13g2_and3_2 _13525_ (.X(_05516_),
    .A(net2169),
    .B(_04611_),
    .C(_04713_));
 sg13g2_nand3_1 _13526_ (.B(_04611_),
    .C(_04713_),
    .A(net2170),
    .Y(_05517_));
 sg13g2_nand2_1 _13527_ (.Y(_05518_),
    .A(net4409),
    .B(net1841));
 sg13g2_a22oi_1 _13528_ (.Y(_05519_),
    .B1(_05516_),
    .B2(net1842),
    .A2(_05514_),
    .A1(_05455_));
 sg13g2_a21oi_1 _13529_ (.A1(_05518_),
    .A2(_05519_),
    .Y(_00672_),
    .B1(net2442));
 sg13g2_nand3b_1 _13530_ (.B(_04645_),
    .C(_05465_),
    .Y(_05520_),
    .A_N(_04637_));
 sg13g2_inv_1 _13531_ (.Y(_05521_),
    .A(_05520_));
 sg13g2_nor3_1 _13532_ (.A(_04631_),
    .B(net1840),
    .C(_05521_),
    .Y(_05522_));
 sg13g2_a21oi_1 _13533_ (.A1(net5214),
    .A2(net1840),
    .Y(_05523_),
    .B1(_05522_));
 sg13g2_nand3_1 _13534_ (.B(_05455_),
    .C(_05489_),
    .A(_04717_),
    .Y(_05524_));
 sg13g2_a21oi_1 _13535_ (.A1(_05523_),
    .A2(_05524_),
    .Y(_00673_),
    .B1(net2442));
 sg13g2_o21ai_1 _13536_ (.B1(net2500),
    .Y(_05525_),
    .A1(_04720_),
    .A2(net1841));
 sg13g2_a21oi_1 _13537_ (.A1(_01964_),
    .A2(net1841),
    .Y(_00674_),
    .B1(_05525_));
 sg13g2_nand2_2 _13538_ (.Y(_05526_),
    .A(_05478_),
    .B(_05481_));
 sg13g2_nand2_1 _13539_ (.Y(_05527_),
    .A(_04715_),
    .B(_05517_));
 sg13g2_or2_1 _13540_ (.X(_05528_),
    .B(_05527_),
    .A(_05526_));
 sg13g2_nand2_1 _13541_ (.Y(_05529_),
    .A(_04613_),
    .B(_05470_));
 sg13g2_nor2_2 _13542_ (.A(net2171),
    .B(_05529_),
    .Y(_05530_));
 sg13g2_or2_1 _13543_ (.X(_05531_),
    .B(_05529_),
    .A(net2172));
 sg13g2_and2_1 _13544_ (.A(_05456_),
    .B(_05462_),
    .X(_05532_));
 sg13g2_nor2_2 _13545_ (.A(_05530_),
    .B(_05532_),
    .Y(_05533_));
 sg13g2_o21ai_1 _13546_ (.B1(_05471_),
    .Y(_05534_),
    .A1(_04615_),
    .A2(_04711_));
 sg13g2_nor4_1 _13547_ (.A(_05457_),
    .B(_05460_),
    .C(_05463_),
    .D(_05534_),
    .Y(_05535_));
 sg13g2_nand2_1 _13548_ (.Y(_05536_),
    .A(_05533_),
    .B(_05535_));
 sg13g2_nor2_1 _13549_ (.A(_05528_),
    .B(_05536_),
    .Y(_05537_));
 sg13g2_nor3_1 _13550_ (.A(net2172),
    .B(_05528_),
    .C(_05536_),
    .Y(_05538_));
 sg13g2_nor3_1 _13551_ (.A(net2103),
    .B(_04716_),
    .C(_05485_),
    .Y(_05539_));
 sg13g2_nand2_1 _13552_ (.Y(_05540_),
    .A(_04616_),
    .B(_05521_));
 sg13g2_nor2_1 _13553_ (.A(_04631_),
    .B(_05520_),
    .Y(_05541_));
 sg13g2_nor3_1 _13554_ (.A(_05538_),
    .B(_05539_),
    .C(_05541_),
    .Y(_05542_));
 sg13g2_o21ai_1 _13555_ (.B1(net2495),
    .Y(_05543_),
    .A1(net5062),
    .A2(net1843));
 sg13g2_a21oi_1 _13556_ (.A1(net1843),
    .A2(_05542_),
    .Y(_00675_),
    .B1(_05543_));
 sg13g2_nor2_1 _13557_ (.A(net4770),
    .B(net1843),
    .Y(_05544_));
 sg13g2_nor3_1 _13558_ (.A(net2442),
    .B(_05455_),
    .C(_05544_),
    .Y(_00676_));
 sg13g2_nand2_1 _13559_ (.Y(_05545_),
    .A(net4838),
    .B(net1841));
 sg13g2_nand3b_1 _13560_ (.B(_05545_),
    .C(net2495),
    .Y(_00677_),
    .A_N(_05455_));
 sg13g2_nor2_2 _13561_ (.A(net2107),
    .B(_05492_),
    .Y(_05546_));
 sg13g2_nand2_1 _13562_ (.Y(_05547_),
    .A(net2109),
    .B(net2052));
 sg13g2_nand2_1 _13563_ (.Y(_05548_),
    .A(_04644_),
    .B(_05499_));
 sg13g2_mux4_1 _13564_ (.S0(net2236),
    .A0(\i_tinyqv.cpu.instr_data[1][4] ),
    .A1(\i_tinyqv.cpu.instr_data[3][4] ),
    .A2(\i_tinyqv.cpu.instr_data[2][4] ),
    .A3(\i_tinyqv.cpu.instr_data[0][4] ),
    .S1(net2290),
    .X(_05549_));
 sg13g2_nand3_1 _13565_ (.B(net2051),
    .C(_05549_),
    .A(_04719_),
    .Y(_05550_));
 sg13g2_nand2_1 _13566_ (.Y(_05551_),
    .A(_05548_),
    .B(_05550_));
 sg13g2_nand3b_1 _13567_ (.B(_05463_),
    .C(net2162),
    .Y(_05552_),
    .A_N(net2159));
 sg13g2_nor2_1 _13568_ (.A(net2056),
    .B(_05481_),
    .Y(_05553_));
 sg13g2_nand2_2 _13569_ (.Y(_05554_),
    .A(_05482_),
    .B(_05553_));
 sg13g2_nand2_1 _13570_ (.Y(_05555_),
    .A(net2055),
    .B(_05482_));
 sg13g2_a22oi_1 _13571_ (.Y(_05556_),
    .B1(net1958),
    .B2(_05551_),
    .A2(_05526_),
    .A1(net2164));
 sg13g2_nand4_1 _13572_ (.B(_05552_),
    .C(_05554_),
    .A(_05540_),
    .Y(_05557_),
    .D(_05556_));
 sg13g2_mux2_1 _13573_ (.A0(net5298),
    .A1(_05557_),
    .S(net1823),
    .X(_00678_));
 sg13g2_a21oi_1 _13574_ (.A1(net2166),
    .A2(_05463_),
    .Y(_05558_),
    .B1(_05537_));
 sg13g2_a21oi_1 _13575_ (.A1(_05554_),
    .A2(_05558_),
    .Y(_05559_),
    .B1(net2108));
 sg13g2_mux4_1 _13576_ (.S0(net2235),
    .A0(\i_tinyqv.cpu.instr_data[1][5] ),
    .A1(\i_tinyqv.cpu.instr_data[3][5] ),
    .A2(\i_tinyqv.cpu.instr_data[2][5] ),
    .A3(\i_tinyqv.cpu.instr_data[0][5] ),
    .S1(net2289),
    .X(_05560_));
 sg13g2_mux2_1 _13577_ (.A0(_04635_),
    .A1(_05560_),
    .S(net2051),
    .X(_05561_));
 sg13g2_nand2_1 _13578_ (.Y(_05562_),
    .A(net2104),
    .B(net2165));
 sg13g2_inv_1 _13579_ (.Y(_05563_),
    .A(_05562_));
 sg13g2_a221oi_1 _13580_ (.B2(_05528_),
    .C1(_05559_),
    .B1(_05563_),
    .A1(net1958),
    .Y(_05564_),
    .A2(_05561_));
 sg13g2_nor2_1 _13581_ (.A(net5235),
    .B(net1818),
    .Y(_05565_));
 sg13g2_a21oi_1 _13582_ (.A1(net1818),
    .A2(_05564_),
    .Y(_00679_),
    .B1(_05565_));
 sg13g2_nand2b_1 _13583_ (.Y(_05566_),
    .B(_05554_),
    .A_N(net2163));
 sg13g2_mux4_1 _13584_ (.S0(net2236),
    .A0(\i_tinyqv.cpu.instr_data[1][6] ),
    .A1(\i_tinyqv.cpu.instr_data[3][6] ),
    .A2(\i_tinyqv.cpu.instr_data[2][6] ),
    .A3(\i_tinyqv.cpu.instr_data[0][6] ),
    .S1(net2290),
    .X(_05567_));
 sg13g2_inv_1 _13585_ (.Y(_05568_),
    .A(_05567_));
 sg13g2_a21oi_1 _13586_ (.A1(_05498_),
    .A2(_05568_),
    .Y(_05569_),
    .B1(_05547_));
 sg13g2_o21ai_1 _13587_ (.B1(_05569_),
    .Y(_05570_),
    .A1(_04633_),
    .A2(net2051));
 sg13g2_o21ai_1 _13588_ (.B1(net2162),
    .Y(_05571_),
    .A1(_05460_),
    .A2(_05532_));
 sg13g2_nand2_2 _13589_ (.Y(_05572_),
    .A(net2169),
    .B(_05457_));
 sg13g2_nand2_2 _13590_ (.Y(_05573_),
    .A(net2103),
    .B(net2163));
 sg13g2_or2_1 _13591_ (.X(_05574_),
    .B(_05573_),
    .A(_05572_));
 sg13g2_nand2_2 _13592_ (.Y(_05575_),
    .A(net2169),
    .B(_04614_));
 sg13g2_inv_1 _13593_ (.Y(_05576_),
    .A(_05575_));
 sg13g2_a22oi_1 _13594_ (.Y(_05577_),
    .B1(_05576_),
    .B2(_04633_),
    .A2(_05566_),
    .A1(_05528_));
 sg13g2_nand4_1 _13595_ (.B(_05571_),
    .C(_05574_),
    .A(_05570_),
    .Y(_05578_),
    .D(_05577_));
 sg13g2_mux2_1 _13596_ (.A0(net5279),
    .A1(_05578_),
    .S(net1828),
    .X(_00680_));
 sg13g2_nand4_1 _13597_ (.B(_05476_),
    .C(_05481_),
    .A(_04715_),
    .Y(_05579_),
    .D(_05572_));
 sg13g2_nand2b_2 _13598_ (.Y(_05580_),
    .B(_05517_),
    .A_N(_05460_));
 sg13g2_o21ai_1 _13599_ (.B1(net2159),
    .Y(_05581_),
    .A1(_05576_),
    .A2(_05580_));
 sg13g2_mux4_1 _13600_ (.S0(net2235),
    .A0(\i_tinyqv.cpu.instr_data[1][7] ),
    .A1(\i_tinyqv.cpu.instr_data[3][7] ),
    .A2(\i_tinyqv.cpu.instr_data[2][7] ),
    .A3(\i_tinyqv.cpu.instr_data[0][7] ),
    .S1(net2289),
    .X(_05582_));
 sg13g2_mux2_1 _13601_ (.A0(net2159),
    .A1(_05582_),
    .S(net2051),
    .X(_05583_));
 sg13g2_a22oi_1 _13602_ (.Y(_05584_),
    .B1(_05583_),
    .B2(net1958),
    .A2(_05579_),
    .A1(net2166));
 sg13g2_nand4_1 _13603_ (.B(_05554_),
    .C(_05581_),
    .A(net1819),
    .Y(_05585_),
    .D(_05584_));
 sg13g2_o21ai_1 _13604_ (.B1(_05585_),
    .Y(_05586_),
    .A1(net5325),
    .A2(net1818));
 sg13g2_inv_1 _13605_ (.Y(_00681_),
    .A(_05586_));
 sg13g2_nand2_1 _13606_ (.Y(_05587_),
    .A(_04715_),
    .B(_05533_));
 sg13g2_nand2_1 _13607_ (.Y(_05588_),
    .A(_05533_),
    .B(_05575_));
 sg13g2_nand3_1 _13608_ (.B(_05533_),
    .C(_05575_),
    .A(_04715_),
    .Y(_05589_));
 sg13g2_or2_1 _13609_ (.X(_05590_),
    .B(_05589_),
    .A(_05580_));
 sg13g2_nand2_1 _13610_ (.Y(_05591_),
    .A(net2162),
    .B(_05473_));
 sg13g2_nor2_1 _13611_ (.A(_05459_),
    .B(_05526_),
    .Y(_05592_));
 sg13g2_a22oi_1 _13612_ (.Y(_05593_),
    .B1(_05591_),
    .B2(_05592_),
    .A2(_05554_),
    .A1(_04627_));
 sg13g2_mux4_1 _13613_ (.S0(net2236),
    .A0(\i_tinyqv.cpu.instr_data[1][8] ),
    .A1(\i_tinyqv.cpu.instr_data[3][8] ),
    .A2(\i_tinyqv.cpu.instr_data[2][8] ),
    .A3(\i_tinyqv.cpu.instr_data[0][8] ),
    .S1(net2290),
    .X(_05594_));
 sg13g2_nand2_1 _13614_ (.Y(_05595_),
    .A(net2051),
    .B(_05594_));
 sg13g2_o21ai_1 _13615_ (.B1(_05595_),
    .Y(_05596_),
    .A1(_05465_),
    .A2(net2051));
 sg13g2_a221oi_1 _13616_ (.B2(net1958),
    .C1(_05593_),
    .B1(_05596_),
    .A1(_05464_),
    .Y(_05597_),
    .A2(_05590_));
 sg13g2_nor2_1 _13617_ (.A(net5149),
    .B(net1818),
    .Y(_05598_));
 sg13g2_a21oi_1 _13618_ (.A1(net1818),
    .A2(_05597_),
    .Y(_00682_),
    .B1(_05598_));
 sg13g2_nor2_2 _13619_ (.A(_04712_),
    .B(_05458_),
    .Y(_05599_));
 sg13g2_nand2_2 _13620_ (.Y(_05600_),
    .A(_04711_),
    .B(_05457_));
 sg13g2_nand2_2 _13621_ (.Y(_05601_),
    .A(_05474_),
    .B(_05600_));
 sg13g2_o21ai_1 _13622_ (.B1(net2164),
    .Y(_05602_),
    .A1(_05527_),
    .A2(_05601_));
 sg13g2_nand2_1 _13623_ (.Y(_05603_),
    .A(_05572_),
    .B(_05575_));
 sg13g2_mux4_1 _13624_ (.S0(net2235),
    .A0(\i_tinyqv.cpu.instr_data[1][9] ),
    .A1(\i_tinyqv.cpu.instr_data[3][9] ),
    .A2(\i_tinyqv.cpu.instr_data[2][9] ),
    .A3(\i_tinyqv.cpu.instr_data[0][9] ),
    .S1(net2289),
    .X(_05604_));
 sg13g2_nor4_1 _13625_ (.A(_05460_),
    .B(_05526_),
    .C(_05532_),
    .D(_05603_),
    .Y(_05605_));
 sg13g2_o21ai_1 _13626_ (.B1(_05602_),
    .Y(_05606_),
    .A1(net2056),
    .A2(_05605_));
 sg13g2_a221oi_1 _13627_ (.B2(_05604_),
    .C1(_05606_),
    .B1(net1958),
    .A1(net2159),
    .Y(_05607_),
    .A2(_05530_));
 sg13g2_nor2_1 _13628_ (.A(net5128),
    .B(net1826),
    .Y(_05608_));
 sg13g2_a21oi_1 _13629_ (.A1(net1826),
    .A2(_05607_),
    .Y(_00683_),
    .B1(_05608_));
 sg13g2_o21ai_1 _13630_ (.B1(net2166),
    .Y(_05609_),
    .A1(_05580_),
    .A2(_05601_));
 sg13g2_nand2_1 _13631_ (.Y(_05610_),
    .A(_04644_),
    .B(_05589_));
 sg13g2_nor2b_1 _13632_ (.A(_05572_),
    .B_N(net2164),
    .Y(_05611_));
 sg13g2_mux4_1 _13633_ (.S0(net2236),
    .A0(\i_tinyqv.cpu.instr_data[1][10] ),
    .A1(\i_tinyqv.cpu.instr_data[3][10] ),
    .A2(\i_tinyqv.cpu.instr_data[2][10] ),
    .A3(\i_tinyqv.cpu.instr_data[0][10] ),
    .S1(net2290),
    .X(_05612_));
 sg13g2_a221oi_1 _13634_ (.B2(_05612_),
    .C1(_05611_),
    .B1(net1958),
    .A1(net2055),
    .Y(_05613_),
    .A2(_05526_));
 sg13g2_nand4_1 _13635_ (.B(_05609_),
    .C(_05610_),
    .A(net1819),
    .Y(_05614_),
    .D(_05613_));
 sg13g2_o21ai_1 _13636_ (.B1(_05614_),
    .Y(_05615_),
    .A1(net5324),
    .A2(net1818));
 sg13g2_inv_1 _13637_ (.Y(_00684_),
    .A(_05615_));
 sg13g2_o21ai_1 _13638_ (.B1(net2165),
    .Y(_05616_),
    .A1(_05459_),
    .A2(_05473_));
 sg13g2_mux4_1 _13639_ (.S0(net2235),
    .A0(\i_tinyqv.cpu.instr_data[1][11] ),
    .A1(\i_tinyqv.cpu.instr_data[3][11] ),
    .A2(\i_tinyqv.cpu.instr_data[2][11] ),
    .A3(\i_tinyqv.cpu.instr_data[0][11] ),
    .S1(net2289),
    .X(_05617_));
 sg13g2_a22oi_1 _13640_ (.Y(_05618_),
    .B1(_05527_),
    .B2(net2161),
    .A2(_05526_),
    .A1(net2055));
 sg13g2_a22oi_1 _13641_ (.Y(_05619_),
    .B1(_05617_),
    .B2(net1958),
    .A2(_05588_),
    .A1(_04635_));
 sg13g2_nand4_1 _13642_ (.B(_05616_),
    .C(_05618_),
    .A(net1819),
    .Y(_05620_),
    .D(_05619_));
 sg13g2_o21ai_1 _13643_ (.B1(_05620_),
    .Y(_05621_),
    .A1(net5308),
    .A2(net1819));
 sg13g2_inv_1 _13644_ (.Y(_00685_),
    .A(_05621_));
 sg13g2_mux4_1 _13645_ (.S0(net2235),
    .A0(\i_tinyqv.cpu.instr_data[1][12] ),
    .A1(\i_tinyqv.cpu.instr_data[3][12] ),
    .A2(\i_tinyqv.cpu.instr_data[2][12] ),
    .A3(\i_tinyqv.cpu.instr_data[0][12] ),
    .S1(net2289),
    .X(_05622_));
 sg13g2_nand2_1 _13646_ (.Y(_05623_),
    .A(_05546_),
    .B(_05622_));
 sg13g2_nand2_1 _13647_ (.Y(_05624_),
    .A(_05482_),
    .B(_05490_));
 sg13g2_o21ai_1 _13648_ (.B1(_05553_),
    .Y(_05625_),
    .A1(net2165),
    .A2(_05624_));
 sg13g2_a21o_1 _13649_ (.A2(_05517_),
    .A1(_05478_),
    .B1(net2056),
    .X(_05626_));
 sg13g2_a22oi_1 _13650_ (.Y(_05627_),
    .B1(_05601_),
    .B2(_04623_),
    .A2(_05587_),
    .A1(_04633_));
 sg13g2_nand4_1 _13651_ (.B(_05625_),
    .C(_05626_),
    .A(_05623_),
    .Y(_05628_),
    .D(_05627_));
 sg13g2_mux2_1 _13652_ (.A0(net5337),
    .A1(_05628_),
    .S(net1819),
    .X(_00686_));
 sg13g2_o21ai_1 _13653_ (.B1(_05626_),
    .Y(_05629_),
    .A1(net2056),
    .A2(_05600_));
 sg13g2_nand2_1 _13654_ (.Y(_05630_),
    .A(_05474_),
    .B(_05531_));
 sg13g2_nand2_1 _13655_ (.Y(_05631_),
    .A(net2055),
    .B(_05630_));
 sg13g2_nand2_1 _13656_ (.Y(_05632_),
    .A(_05625_),
    .B(_05631_));
 sg13g2_nor2_1 _13657_ (.A(_05629_),
    .B(_05632_),
    .Y(_05633_));
 sg13g2_mux4_1 _13658_ (.S0(net2236),
    .A0(\i_tinyqv.cpu.instr_data[1][13] ),
    .A1(\i_tinyqv.cpu.instr_data[3][13] ),
    .A2(\i_tinyqv.cpu.instr_data[2][13] ),
    .A3(\i_tinyqv.cpu.instr_data[0][13] ),
    .S1(net2290),
    .X(_05634_));
 sg13g2_nand2_1 _13659_ (.Y(_05635_),
    .A(net2108),
    .B(_05634_));
 sg13g2_nand2b_1 _13660_ (.Y(_05636_),
    .B(net2052),
    .A_N(_05635_));
 sg13g2_o21ai_1 _13661_ (.B1(net2159),
    .Y(_05637_),
    .A1(_04714_),
    .A2(_05532_));
 sg13g2_nand4_1 _13662_ (.B(_05633_),
    .C(_05636_),
    .A(net1819),
    .Y(_05638_),
    .D(_05637_));
 sg13g2_o21ai_1 _13663_ (.B1(_05638_),
    .Y(_05639_),
    .A1(net5359),
    .A2(net1823));
 sg13g2_inv_1 _13664_ (.Y(_00687_),
    .A(_05639_));
 sg13g2_mux4_1 _13665_ (.S0(net2239),
    .A0(\i_tinyqv.cpu.instr_data[1][14] ),
    .A1(\i_tinyqv.cpu.instr_data[3][14] ),
    .A2(\i_tinyqv.cpu.instr_data[2][14] ),
    .A3(\i_tinyqv.cpu.instr_data[0][14] ),
    .S1(net2291),
    .X(_05640_));
 sg13g2_a22oi_1 _13666_ (.Y(_05641_),
    .B1(net1958),
    .B2(_05640_),
    .A2(_04714_),
    .A1(_04635_));
 sg13g2_nand3_1 _13667_ (.B(_05633_),
    .C(_05641_),
    .A(net1819),
    .Y(_05642_));
 sg13g2_o21ai_1 _13668_ (.B1(_05642_),
    .Y(_05643_),
    .A1(net2531),
    .A2(net1818));
 sg13g2_inv_1 _13669_ (.Y(_00688_),
    .A(_05643_));
 sg13g2_o21ai_1 _13670_ (.B1(_05633_),
    .Y(_05644_),
    .A1(_04642_),
    .A2(_04715_));
 sg13g2_mux4_1 _13671_ (.S0(net2238),
    .A0(\i_tinyqv.cpu.instr_data[1][15] ),
    .A1(\i_tinyqv.cpu.instr_data[3][15] ),
    .A2(\i_tinyqv.cpu.instr_data[2][15] ),
    .A3(\i_tinyqv.cpu.instr_data[0][15] ),
    .S1(net2291),
    .X(_05645_));
 sg13g2_and2_1 _13672_ (.A(_04719_),
    .B(_05645_),
    .X(_05646_));
 sg13g2_nand3_1 _13673_ (.B(_04718_),
    .C(_05549_),
    .A(_04620_),
    .Y(_05647_));
 sg13g2_nor2_1 _13674_ (.A(_05514_),
    .B(_05646_),
    .Y(_05648_));
 sg13g2_a221oi_1 _13675_ (.B2(_05648_),
    .C1(_05547_),
    .B1(_05647_),
    .A1(_04645_),
    .Y(_05649_),
    .A2(_05514_));
 sg13g2_o21ai_1 _13676_ (.B1(net1821),
    .Y(_05650_),
    .A1(_05644_),
    .A2(_05649_));
 sg13g2_o21ai_1 _13677_ (.B1(_05650_),
    .Y(_00689_),
    .A1(_01993_),
    .A2(net1826));
 sg13g2_nor2_1 _13678_ (.A(net4554),
    .B(net1826),
    .Y(_05651_));
 sg13g2_nand2_1 _13679_ (.Y(_05652_),
    .A(net2108),
    .B(_05645_));
 sg13g2_nand2_2 _13680_ (.Y(_05653_),
    .A(_04719_),
    .B(net2052));
 sg13g2_nand2_1 _13681_ (.Y(_05654_),
    .A(_05546_),
    .B(_05646_));
 sg13g2_nand2b_1 _13682_ (.Y(_05655_),
    .B(_05654_),
    .A_N(_05644_));
 sg13g2_nor2_1 _13683_ (.A(net2105),
    .B(net2056),
    .Y(_05656_));
 sg13g2_a221oi_1 _13684_ (.B2(_05656_),
    .C1(_05655_),
    .B1(_05653_),
    .A1(_04621_),
    .Y(_05657_),
    .A2(_05510_));
 sg13g2_a21oi_1 _13685_ (.A1(net1826),
    .A2(_05657_),
    .Y(_00690_),
    .B1(_05651_));
 sg13g2_nor2_1 _13686_ (.A(net4447),
    .B(net1825),
    .Y(_05658_));
 sg13g2_and2_1 _13687_ (.A(net2108),
    .B(net2168),
    .X(_05659_));
 sg13g2_a221oi_1 _13688_ (.B2(_05659_),
    .C1(_05655_),
    .B1(_05653_),
    .A1(_04620_),
    .Y(_05660_),
    .A2(_05510_));
 sg13g2_a21oi_1 _13689_ (.A1(net1825),
    .A2(_05660_),
    .Y(_00691_),
    .B1(_05658_));
 sg13g2_a21o_1 _13690_ (.A2(_05646_),
    .A1(net2052),
    .B1(net2107),
    .X(_05661_));
 sg13g2_a21oi_1 _13691_ (.A1(net2170),
    .A2(_05653_),
    .Y(_05662_),
    .B1(_05661_));
 sg13g2_a21oi_1 _13692_ (.A1(_04623_),
    .A2(_05510_),
    .Y(_05663_),
    .B1(_05644_));
 sg13g2_a21oi_1 _13693_ (.A1(net2107),
    .A2(_05663_),
    .Y(_05664_),
    .B1(_05662_));
 sg13g2_mux2_1 _13694_ (.A0(net4846),
    .A1(_05664_),
    .S(net1820),
    .X(_00692_));
 sg13g2_nor2_1 _13695_ (.A(net2104),
    .B(_04612_),
    .Y(_05665_));
 sg13g2_a221oi_1 _13696_ (.B2(_05665_),
    .C1(_05655_),
    .B1(_05653_),
    .A1(_04618_),
    .Y(_05666_),
    .A2(_05510_));
 sg13g2_nor2_1 _13697_ (.A(net4553),
    .B(net1825),
    .Y(_05667_));
 sg13g2_a21oi_1 _13698_ (.A1(net1825),
    .A2(_05666_),
    .Y(_00693_),
    .B1(_05667_));
 sg13g2_mux4_1 _13699_ (.S0(_04583_),
    .A0(\i_tinyqv.cpu.instr_data[0][0] ),
    .A1(\i_tinyqv.cpu.instr_data[2][0] ),
    .A2(\i_tinyqv.cpu.instr_data[3][0] ),
    .A3(\i_tinyqv.cpu.instr_data[1][0] ),
    .S1(net2288),
    .X(_05668_));
 sg13g2_a21oi_1 _13700_ (.A1(_05653_),
    .A2(_05668_),
    .Y(_05669_),
    .B1(_05661_));
 sg13g2_a22oi_1 _13701_ (.Y(_05670_),
    .B1(_05553_),
    .B2(_05624_),
    .A2(_04714_),
    .A1(net2055));
 sg13g2_nand2b_1 _13702_ (.Y(_05671_),
    .B(_05670_),
    .A_N(_05629_));
 sg13g2_a221oi_1 _13703_ (.B2(_04643_),
    .C1(_05671_),
    .B1(_05630_),
    .A1(net2161),
    .Y(_05672_),
    .A2(_05510_));
 sg13g2_a21oi_1 _13704_ (.A1(net2107),
    .A2(_05672_),
    .Y(_05673_),
    .B1(_05669_));
 sg13g2_mux2_1 _13705_ (.A0(net4858),
    .A1(_05673_),
    .S(net1821),
    .X(_00694_));
 sg13g2_nand2_1 _13706_ (.Y(_05674_),
    .A(_05471_),
    .B(_05531_));
 sg13g2_a21oi_1 _13707_ (.A1(_04643_),
    .A2(_05674_),
    .Y(_05675_),
    .B1(_05671_));
 sg13g2_nand2_1 _13708_ (.Y(_05676_),
    .A(_05654_),
    .B(_05675_));
 sg13g2_mux4_1 _13709_ (.S0(net2238),
    .A0(_02008_),
    .A1(_02010_),
    .A2(_02011_),
    .A3(_02009_),
    .S1(net2291),
    .X(_05677_));
 sg13g2_nor2_1 _13710_ (.A(_04588_),
    .B(_05677_),
    .Y(_05678_));
 sg13g2_a21oi_1 _13711_ (.A1(_05653_),
    .A2(_05678_),
    .Y(_05679_),
    .B1(_05676_));
 sg13g2_nor2_1 _13712_ (.A(net4472),
    .B(net1825),
    .Y(_05680_));
 sg13g2_a21oi_1 _13713_ (.A1(net1825),
    .A2(_05679_),
    .Y(_00695_),
    .B1(_05680_));
 sg13g2_mux4_1 _13714_ (.S0(_04583_),
    .A0(\i_tinyqv.cpu.instr_data[0][2] ),
    .A1(\i_tinyqv.cpu.instr_data[2][2] ),
    .A2(\i_tinyqv.cpu.instr_data[3][2] ),
    .A3(\i_tinyqv.cpu.instr_data[1][2] ),
    .S1(_04581_),
    .X(_05681_));
 sg13g2_and2_1 _13715_ (.A(net2108),
    .B(_05681_),
    .X(_05682_));
 sg13g2_a21oi_1 _13716_ (.A1(_05653_),
    .A2(_05682_),
    .Y(_05683_),
    .B1(_05676_));
 sg13g2_nor2_1 _13717_ (.A(net4406),
    .B(net1827),
    .Y(_05684_));
 sg13g2_a21oi_1 _13718_ (.A1(net1827),
    .A2(_05683_),
    .Y(_00696_),
    .B1(_05684_));
 sg13g2_mux4_1 _13719_ (.S0(_04583_),
    .A0(\i_tinyqv.cpu.instr_data[0][3] ),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .A2(\i_tinyqv.cpu.instr_data[3][3] ),
    .A3(\i_tinyqv.cpu.instr_data[1][3] ),
    .S1(net2288),
    .X(_05685_));
 sg13g2_nand3_1 _13720_ (.B(_05653_),
    .C(_05685_),
    .A(_04587_),
    .Y(_05686_));
 sg13g2_nor2b_1 _13721_ (.A(_05676_),
    .B_N(_05686_),
    .Y(_05687_));
 sg13g2_nor2_1 _13722_ (.A(net4533),
    .B(net1826),
    .Y(_05688_));
 sg13g2_a21oi_1 _13723_ (.A1(net1826),
    .A2(_05687_),
    .Y(_00697_),
    .B1(_05688_));
 sg13g2_a221oi_1 _13724_ (.B2(_04643_),
    .C1(_05671_),
    .B1(_05674_),
    .A1(_05546_),
    .Y(_05689_),
    .A2(_05645_));
 sg13g2_o21ai_1 _13725_ (.B1(_05675_),
    .Y(_05690_),
    .A1(_05492_),
    .A2(_05652_));
 sg13g2_nand2_1 _13726_ (.Y(_05691_),
    .A(net2109),
    .B(_05549_));
 sg13g2_o21ai_1 _13727_ (.B1(_05689_),
    .Y(_05692_),
    .A1(net2053),
    .A2(_05691_));
 sg13g2_mux2_1 _13728_ (.A0(net4746),
    .A1(_05692_),
    .S(net1824),
    .X(_00698_));
 sg13g2_nand2_1 _13729_ (.Y(_05693_),
    .A(net2108),
    .B(_05560_));
 sg13g2_o21ai_1 _13730_ (.B1(_05689_),
    .Y(_05694_),
    .A1(net2053),
    .A2(_05693_));
 sg13g2_mux2_1 _13731_ (.A0(net4831),
    .A1(_05694_),
    .S(net1824),
    .X(_00699_));
 sg13g2_nand2_1 _13732_ (.Y(_05695_),
    .A(net2108),
    .B(_05567_));
 sg13g2_o21ai_1 _13733_ (.B1(_05689_),
    .Y(_05696_),
    .A1(net2052),
    .A2(_05695_));
 sg13g2_mux2_1 _13734_ (.A0(net4932),
    .A1(_05696_),
    .S(net1826),
    .X(_00700_));
 sg13g2_nand2_1 _13735_ (.Y(_05697_),
    .A(net2108),
    .B(_05582_));
 sg13g2_o21ai_1 _13736_ (.B1(_05689_),
    .Y(_05698_),
    .A1(net2052),
    .A2(_05697_));
 sg13g2_mux2_1 _13737_ (.A0(net4835),
    .A1(_05698_),
    .S(net1821),
    .X(_00701_));
 sg13g2_a21oi_1 _13738_ (.A1(_05511_),
    .A2(_05594_),
    .Y(_05699_),
    .B1(_05690_));
 sg13g2_nor2_1 _13739_ (.A(net4287),
    .B(net1822),
    .Y(_05700_));
 sg13g2_a21oi_1 _13740_ (.A1(net1822),
    .A2(_05699_),
    .Y(_00702_),
    .B1(_05700_));
 sg13g2_a21oi_1 _13741_ (.A1(_05511_),
    .A2(_05604_),
    .Y(_05701_),
    .B1(_05690_));
 sg13g2_nor2_1 _13742_ (.A(net4361),
    .B(net1820),
    .Y(_05702_));
 sg13g2_a21oi_1 _13743_ (.A1(net1818),
    .A2(_05701_),
    .Y(_00703_),
    .B1(_05702_));
 sg13g2_a21oi_1 _13744_ (.A1(_05511_),
    .A2(_05612_),
    .Y(_05703_),
    .B1(_05690_));
 sg13g2_nor2_1 _13745_ (.A(net4376),
    .B(net1820),
    .Y(_05704_));
 sg13g2_a21oi_1 _13746_ (.A1(net1820),
    .A2(_05703_),
    .Y(_00704_),
    .B1(_05704_));
 sg13g2_a21oi_1 _13747_ (.A1(_05511_),
    .A2(_05617_),
    .Y(_05705_),
    .B1(_05690_));
 sg13g2_nor2_1 _13748_ (.A(net3843),
    .B(net1825),
    .Y(_05706_));
 sg13g2_a21oi_1 _13749_ (.A1(net1825),
    .A2(_05705_),
    .Y(_00705_),
    .B1(_05706_));
 sg13g2_a21oi_1 _13750_ (.A1(_05511_),
    .A2(_05622_),
    .Y(_05707_),
    .B1(_05690_));
 sg13g2_nor2_1 _13751_ (.A(net4291),
    .B(net1821),
    .Y(_05708_));
 sg13g2_a21oi_1 _13752_ (.A1(net1821),
    .A2(_05707_),
    .Y(_00706_),
    .B1(_05708_));
 sg13g2_o21ai_1 _13753_ (.B1(_05689_),
    .Y(_05709_),
    .A1(net2053),
    .A2(_05635_));
 sg13g2_mux2_1 _13754_ (.A0(net4257),
    .A1(_05709_),
    .S(net1821),
    .X(_00707_));
 sg13g2_a21oi_1 _13755_ (.A1(_05511_),
    .A2(_05640_),
    .Y(_05710_),
    .B1(_05690_));
 sg13g2_nor2_1 _13756_ (.A(net4515),
    .B(net1820),
    .Y(_05711_));
 sg13g2_a21oi_1 _13757_ (.A1(net1820),
    .A2(_05710_),
    .Y(_00708_),
    .B1(_05711_));
 sg13g2_nand3_1 _13758_ (.B(_05652_),
    .C(_05675_),
    .A(net1820),
    .Y(_05712_));
 sg13g2_o21ai_1 _13759_ (.B1(_05712_),
    .Y(_05713_),
    .A1(net4797),
    .A2(net1820));
 sg13g2_inv_1 _13760_ (.Y(_00709_),
    .A(_05713_));
 sg13g2_nand2_2 _13761_ (.Y(_05714_),
    .A(_05502_),
    .B(_05612_));
 sg13g2_nand2_1 _13762_ (.Y(_05715_),
    .A(_05515_),
    .B(_05714_));
 sg13g2_nor4_2 _13763_ (.A(net2103),
    .B(_04628_),
    .C(_04718_),
    .Y(_05716_),
    .D(_05493_));
 sg13g2_mux2_1 _13764_ (.A0(net2055),
    .A1(net2167),
    .S(_05715_),
    .X(_05717_));
 sg13g2_o21ai_1 _13765_ (.B1(_05480_),
    .Y(_05718_),
    .A1(_05490_),
    .A2(_05555_));
 sg13g2_a21oi_1 _13766_ (.A1(_04716_),
    .A2(_05483_),
    .Y(_05719_),
    .B1(_05718_));
 sg13g2_a21o_1 _13767_ (.A2(_05717_),
    .A1(_05716_),
    .B1(_05719_),
    .X(_05720_));
 sg13g2_o21ai_1 _13768_ (.B1(net1823),
    .Y(_05721_),
    .A1(_05477_),
    .A2(_05720_));
 sg13g2_o21ai_1 _13769_ (.B1(_05721_),
    .Y(_00710_),
    .A1(_02001_),
    .A2(net1829));
 sg13g2_nor2_1 _13770_ (.A(net2167),
    .B(_05715_),
    .Y(_05722_));
 sg13g2_nor2_1 _13771_ (.A(_05617_),
    .B(_05714_),
    .Y(_05723_));
 sg13g2_a21oi_1 _13772_ (.A1(_04607_),
    .A2(_05714_),
    .Y(_05724_),
    .B1(_05723_));
 sg13g2_o21ai_1 _13773_ (.B1(_05716_),
    .Y(_05725_),
    .A1(net2169),
    .A2(_05515_));
 sg13g2_nor2_1 _13774_ (.A(_05722_),
    .B(_05725_),
    .Y(_05726_));
 sg13g2_a21oi_1 _13775_ (.A1(_04627_),
    .A2(_05483_),
    .Y(_05727_),
    .B1(_05465_));
 sg13g2_nor2b_1 _13776_ (.A(_05718_),
    .B_N(_05727_),
    .Y(_05728_));
 sg13g2_nor3_1 _13777_ (.A(_05506_),
    .B(_05726_),
    .C(_05728_),
    .Y(_05729_));
 sg13g2_nor2_1 _13778_ (.A(net4352),
    .B(net1823),
    .Y(_05730_));
 sg13g2_a21oi_1 _13779_ (.A1(net1823),
    .A2(_05729_),
    .Y(_00711_),
    .B1(_05730_));
 sg13g2_nand2b_1 _13780_ (.Y(_05731_),
    .B(_05483_),
    .A_N(_04629_));
 sg13g2_xnor2_1 _13781_ (.Y(_05732_),
    .A(_05515_),
    .B(_05724_));
 sg13g2_a221oi_1 _13782_ (.B2(_05716_),
    .C1(_05516_),
    .B1(_05732_),
    .A1(_05480_),
    .Y(_05733_),
    .A2(_05731_));
 sg13g2_nor2_1 _13783_ (.A(net2526),
    .B(net1823),
    .Y(_05734_));
 sg13g2_a21oi_1 _13784_ (.A1(net1823),
    .A2(_05733_),
    .Y(_00712_),
    .B1(_05734_));
 sg13g2_o21ai_1 _13785_ (.B1(_04619_),
    .Y(_05735_),
    .A1(net2168),
    .A2(net2056));
 sg13g2_nand2_1 _13786_ (.Y(_05736_),
    .A(_05640_),
    .B(_05735_));
 sg13g2_a21oi_1 _13787_ (.A1(_05714_),
    .A2(_05736_),
    .Y(_05737_),
    .B1(_05514_));
 sg13g2_nand2_1 _13788_ (.Y(_05738_),
    .A(net2159),
    .B(_05465_));
 sg13g2_a21oi_1 _13789_ (.A1(_05731_),
    .A2(_05738_),
    .Y(_05739_),
    .B1(_05481_));
 sg13g2_a221oi_1 _13790_ (.B2(_05737_),
    .C1(_05739_),
    .B1(_05716_),
    .A1(_04614_),
    .Y(_05740_),
    .A2(_04711_));
 sg13g2_nor2_1 _13791_ (.A(net5189),
    .B(net1824),
    .Y(_05741_));
 sg13g2_a21oi_1 _13792_ (.A1(net1828),
    .A2(_05740_),
    .Y(_00713_),
    .B1(_05741_));
 sg13g2_nand3_1 _13793_ (.B(_04628_),
    .C(net2055),
    .A(net2168),
    .Y(_05742_));
 sg13g2_nand2_1 _13794_ (.Y(_05743_),
    .A(_05461_),
    .B(_05496_));
 sg13g2_nor2_1 _13795_ (.A(_05516_),
    .B(_05743_),
    .Y(_05744_));
 sg13g2_a22oi_1 _13796_ (.Y(_05745_),
    .B1(_05744_),
    .B2(net2160),
    .A2(_05516_),
    .A1(net2168));
 sg13g2_inv_1 _13797_ (.Y(_05746_),
    .A(_05745_));
 sg13g2_a22oi_1 _13798_ (.Y(_05747_),
    .B1(_05746_),
    .B2(net2105),
    .A2(_05742_),
    .A1(_05656_));
 sg13g2_nor2_1 _13799_ (.A(net4966),
    .B(net1829),
    .Y(_05748_));
 sg13g2_a21oi_1 _13800_ (.A1(net1829),
    .A2(_05747_),
    .Y(_00714_),
    .B1(_05748_));
 sg13g2_nor2_2 _13801_ (.A(_05659_),
    .B(_05743_),
    .Y(_05749_));
 sg13g2_nor2_1 _13802_ (.A(net4816),
    .B(net1829),
    .Y(_05750_));
 sg13g2_a21oi_1 _13803_ (.A1(net1829),
    .A2(_05749_),
    .Y(_00715_),
    .B1(_05750_));
 sg13g2_nand2_1 _13804_ (.Y(_05751_),
    .A(net2109),
    .B(net2170));
 sg13g2_nand3_1 _13805_ (.B(_05470_),
    .C(_05499_),
    .A(_04642_),
    .Y(_05752_));
 sg13g2_nand2_1 _13806_ (.Y(_05753_),
    .A(_05742_),
    .B(_05752_));
 sg13g2_a21oi_1 _13807_ (.A1(net2162),
    .A2(net2160),
    .Y(_05754_),
    .B1(_05464_));
 sg13g2_nand3_1 _13808_ (.B(_05744_),
    .C(_05754_),
    .A(net2105),
    .Y(_05755_));
 sg13g2_o21ai_1 _13809_ (.B1(_05755_),
    .Y(_05756_),
    .A1(_05751_),
    .A2(_05753_));
 sg13g2_mux2_1 _13810_ (.A0(net4338),
    .A1(_05756_),
    .S(net1829),
    .X(_00716_));
 sg13g2_nor2_1 _13811_ (.A(net5226),
    .B(net1824),
    .Y(_05757_));
 sg13g2_nand2_1 _13812_ (.Y(_05758_),
    .A(_04609_),
    .B(_05469_));
 sg13g2_a21o_2 _13813_ (.A2(_05462_),
    .A1(_04611_),
    .B1(_05580_),
    .X(_05759_));
 sg13g2_nor2_1 _13814_ (.A(_04617_),
    .B(net2056),
    .Y(_05760_));
 sg13g2_nor4_1 _13815_ (.A(_05477_),
    .B(_05506_),
    .C(_05759_),
    .D(_05760_),
    .Y(_05761_));
 sg13g2_nand3_1 _13816_ (.B(_05758_),
    .C(_05761_),
    .A(_04631_),
    .Y(_05762_));
 sg13g2_nand2_1 _13817_ (.Y(_05763_),
    .A(_05531_),
    .B(_05600_));
 sg13g2_a221oi_1 _13818_ (.B2(_05762_),
    .C1(_05763_),
    .B1(_04644_),
    .A1(net2109),
    .Y(_05764_),
    .A2(_04611_));
 sg13g2_a21oi_1 _13819_ (.A1(net1824),
    .A2(_05764_),
    .Y(_00717_),
    .B1(_05757_));
 sg13g2_nor2_1 _13820_ (.A(net2106),
    .B(_05668_),
    .Y(_05765_));
 sg13g2_nand2_1 _13821_ (.Y(_05766_),
    .A(_04635_),
    .B(_05762_));
 sg13g2_nand2_1 _13822_ (.Y(_05767_),
    .A(net2104),
    .B(_05471_));
 sg13g2_a21oi_1 _13823_ (.A1(_05572_),
    .A2(_05575_),
    .Y(_05768_),
    .B1(net2168));
 sg13g2_nor4_1 _13824_ (.A(_05532_),
    .B(_05763_),
    .C(_05767_),
    .D(_05768_),
    .Y(_05769_));
 sg13g2_a21oi_2 _13825_ (.B1(_05765_),
    .Y(_05770_),
    .A2(_05769_),
    .A1(_05766_));
 sg13g2_mux2_1 _13826_ (.A0(net5060),
    .A1(_05770_),
    .S(net1829),
    .X(_00718_));
 sg13g2_a22oi_1 _13827_ (.Y(_05771_),
    .B1(_05762_),
    .B2(_04633_),
    .A2(_05470_),
    .A1(net2173));
 sg13g2_nor2_1 _13828_ (.A(net2109),
    .B(_05771_),
    .Y(_05772_));
 sg13g2_or2_1 _13829_ (.X(_05773_),
    .B(_05772_),
    .A(_05678_));
 sg13g2_mux2_1 _13830_ (.A0(net5044),
    .A1(_05773_),
    .S(net1830),
    .X(_00719_));
 sg13g2_o21ai_1 _13831_ (.B1(net2103),
    .Y(_05774_),
    .A1(net2160),
    .A2(_05759_));
 sg13g2_inv_1 _13832_ (.Y(_05775_),
    .A(_05774_));
 sg13g2_a21oi_1 _13833_ (.A1(_05762_),
    .A2(_05775_),
    .Y(_05776_),
    .B1(_05682_));
 sg13g2_nor2_1 _13834_ (.A(net5250),
    .B(net1824),
    .Y(_05777_));
 sg13g2_a21oi_1 _13835_ (.A1(net1824),
    .A2(_05776_),
    .Y(_00720_),
    .B1(_05777_));
 sg13g2_a21oi_2 _13836_ (.B1(_05452_),
    .Y(_05778_),
    .A2(_02824_),
    .A1(_02814_));
 sg13g2_inv_4 _13837_ (.A(_05778_),
    .Y(_05779_));
 sg13g2_nand2_1 _13838_ (.Y(_05780_),
    .A(net2499),
    .B(_05779_));
 sg13g2_nand3_1 _13839_ (.B(net2164),
    .C(_05517_),
    .A(net2104),
    .Y(_05781_));
 sg13g2_xor2_1 _13840_ (.B(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A(net3944),
    .X(_05782_));
 sg13g2_nand4_1 _13841_ (.B(_05531_),
    .C(_05691_),
    .A(net1875),
    .Y(_05783_),
    .D(_05781_));
 sg13g2_o21ai_1 _13842_ (.B1(_05783_),
    .Y(_05784_),
    .A1(net1874),
    .A2(_05782_));
 sg13g2_nand2_1 _13843_ (.Y(_05785_),
    .A(net3944),
    .B(net1809));
 sg13g2_o21ai_1 _13844_ (.B1(_05785_),
    .Y(_00721_),
    .A1(net1809),
    .A2(_05784_));
 sg13g2_nand3_1 _13845_ (.B(net2517),
    .C(net4397),
    .A(net2515),
    .Y(_05786_));
 sg13g2_a21o_1 _13846_ (.A2(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A1(net2517),
    .B1(net2515),
    .X(_05787_));
 sg13g2_and2_1 _13847_ (.A(_05786_),
    .B(_05787_),
    .X(_05788_));
 sg13g2_nor3_1 _13848_ (.A(_04614_),
    .B(_05516_),
    .C(_05530_),
    .Y(_05789_));
 sg13g2_nor2_1 _13849_ (.A(net2172),
    .B(_05789_),
    .Y(_05790_));
 sg13g2_o21ai_1 _13850_ (.B1(_05693_),
    .Y(_05791_),
    .A1(_05562_),
    .A2(_05790_));
 sg13g2_mux2_1 _13851_ (.A0(_05788_),
    .A1(_05791_),
    .S(net1873),
    .X(_05792_));
 sg13g2_nor2_1 _13852_ (.A(net1809),
    .B(_05792_),
    .Y(_05793_));
 sg13g2_a21oi_1 _13853_ (.A1(_01995_),
    .A2(net1808),
    .Y(_00722_),
    .B1(_05793_));
 sg13g2_or2_1 _13854_ (.X(_05794_),
    .B(_05786_),
    .A(_01994_));
 sg13g2_xnor2_1 _13855_ (.Y(_05795_),
    .A(_01994_),
    .B(_05786_));
 sg13g2_o21ai_1 _13856_ (.B1(_05695_),
    .Y(_05796_),
    .A1(_05573_),
    .A2(_05790_));
 sg13g2_nor2_1 _13857_ (.A(net1873),
    .B(_05795_),
    .Y(_05797_));
 sg13g2_a21oi_1 _13858_ (.A1(net1873),
    .A2(_05796_),
    .Y(_05798_),
    .B1(_05797_));
 sg13g2_nand2_1 _13859_ (.Y(_05799_),
    .A(net2514),
    .B(net1808));
 sg13g2_o21ai_1 _13860_ (.B1(_05799_),
    .Y(_00723_),
    .A1(net1809),
    .A2(_05798_));
 sg13g2_a21oi_1 _13861_ (.A1(_04615_),
    .A2(_05529_),
    .Y(_05800_),
    .B1(_04619_));
 sg13g2_o21ai_1 _13862_ (.B1(net2104),
    .Y(_05801_),
    .A1(_05789_),
    .A2(_05800_));
 sg13g2_nand2_2 _13863_ (.Y(_05802_),
    .A(_05697_),
    .B(_05801_));
 sg13g2_xor2_1 _13864_ (.B(_05794_),
    .A(net2513),
    .X(_05803_));
 sg13g2_nor2_1 _13865_ (.A(net1874),
    .B(_05803_),
    .Y(_05804_));
 sg13g2_a21oi_1 _13866_ (.A1(net1873),
    .A2(_05802_),
    .Y(_05805_),
    .B1(_05804_));
 sg13g2_nand2_1 _13867_ (.Y(_05806_),
    .A(net2513),
    .B(net1808));
 sg13g2_o21ai_1 _13868_ (.B1(_05806_),
    .Y(_00724_),
    .A1(net1809),
    .A2(_05805_));
 sg13g2_a22oi_1 _13869_ (.Y(_05807_),
    .B1(_05599_),
    .B2(_04644_),
    .A2(_05530_),
    .A1(net2164));
 sg13g2_nand2_1 _13870_ (.Y(_05808_),
    .A(net2109),
    .B(_05753_));
 sg13g2_a21oi_1 _13871_ (.A1(_05807_),
    .A2(_05808_),
    .Y(_05809_),
    .B1(net1840));
 sg13g2_nand2_1 _13872_ (.Y(_05810_),
    .A(net5352),
    .B(_05778_));
 sg13g2_o21ai_1 _13873_ (.B1(_05810_),
    .Y(_05811_),
    .A1(net5352),
    .A2(net1875));
 sg13g2_o21ai_1 _13874_ (.B1(net2495),
    .Y(_05812_),
    .A1(_05809_),
    .A2(_05811_));
 sg13g2_inv_1 _13875_ (.Y(_00725_),
    .A(_05812_));
 sg13g2_xnor2_1 _13876_ (.Y(_05813_),
    .A(net5050),
    .B(\i_tinyqv.cpu.additional_mem_ops[0] ));
 sg13g2_nor2_2 _13877_ (.A(net2105),
    .B(_05752_),
    .Y(_05814_));
 sg13g2_a221oi_1 _13878_ (.B2(_04635_),
    .C1(_05814_),
    .B1(_05599_),
    .A1(net2165),
    .Y(_05815_),
    .A2(_05530_));
 sg13g2_o21ai_1 _13879_ (.B1(_05815_),
    .Y(_05816_),
    .A1(_05742_),
    .A2(_05751_));
 sg13g2_nand2b_1 _13880_ (.Y(_05817_),
    .B(net1875),
    .A_N(_05816_));
 sg13g2_o21ai_1 _13881_ (.B1(_05817_),
    .Y(_05818_),
    .A1(net1875),
    .A2(_05813_));
 sg13g2_o21ai_1 _13882_ (.B1(net2494),
    .Y(_05819_),
    .A1(net5050),
    .A2(_05779_));
 sg13g2_a21oi_1 _13883_ (.A1(_05779_),
    .A2(_05818_),
    .Y(_00726_),
    .B1(_05819_));
 sg13g2_a22oi_1 _13884_ (.Y(_05820_),
    .B1(_05599_),
    .B2(_04633_),
    .A2(_05530_),
    .A1(net2163));
 sg13g2_nand2b_1 _13885_ (.Y(_05821_),
    .B(net1824),
    .A_N(_05820_));
 sg13g2_o21ai_1 _13886_ (.B1(_05779_),
    .Y(_05822_),
    .A1(_02815_),
    .A2(_02822_));
 sg13g2_nand3_1 _13887_ (.B(net4315),
    .C(_05822_),
    .A(net2494),
    .Y(_05823_));
 sg13g2_nand2_1 _13888_ (.Y(_00727_),
    .A(_05821_),
    .B(net4316));
 sg13g2_nor2_1 _13889_ (.A(net4397),
    .B(net1830),
    .Y(_05824_));
 sg13g2_a21oi_1 _13890_ (.A1(net1829),
    .A2(_05814_),
    .Y(_00728_),
    .B1(_05824_));
 sg13g2_nand2_1 _13891_ (.Y(_05825_),
    .A(_04578_),
    .B(net1875));
 sg13g2_nand2_1 _13892_ (.Y(_05826_),
    .A(net4937),
    .B(_05451_));
 sg13g2_a21oi_1 _13893_ (.A1(_05825_),
    .A2(_05826_),
    .Y(_00729_),
    .B1(net2444));
 sg13g2_nand2_1 _13894_ (.Y(_05827_),
    .A(_05451_),
    .B(_05825_));
 sg13g2_nand2b_1 _13895_ (.Y(_05828_),
    .B(_04602_),
    .A_N(_04646_));
 sg13g2_o21ai_1 _13896_ (.B1(net2500),
    .Y(_05829_),
    .A1(net2512),
    .A2(_05827_));
 sg13g2_a21oi_1 _13897_ (.A1(_05827_),
    .A2(_05828_),
    .Y(_00730_),
    .B1(_05829_));
 sg13g2_nor2b_1 _13898_ (.A(_04651_),
    .B_N(_04765_),
    .Y(_00731_));
 sg13g2_nor3_1 _13899_ (.A(net5068),
    .B(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .C(net2321),
    .Y(_05830_));
 sg13g2_o21ai_1 _13900_ (.B1(net5234),
    .Y(_05831_),
    .A1(net5068),
    .A2(net2321));
 sg13g2_nand2_1 _13901_ (.Y(_05832_),
    .A(net2498),
    .B(_05831_));
 sg13g2_nor2_1 _13902_ (.A(net5069),
    .B(_05832_),
    .Y(_00732_));
 sg13g2_and2_1 _13903_ (.A(_02034_),
    .B(_05831_),
    .X(_05833_));
 sg13g2_nor2_1 _13904_ (.A(_02034_),
    .B(_05831_),
    .Y(_05834_));
 sg13g2_nor3_1 _13905_ (.A(net2450),
    .B(_05833_),
    .C(net4868),
    .Y(_00733_));
 sg13g2_nor2_1 _13906_ (.A(net4841),
    .B(_05834_),
    .Y(_05835_));
 sg13g2_and2_1 _13907_ (.A(net4841),
    .B(_05834_),
    .X(_05836_));
 sg13g2_nor3_1 _13908_ (.A(net2450),
    .B(net4842),
    .C(_05836_),
    .Y(_00734_));
 sg13g2_o21ai_1 _13909_ (.B1(net2498),
    .Y(_05837_),
    .A1(net4398),
    .A2(_05836_));
 sg13g2_a21oi_1 _13910_ (.A1(net4398),
    .A2(_05836_),
    .Y(_00735_),
    .B1(_05837_));
 sg13g2_mux2_1 _13911_ (.A0(\i_tinyqv.cpu.i_core.i_instrret.add ),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.cy ),
    .S(net2319),
    .X(_05838_));
 sg13g2_and2_1 _13912_ (.A(net5090),
    .B(_05838_),
    .X(_05839_));
 sg13g2_and2_1 _13913_ (.A(net5065),
    .B(_05839_),
    .X(_05840_));
 sg13g2_nand2_1 _13914_ (.Y(_05841_),
    .A(net5135),
    .B(_05840_));
 sg13g2_nor3_1 _13915_ (.A(net2450),
    .B(_02081_),
    .C(_05841_),
    .Y(_00736_));
 sg13g2_nand2_1 _13916_ (.Y(_05842_),
    .A(net2322),
    .B(_02817_));
 sg13g2_mux2_1 _13917_ (.A0(_02719_),
    .A1(_02730_),
    .S(_02791_),
    .X(_05843_));
 sg13g2_mux2_1 _13918_ (.A0(_05843_),
    .A1(net4672),
    .S(_05842_),
    .X(_00737_));
 sg13g2_and3_1 _13919_ (.X(_00738_),
    .A(net2498),
    .B(net4398),
    .C(_05836_));
 sg13g2_o21ai_1 _13920_ (.B1(net2498),
    .Y(_05844_),
    .A1(net5090),
    .A2(_05838_));
 sg13g2_nor2_1 _13921_ (.A(_05839_),
    .B(net5091),
    .Y(_00739_));
 sg13g2_o21ai_1 _13922_ (.B1(net2498),
    .Y(_05845_),
    .A1(net5065),
    .A2(_05839_));
 sg13g2_nor2_1 _13923_ (.A(_05840_),
    .B(net5066),
    .Y(_00740_));
 sg13g2_o21ai_1 _13924_ (.B1(net2498),
    .Y(_05846_),
    .A1(net5135),
    .A2(_05840_));
 sg13g2_nor2b_1 _13925_ (.A(_05846_),
    .B_N(_05841_),
    .Y(_00741_));
 sg13g2_xnor2_1 _13926_ (.Y(_05847_),
    .A(_02081_),
    .B(_05841_));
 sg13g2_nor2_1 _13927_ (.A(net2450),
    .B(_05847_),
    .Y(_00742_));
 sg13g2_nand2_1 _13928_ (.Y(_05848_),
    .A(net4278),
    .B(net2341));
 sg13g2_nor2_2 _13929_ (.A(_02473_),
    .B(net2341),
    .Y(_05849_));
 sg13g2_nand3_1 _13930_ (.B(net2081),
    .C(_05849_),
    .A(net2549),
    .Y(_05850_));
 sg13g2_and3_2 _13931_ (.X(_05851_),
    .A(net2638),
    .B(_05848_),
    .C(_05850_));
 sg13g2_nand3_1 _13932_ (.B(_05848_),
    .C(_05850_),
    .A(net2638),
    .Y(_05852_));
 sg13g2_nand2_1 _13933_ (.Y(_05853_),
    .A(net4943),
    .B(net2308));
 sg13g2_nand2_1 _13934_ (.Y(_05854_),
    .A(\crc16_read[9] ),
    .B(net2306));
 sg13g2_nand3_1 _13935_ (.B(_05853_),
    .C(_05854_),
    .A(_05851_),
    .Y(_00743_));
 sg13g2_nand2_1 _13936_ (.Y(_05855_),
    .A(net5099),
    .B(net2308));
 sg13g2_nand2_1 _13937_ (.Y(_05856_),
    .A(net4981),
    .B(net2306));
 sg13g2_nand3_1 _13938_ (.B(_05855_),
    .C(_05856_),
    .A(_05851_),
    .Y(_00744_));
 sg13g2_nand2_1 _13939_ (.Y(_05857_),
    .A(net4981),
    .B(net2309));
 sg13g2_nand2_1 _13940_ (.Y(_05858_),
    .A(net4938),
    .B(net2307));
 sg13g2_nand3_1 _13941_ (.B(_05857_),
    .C(_05858_),
    .A(_05851_),
    .Y(_00745_));
 sg13g2_nand2_1 _13942_ (.Y(_05859_),
    .A(net4938),
    .B(net2308));
 sg13g2_nand2_1 _13943_ (.Y(_05860_),
    .A(\crc16_read[12] ),
    .B(net2306));
 sg13g2_nand3_1 _13944_ (.B(_05859_),
    .C(_05860_),
    .A(_05851_),
    .Y(_00746_));
 sg13g2_nand2_1 _13945_ (.Y(_05861_),
    .A(\crc16_read[12] ),
    .B(net2309));
 sg13g2_nand2_1 _13946_ (.Y(_05862_),
    .A(net4751),
    .B(_03538_));
 sg13g2_nand3_1 _13947_ (.B(_05861_),
    .C(net4752),
    .A(_05851_),
    .Y(_00747_));
 sg13g2_xor2_1 _13948_ (.B(net4785),
    .A(net4832),
    .X(_05863_));
 sg13g2_nand2_1 _13949_ (.Y(_05864_),
    .A(_01941_),
    .B(net2309));
 sg13g2_o21ai_1 _13950_ (.B1(_05864_),
    .Y(_05865_),
    .A1(net2309),
    .A2(_05863_));
 sg13g2_nand2_1 _13951_ (.Y(_00748_),
    .A(_05851_),
    .B(_05865_));
 sg13g2_nand2_1 _13952_ (.Y(_05866_),
    .A(net4785),
    .B(net2309));
 sg13g2_nand2_1 _13953_ (.Y(_05867_),
    .A(\crc16_read[15] ),
    .B(net2307));
 sg13g2_nand3_1 _13954_ (.B(_05866_),
    .C(_05867_),
    .A(_05851_),
    .Y(_00749_));
 sg13g2_nand2_1 _13955_ (.Y(_05868_),
    .A(net4850),
    .B(net2308));
 sg13g2_nand2_1 _13956_ (.Y(_05869_),
    .A(net4832),
    .B(net2307));
 sg13g2_nand3_1 _13957_ (.B(_05868_),
    .C(_05869_),
    .A(_05851_),
    .Y(_00750_));
 sg13g2_nor2_2 _13958_ (.A(net2318),
    .B(_02818_),
    .Y(_05870_));
 sg13g2_nor2_1 _13959_ (.A(net3866),
    .B(net2320),
    .Y(_05871_));
 sg13g2_nor3_1 _13960_ (.A(_03135_),
    .B(_05870_),
    .C(_05871_),
    .Y(_00751_));
 sg13g2_and2_1 _13961_ (.A(net2500),
    .B(_03151_),
    .X(_05872_));
 sg13g2_nand4_1 _13962_ (.B(_02802_),
    .C(_02812_),
    .A(net2317),
    .Y(_05873_),
    .D(_05872_));
 sg13g2_o21ai_1 _13963_ (.B1(_05873_),
    .Y(_00752_),
    .A1(_01962_),
    .A2(_05276_));
 sg13g2_a21oi_1 _13964_ (.A1(\i_tinyqv.cpu.i_core.cycle[0] ),
    .A2(net2317),
    .Y(_05874_),
    .B1(net4136));
 sg13g2_nor3_1 _13965_ (.A(net2444),
    .B(_02813_),
    .C(net4137),
    .Y(_00753_));
 sg13g2_nor2_1 _13966_ (.A(_05386_),
    .B(_05390_),
    .Y(_05875_));
 sg13g2_and4_1 _13967_ (.A(_05369_),
    .B(_05378_),
    .C(_05395_),
    .D(_05430_),
    .X(_05876_));
 sg13g2_nand3_1 _13968_ (.B(_05358_),
    .C(_05394_),
    .A(_05356_),
    .Y(_05877_));
 sg13g2_a22oi_1 _13969_ (.Y(_05878_),
    .B1(_05387_),
    .B2(net2543),
    .A2(_05360_),
    .A1(_05359_));
 sg13g2_nand2_1 _13970_ (.Y(_05879_),
    .A(_05877_),
    .B(_05878_));
 sg13g2_a21oi_1 _13971_ (.A1(_05875_),
    .A2(_05876_),
    .Y(_05880_),
    .B1(_05879_));
 sg13g2_a21oi_1 _13972_ (.A1(_05357_),
    .A2(_05394_),
    .Y(_05881_),
    .B1(_05374_));
 sg13g2_nand4_1 _13973_ (.B(_05437_),
    .C(_05880_),
    .A(_05428_),
    .Y(_05882_),
    .D(_05881_));
 sg13g2_or2_1 _13974_ (.X(_05883_),
    .B(_05882_),
    .A(_05875_));
 sg13g2_inv_1 _13975_ (.Y(_05884_),
    .A(_05883_));
 sg13g2_nand2_1 _13976_ (.Y(_05885_),
    .A(net2507),
    .B(_05882_));
 sg13g2_o21ai_1 _13977_ (.B1(_05885_),
    .Y(_00754_),
    .A1(net2508),
    .A2(_05883_));
 sg13g2_nand2_1 _13978_ (.Y(_05886_),
    .A(net2506),
    .B(_05882_));
 sg13g2_xor2_1 _13979_ (.B(net2506),
    .A(net2507),
    .X(_05887_));
 sg13g2_o21ai_1 _13980_ (.B1(_05886_),
    .Y(_00755_),
    .A1(_05883_),
    .A2(_05887_));
 sg13g2_nand2_1 _13981_ (.Y(_05888_),
    .A(net4881),
    .B(_05882_));
 sg13g2_xnor2_1 _13982_ (.Y(_05889_),
    .A(net4881),
    .B(_05380_));
 sg13g2_o21ai_1 _13983_ (.B1(_05888_),
    .Y(_00756_),
    .A1(_05883_),
    .A2(_05889_));
 sg13g2_xnor2_1 _13984_ (.Y(_05890_),
    .A(net4865),
    .B(_05381_));
 sg13g2_a22oi_1 _13985_ (.Y(_00757_),
    .B1(_05884_),
    .B2(_05890_),
    .A2(_05882_),
    .A1(_02023_));
 sg13g2_nand2_1 _13986_ (.Y(_05891_),
    .A(net3614),
    .B(net2319));
 sg13g2_o21ai_1 _13987_ (.B1(_05891_),
    .Y(_00758_),
    .A1(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .A2(_04545_));
 sg13g2_and3_1 _13988_ (.X(_05892_),
    .A(net4398),
    .B(net2317),
    .C(_05836_));
 sg13g2_and2_1 _13989_ (.A(net4810),
    .B(_05892_),
    .X(_05893_));
 sg13g2_o21ai_1 _13990_ (.B1(net2498),
    .Y(_05894_),
    .A1(net4810),
    .A2(_05892_));
 sg13g2_nor2_1 _13991_ (.A(_05893_),
    .B(_05894_),
    .Y(_00759_));
 sg13g2_nand2_1 _13992_ (.Y(_05895_),
    .A(net4946),
    .B(_05893_));
 sg13g2_o21ai_1 _13993_ (.B1(net2499),
    .Y(_05896_),
    .A1(net4946),
    .A2(_05893_));
 sg13g2_nor2b_1 _13994_ (.A(_05896_),
    .B_N(_05895_),
    .Y(_00760_));
 sg13g2_o21ai_1 _13995_ (.B1(net2499),
    .Y(_05897_),
    .A1(_01961_),
    .A2(_05895_));
 sg13g2_a21oi_1 _13996_ (.A1(_01961_),
    .A2(_05895_),
    .Y(_00761_),
    .B1(_05897_));
 sg13g2_o21ai_1 _13997_ (.B1(net2499),
    .Y(_05898_),
    .A1(net4945),
    .A2(_04545_));
 sg13g2_nor2_1 _13998_ (.A(net3614),
    .B(_05898_),
    .Y(_05899_));
 sg13g2_or2_1 _13999_ (.X(_05900_),
    .B(_05898_),
    .A(net3614));
 sg13g2_nand2_1 _14000_ (.Y(_05901_),
    .A(_02550_),
    .B(_05899_));
 sg13g2_mux2_1 _14001_ (.A0(\dio1_sync[1] ),
    .A1(net4151),
    .S(_05901_),
    .X(_00762_));
 sg13g2_mux2_1 _14002_ (.A0(timer_irq),
    .A1(net4205),
    .S(_05901_),
    .X(_00763_));
 sg13g2_nand2_1 _14003_ (.Y(_05902_),
    .A(net4061),
    .B(_03387_));
 sg13g2_nand2_2 _14004_ (.Y(_05903_),
    .A(net2500),
    .B(net2355));
 sg13g2_nor2_2 _14005_ (.A(_02794_),
    .B(_02810_),
    .Y(_05904_));
 sg13g2_or4_1 _14006_ (.A(_02794_),
    .B(_02810_),
    .C(_03377_),
    .D(_03385_),
    .X(_05905_));
 sg13g2_o21ai_1 _14007_ (.B1(_04548_),
    .Y(_05906_),
    .A1(_02703_),
    .A2(_05905_));
 sg13g2_a21oi_1 _14008_ (.A1(_02061_),
    .A2(_05905_),
    .Y(_05907_),
    .B1(_05906_));
 sg13g2_a21oi_1 _14009_ (.A1(_02711_),
    .A2(_04549_),
    .Y(_05908_),
    .B1(_05907_));
 sg13g2_o21ai_1 _14010_ (.B1(_05902_),
    .Y(_00764_),
    .A1(_05903_),
    .A2(_05908_));
 sg13g2_mux2_1 _14011_ (.A0(_02667_),
    .A1(\i_tinyqv.cpu.i_core.mepc[1] ),
    .S(_05905_),
    .X(_05909_));
 sg13g2_a21oi_1 _14012_ (.A1(_02671_),
    .A2(_04549_),
    .Y(_05910_),
    .B1(_05903_));
 sg13g2_o21ai_1 _14013_ (.B1(_05910_),
    .Y(_05911_),
    .A1(_04549_),
    .A2(_05909_));
 sg13g2_o21ai_1 _14014_ (.B1(_05911_),
    .Y(_00765_),
    .A1(_02043_),
    .A2(net2352));
 sg13g2_nand2b_1 _14015_ (.Y(_05912_),
    .B(_02626_),
    .A_N(_05905_));
 sg13g2_a21oi_1 _14016_ (.A1(net4275),
    .A2(_05905_),
    .Y(_05913_),
    .B1(_04549_));
 sg13g2_a21oi_1 _14017_ (.A1(_05912_),
    .A2(_05913_),
    .Y(_05914_),
    .B1(_05903_));
 sg13g2_o21ai_1 _14018_ (.B1(_05914_),
    .Y(_05915_),
    .A1(_02631_),
    .A2(_04548_));
 sg13g2_o21ai_1 _14019_ (.B1(_05915_),
    .Y(_00766_),
    .A1(_02044_),
    .A2(net2354));
 sg13g2_nand2b_1 _14020_ (.Y(_05916_),
    .B(_02537_),
    .A_N(_05905_));
 sg13g2_a21oi_1 _14021_ (.A1(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A2(_05905_),
    .Y(_05917_),
    .B1(_04549_));
 sg13g2_a21oi_1 _14022_ (.A1(_05916_),
    .A2(_05917_),
    .Y(_05918_),
    .B1(_05903_));
 sg13g2_o21ai_1 _14023_ (.B1(_05918_),
    .Y(_05919_),
    .A1(_02553_),
    .A2(_04548_));
 sg13g2_o21ai_1 _14024_ (.B1(_05919_),
    .Y(_00767_),
    .A1(_02045_),
    .A2(net2352));
 sg13g2_o21ai_1 _14025_ (.B1(_04550_),
    .Y(_05920_),
    .A1(net4945),
    .A2(net2298));
 sg13g2_nand2_1 _14026_ (.Y(_00768_),
    .A(_05899_),
    .B(_05920_));
 sg13g2_nor3_1 _14027_ (.A(_03771_),
    .B(_04551_),
    .C(net2298),
    .Y(_05921_));
 sg13g2_nand3_1 _14028_ (.B(_02537_),
    .C(_02809_),
    .A(net2528),
    .Y(_05922_));
 sg13g2_nor4_1 _14029_ (.A(_03770_),
    .B(_04551_),
    .C(net2298),
    .D(_05904_),
    .Y(_05923_));
 sg13g2_and2_1 _14030_ (.A(_05922_),
    .B(_05923_),
    .X(_05924_));
 sg13g2_or2_1 _14031_ (.X(_05925_),
    .B(_05924_),
    .A(_05921_));
 sg13g2_a21oi_2 _14032_ (.B1(_03139_),
    .Y(_05926_),
    .A2(net2530),
    .A1(net2528));
 sg13g2_and3_1 _14033_ (.X(_05927_),
    .A(_02537_),
    .B(_04550_),
    .C(_05926_));
 sg13g2_nor2_1 _14034_ (.A(_04551_),
    .B(net2295),
    .Y(_05928_));
 sg13g2_a21oi_1 _14035_ (.A1(net3964),
    .A2(_05928_),
    .Y(_05929_),
    .B1(_05927_));
 sg13g2_a21oi_1 _14036_ (.A1(net4825),
    .A2(_05925_),
    .Y(_05930_),
    .B1(_05900_));
 sg13g2_o21ai_1 _14037_ (.B1(_05930_),
    .Y(_00769_),
    .A1(_05925_),
    .A2(_05929_));
 sg13g2_a21oi_1 _14038_ (.A1(_03894_),
    .A2(net2295),
    .Y(_05931_),
    .B1(_04551_));
 sg13g2_nor3_1 _14039_ (.A(_02707_),
    .B(_03770_),
    .C(net2298),
    .Y(_05932_));
 sg13g2_or3_1 _14040_ (.A(_05924_),
    .B(_05931_),
    .C(_05932_),
    .X(_05933_));
 sg13g2_a21oi_1 _14041_ (.A1(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .A2(_04551_),
    .Y(_05934_),
    .B1(_05927_));
 sg13g2_nor2b_1 _14042_ (.A(_05933_),
    .B_N(_05934_),
    .Y(_05935_));
 sg13g2_nor2b_1 _14043_ (.A(net3964),
    .B_N(_05933_),
    .Y(_05936_));
 sg13g2_nor3_1 _14044_ (.A(_05900_),
    .B(_05935_),
    .C(_05936_),
    .Y(_00770_));
 sg13g2_nor2b_1 _14045_ (.A(_05506_),
    .B_N(_05478_),
    .Y(_05937_));
 sg13g2_nand3_1 _14046_ (.B(_05572_),
    .C(_05937_),
    .A(_05471_),
    .Y(_05938_));
 sg13g2_or2_1 _14047_ (.X(_05939_),
    .B(_05938_),
    .A(_05504_));
 sg13g2_nand2b_2 _14048_ (.Y(_05940_),
    .B(_05481_),
    .A_N(_05939_));
 sg13g2_nor3_1 _14049_ (.A(_04616_),
    .B(_05457_),
    .C(_05475_),
    .Y(_05941_));
 sg13g2_nor3_1 _14050_ (.A(_04714_),
    .B(_05480_),
    .C(_05938_),
    .Y(_05942_));
 sg13g2_nand2_2 _14051_ (.Y(_05943_),
    .A(_05941_),
    .B(_05942_));
 sg13g2_a22oi_1 _14052_ (.Y(_05944_),
    .B1(_05760_),
    .B2(_04630_),
    .A2(_04714_),
    .A1(_04612_));
 sg13g2_nand2_1 _14053_ (.Y(_05945_),
    .A(_05600_),
    .B(_05944_));
 sg13g2_mux2_1 _14054_ (.A0(_04621_),
    .A1(_05945_),
    .S(_05943_),
    .X(_05946_));
 sg13g2_a22oi_1 _14055_ (.Y(_05947_),
    .B1(_05946_),
    .B2(net2105),
    .A2(_05940_),
    .A1(_04644_));
 sg13g2_mux2_1 _14056_ (.A0(net4426),
    .A1(_05947_),
    .S(net1874),
    .X(_05948_));
 sg13g2_nand2_1 _14057_ (.Y(_05949_),
    .A(net4426),
    .B(net1809));
 sg13g2_o21ai_1 _14058_ (.B1(_05949_),
    .Y(_00771_),
    .A1(net1809),
    .A2(_05948_));
 sg13g2_nand2_1 _14059_ (.Y(_05950_),
    .A(_04635_),
    .B(_05940_));
 sg13g2_o21ai_1 _14060_ (.B1(_05950_),
    .Y(_05951_),
    .A1(_05562_),
    .A2(_05943_));
 sg13g2_nor3_1 _14061_ (.A(_03148_),
    .B(_04017_),
    .C(net1873),
    .Y(_05952_));
 sg13g2_a21oi_1 _14062_ (.A1(net1873),
    .A2(_05951_),
    .Y(_05953_),
    .B1(_05952_));
 sg13g2_nand2_1 _14063_ (.Y(_05954_),
    .A(net4105),
    .B(net1808));
 sg13g2_o21ai_1 _14064_ (.B1(_05954_),
    .Y(_00772_),
    .A1(net1808),
    .A2(_05953_));
 sg13g2_nor2_1 _14065_ (.A(_05573_),
    .B(_05943_),
    .Y(_05955_));
 sg13g2_a21oi_2 _14066_ (.B1(_05955_),
    .Y(_05956_),
    .A2(_05940_),
    .A1(_04633_));
 sg13g2_xor2_1 _14067_ (.B(_03148_),
    .A(net2505),
    .X(_05957_));
 sg13g2_nand2_1 _14068_ (.Y(_05958_),
    .A(net1874),
    .B(_05956_));
 sg13g2_o21ai_1 _14069_ (.B1(_05958_),
    .Y(_05959_),
    .A1(net1873),
    .A2(_05957_));
 sg13g2_nand2_1 _14070_ (.Y(_05960_),
    .A(net2505),
    .B(net1808));
 sg13g2_o21ai_1 _14071_ (.B1(_05960_),
    .Y(_00773_),
    .A1(net1808),
    .A2(_05959_));
 sg13g2_o21ai_1 _14072_ (.B1(net2160),
    .Y(_05961_),
    .A1(_05599_),
    .A2(_05939_));
 sg13g2_o21ai_1 _14073_ (.B1(_05961_),
    .Y(_05962_),
    .A1(net2109),
    .A2(_05943_));
 sg13g2_o21ai_1 _14074_ (.B1(net1875),
    .Y(_05963_),
    .A1(_05480_),
    .A2(_05962_));
 sg13g2_xor2_1 _14075_ (.B(_03149_),
    .A(net2504),
    .X(_05964_));
 sg13g2_o21ai_1 _14076_ (.B1(_05963_),
    .Y(_05965_),
    .A1(net1873),
    .A2(_05964_));
 sg13g2_mux2_1 _14077_ (.A0(_05965_),
    .A1(net2504),
    .S(net1808),
    .X(_00774_));
 sg13g2_nor2_1 _14078_ (.A(net4402),
    .B(net1855),
    .Y(_05966_));
 sg13g2_and3_1 _14079_ (.X(_05967_),
    .A(net2573),
    .B(net2574),
    .C(\i_tinyqv.cpu.instr_write_offset[3] ));
 sg13g2_a21oi_1 _14080_ (.A1(net2574),
    .A2(\i_tinyqv.cpu.instr_write_offset[3] ),
    .Y(_05968_),
    .B1(net2573));
 sg13g2_or3_1 _14081_ (.A(net2563),
    .B(_05967_),
    .C(_05968_),
    .X(_05969_));
 sg13g2_o21ai_1 _14082_ (.B1(_05969_),
    .Y(_05970_),
    .A1(_01967_),
    .A2(_05031_));
 sg13g2_o21ai_1 _14083_ (.B1(net1833),
    .Y(_05971_),
    .A1(net1860),
    .A2(_05970_));
 sg13g2_nor3_2 _14084_ (.A(net2607),
    .B(_01982_),
    .C(_04039_),
    .Y(_05972_));
 sg13g2_nand2_2 _14085_ (.Y(_05973_),
    .A(net4625),
    .B(_04040_));
 sg13g2_nor2_2 _14086_ (.A(net1831),
    .B(net2281),
    .Y(_05974_));
 sg13g2_a22oi_1 _14087_ (.Y(_05975_),
    .B1(net1806),
    .B2(net3828),
    .A2(net2282),
    .A1(net3479));
 sg13g2_o21ai_1 _14088_ (.B1(_05975_),
    .Y(_00775_),
    .A1(_05966_),
    .A2(_05971_));
 sg13g2_nor2_1 _14089_ (.A(\addr[5] ),
    .B(net1855),
    .Y(_05976_));
 sg13g2_nor2_1 _14090_ (.A(_01967_),
    .B(_05038_),
    .Y(_05977_));
 sg13g2_and2_1 _14091_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(_05967_),
    .X(_05978_));
 sg13g2_o21ai_1 _14092_ (.B1(net2441),
    .Y(_05979_),
    .A1(\i_tinyqv.cpu.instr_data_start[5] ),
    .A2(_05967_));
 sg13g2_o21ai_1 _14093_ (.B1(net1856),
    .Y(_05980_),
    .A1(_05978_),
    .A2(_05979_));
 sg13g2_o21ai_1 _14094_ (.B1(net1833),
    .Y(_05981_),
    .A1(_05977_),
    .A2(_05980_));
 sg13g2_a22oi_1 _14095_ (.Y(_05982_),
    .B1(net1806),
    .B2(net4211),
    .A2(net2282),
    .A1(net3942));
 sg13g2_o21ai_1 _14096_ (.B1(_05982_),
    .Y(_00776_),
    .A1(_05976_),
    .A2(_05981_));
 sg13g2_xnor2_1 _14097_ (.Y(_05983_),
    .A(_01977_),
    .B(_05978_));
 sg13g2_nor2_1 _14098_ (.A(net2564),
    .B(_05983_),
    .Y(_05984_));
 sg13g2_a21oi_1 _14099_ (.A1(net2563),
    .A2(_05054_),
    .Y(_05985_),
    .B1(_05984_));
 sg13g2_nand2_1 _14100_ (.Y(_05986_),
    .A(net1856),
    .B(_05985_));
 sg13g2_a21oi_1 _14101_ (.A1(\addr[6] ),
    .A2(net1860),
    .Y(_05987_),
    .B1(net1836));
 sg13g2_nand2_1 _14102_ (.Y(_05988_),
    .A(net3838),
    .B(net2282));
 sg13g2_a21oi_1 _14103_ (.A1(net3602),
    .A2(net2221),
    .Y(_05989_),
    .B1(net1833));
 sg13g2_a22oi_1 _14104_ (.Y(_00777_),
    .B1(_05988_),
    .B2(_05989_),
    .A2(_05987_),
    .A1(_05986_));
 sg13g2_a21o_1 _14105_ (.A2(_05978_),
    .A1(\i_tinyqv.cpu.instr_data_start[6] ),
    .B1(net2572),
    .X(_05990_));
 sg13g2_nand3_1 _14106_ (.B(\i_tinyqv.cpu.instr_data_start[6] ),
    .C(_05978_),
    .A(\i_tinyqv.cpu.instr_data_start[7] ),
    .Y(_05991_));
 sg13g2_a21oi_1 _14107_ (.A1(_05990_),
    .A2(_05991_),
    .Y(_05992_),
    .B1(net2564));
 sg13g2_and2_1 _14108_ (.A(net2564),
    .B(_05062_),
    .X(_05993_));
 sg13g2_o21ai_1 _14109_ (.B1(net1856),
    .Y(_05994_),
    .A1(_05992_),
    .A2(_05993_));
 sg13g2_o21ai_1 _14110_ (.B1(_05994_),
    .Y(_05995_),
    .A1(net4232),
    .A2(net1855));
 sg13g2_a22oi_1 _14111_ (.Y(_05996_),
    .B1(net1806),
    .B2(net4344),
    .A2(_05972_),
    .A1(net3566));
 sg13g2_o21ai_1 _14112_ (.B1(net4345),
    .Y(_00778_),
    .A1(net1836),
    .A2(_05995_));
 sg13g2_or2_1 _14113_ (.X(_05997_),
    .B(_05991_),
    .A(_01976_));
 sg13g2_a21oi_1 _14114_ (.A1(_01976_),
    .A2(_05991_),
    .Y(_05998_),
    .B1(net2563));
 sg13g2_a22oi_1 _14115_ (.Y(_05999_),
    .B1(_05997_),
    .B2(_05998_),
    .A2(_05074_),
    .A1(net2564));
 sg13g2_nand2_1 _14116_ (.Y(_06000_),
    .A(net3828),
    .B(net2282));
 sg13g2_nor2_1 _14117_ (.A(net1859),
    .B(_05999_),
    .Y(_06001_));
 sg13g2_a21oi_1 _14118_ (.A1(\addr[8] ),
    .A2(net1859),
    .Y(_06002_),
    .B1(_06001_));
 sg13g2_a21oi_1 _14119_ (.A1(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .A2(net2221),
    .Y(_06003_),
    .B1(net1833));
 sg13g2_a22oi_1 _14120_ (.Y(_00779_),
    .B1(_06003_),
    .B2(_06000_),
    .A2(_06002_),
    .A1(net1834));
 sg13g2_nand2_1 _14121_ (.Y(_06004_),
    .A(_01975_),
    .B(_05997_));
 sg13g2_nor2_2 _14122_ (.A(_01975_),
    .B(_05997_),
    .Y(_06005_));
 sg13g2_nor2_1 _14123_ (.A(net2563),
    .B(_06005_),
    .Y(_06006_));
 sg13g2_a221oi_1 _14124_ (.B2(_06006_),
    .C1(net1859),
    .B1(_06004_),
    .A1(net2563),
    .Y(_06007_),
    .A2(_05091_));
 sg13g2_o21ai_1 _14125_ (.B1(net1833),
    .Y(_06008_),
    .A1(net4342),
    .A2(net1855));
 sg13g2_a22oi_1 _14126_ (.Y(_06009_),
    .B1(net1806),
    .B2(net4772),
    .A2(net2282),
    .A1(net4211));
 sg13g2_o21ai_1 _14127_ (.B1(_06009_),
    .Y(_00780_),
    .A1(_06007_),
    .A2(_06008_));
 sg13g2_o21ai_1 _14128_ (.B1(_01967_),
    .Y(_06010_),
    .A1(net2570),
    .A2(_06005_));
 sg13g2_a21oi_1 _14129_ (.A1(net2570),
    .A2(_06005_),
    .Y(_06011_),
    .B1(_06010_));
 sg13g2_a21oi_1 _14130_ (.A1(net2563),
    .A2(_05102_),
    .Y(_06012_),
    .B1(_06011_));
 sg13g2_nand2_1 _14131_ (.Y(_06013_),
    .A(net3602),
    .B(_05972_));
 sg13g2_nor2_1 _14132_ (.A(net1859),
    .B(_06012_),
    .Y(_06014_));
 sg13g2_a21oi_1 _14133_ (.A1(\addr[10] ),
    .A2(net1859),
    .Y(_06015_),
    .B1(_06014_));
 sg13g2_a21oi_1 _14134_ (.A1(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .A2(net2221),
    .Y(_06016_),
    .B1(net1832));
 sg13g2_a22oi_1 _14135_ (.Y(_00781_),
    .B1(_06016_),
    .B2(net3603),
    .A2(_06015_),
    .A1(net1833));
 sg13g2_nand3_1 _14136_ (.B(net2570),
    .C(_06005_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .Y(_06017_));
 sg13g2_a21oi_1 _14137_ (.A1(net2570),
    .A2(_06005_),
    .Y(_06018_),
    .B1(\i_tinyqv.cpu.instr_data_start[11] ));
 sg13g2_nor2_1 _14138_ (.A(net2562),
    .B(_06018_),
    .Y(_06019_));
 sg13g2_a22oi_1 _14139_ (.Y(_06020_),
    .B1(_06017_),
    .B2(_06019_),
    .A2(_05112_),
    .A1(net2562));
 sg13g2_a21oi_1 _14140_ (.A1(net1853),
    .A2(_06020_),
    .Y(_06021_),
    .B1(net1836));
 sg13g2_o21ai_1 _14141_ (.B1(_06021_),
    .Y(_06022_),
    .A1(net4225),
    .A2(net1853));
 sg13g2_a22oi_1 _14142_ (.Y(_06023_),
    .B1(net1806),
    .B2(net3625),
    .A2(_05972_),
    .A1(net4344));
 sg13g2_nand2_1 _14143_ (.Y(_00782_),
    .A(_06022_),
    .B(_06023_));
 sg13g2_nor2_1 _14144_ (.A(_01974_),
    .B(_06017_),
    .Y(_06024_));
 sg13g2_xnor2_1 _14145_ (.Y(_06025_),
    .A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(_06017_));
 sg13g2_nand2_1 _14146_ (.Y(_06026_),
    .A(net2562),
    .B(_05127_));
 sg13g2_o21ai_1 _14147_ (.B1(_06026_),
    .Y(_06027_),
    .A1(net2562),
    .A2(_06025_));
 sg13g2_a21oi_1 _14148_ (.A1(\addr[12] ),
    .A2(net1857),
    .Y(_06028_),
    .B1(net1836));
 sg13g2_o21ai_1 _14149_ (.B1(_06028_),
    .Y(_06029_),
    .A1(net1858),
    .A2(_06027_));
 sg13g2_o21ai_1 _14150_ (.B1(_06029_),
    .Y(_06030_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .A2(_05973_));
 sg13g2_a21oi_1 _14151_ (.A1(_02040_),
    .A2(net1807),
    .Y(_00783_),
    .B1(_06030_));
 sg13g2_and2_1 _14152_ (.A(net2569),
    .B(_06024_),
    .X(_06031_));
 sg13g2_xor2_1 _14153_ (.B(_06024_),
    .A(net2569),
    .X(_06032_));
 sg13g2_nor2_1 _14154_ (.A(net2440),
    .B(_05141_),
    .Y(_06033_));
 sg13g2_a21oi_1 _14155_ (.A1(net2440),
    .A2(_06032_),
    .Y(_06034_),
    .B1(_06033_));
 sg13g2_a21oi_1 _14156_ (.A1(\addr[13] ),
    .A2(net1857),
    .Y(_06035_),
    .B1(net1835));
 sg13g2_o21ai_1 _14157_ (.B1(_06035_),
    .Y(_06036_),
    .A1(net1857),
    .A2(_06034_));
 sg13g2_o21ai_1 _14158_ (.B1(_06036_),
    .Y(_06037_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .A2(net2221));
 sg13g2_a21oi_1 _14159_ (.A1(_02041_),
    .A2(net1807),
    .Y(_00784_),
    .B1(_06037_));
 sg13g2_xnor2_1 _14160_ (.Y(_06038_),
    .A(net2568),
    .B(_06031_));
 sg13g2_nand2_1 _14161_ (.Y(_06039_),
    .A(net2440),
    .B(_06038_));
 sg13g2_o21ai_1 _14162_ (.B1(_06039_),
    .Y(_06040_),
    .A1(net2440),
    .A2(_05152_));
 sg13g2_nor2_1 _14163_ (.A(net1857),
    .B(_06040_),
    .Y(_06041_));
 sg13g2_a21oi_1 _14164_ (.A1(net4400),
    .A2(net1857),
    .Y(_06042_),
    .B1(_06041_));
 sg13g2_nand2b_1 _14165_ (.Y(_06043_),
    .B(net1807),
    .A_N(\i_tinyqv.mem.q_ctrl.addr[14] ));
 sg13g2_o21ai_1 _14166_ (.B1(_06043_),
    .Y(_06044_),
    .A1(net4781),
    .A2(net2221));
 sg13g2_a21oi_1 _14167_ (.A1(net1832),
    .A2(_06042_),
    .Y(_00785_),
    .B1(net4782));
 sg13g2_and3_1 _14168_ (.X(_06045_),
    .A(\i_tinyqv.cpu.instr_data_start[15] ),
    .B(net2568),
    .C(_06031_));
 sg13g2_a21oi_1 _14169_ (.A1(net2568),
    .A2(_06031_),
    .Y(_06046_),
    .B1(\i_tinyqv.cpu.instr_data_start[15] ));
 sg13g2_nor3_1 _14170_ (.A(net2561),
    .B(_06045_),
    .C(_06046_),
    .Y(_06047_));
 sg13g2_nor2_1 _14171_ (.A(net2440),
    .B(_05165_),
    .Y(_06048_));
 sg13g2_nand2_1 _14172_ (.Y(_06049_),
    .A(net3625),
    .B(net2282));
 sg13g2_o21ai_1 _14173_ (.B1(net1854),
    .Y(_06050_),
    .A1(_06047_),
    .A2(_06048_));
 sg13g2_a21oi_1 _14174_ (.A1(\addr[15] ),
    .A2(net1858),
    .Y(_06051_),
    .B1(net1835));
 sg13g2_a21oi_1 _14175_ (.A1(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .A2(net2221),
    .Y(_06052_),
    .B1(net1831));
 sg13g2_a22oi_1 _14176_ (.Y(_00786_),
    .B1(_06052_),
    .B2(_06049_),
    .A2(_06051_),
    .A1(_06050_));
 sg13g2_or2_1 _14177_ (.X(_06053_),
    .B(_06045_),
    .A(net2567));
 sg13g2_and2_1 _14178_ (.A(net2567),
    .B(_06045_),
    .X(_06054_));
 sg13g2_nor2_1 _14179_ (.A(net2561),
    .B(_06054_),
    .Y(_06055_));
 sg13g2_a221oi_1 _14180_ (.B2(_06055_),
    .C1(net1857),
    .B1(_06053_),
    .A1(net2560),
    .Y(_06056_),
    .A2(_05177_));
 sg13g2_o21ai_1 _14181_ (.B1(net1831),
    .Y(_06057_),
    .A1(\addr[16] ),
    .A2(net1852));
 sg13g2_a22oi_1 _14182_ (.Y(_06058_),
    .B1(net1807),
    .B2(net4285),
    .A2(net2282),
    .A1(net3627));
 sg13g2_o21ai_1 _14183_ (.B1(_06058_),
    .Y(_00787_),
    .A1(_06056_),
    .A2(_06057_));
 sg13g2_nand2_1 _14184_ (.Y(_06059_),
    .A(net2561),
    .B(_05190_));
 sg13g2_a21oi_1 _14185_ (.A1(net2566),
    .A2(_06054_),
    .Y(_06060_),
    .B1(net2561));
 sg13g2_o21ai_1 _14186_ (.B1(_06060_),
    .Y(_06061_),
    .A1(net2566),
    .A2(_06054_));
 sg13g2_nand3_1 _14187_ (.B(_06059_),
    .C(_06061_),
    .A(net1854),
    .Y(_06062_));
 sg13g2_o21ai_1 _14188_ (.B1(_06062_),
    .Y(_06063_),
    .A1(net4537),
    .A2(net1852));
 sg13g2_a22oi_1 _14189_ (.Y(_06064_),
    .B1(net1807),
    .B2(net3814),
    .A2(net2281),
    .A1(net3749));
 sg13g2_o21ai_1 _14190_ (.B1(_06064_),
    .Y(_00788_),
    .A1(net1835),
    .A2(_06063_));
 sg13g2_and3_2 _14191_ (.X(_06065_),
    .A(\i_tinyqv.cpu.instr_data_start[18] ),
    .B(net2566),
    .C(_06054_));
 sg13g2_a21oi_1 _14192_ (.A1(net2566),
    .A2(_06054_),
    .Y(_06066_),
    .B1(\i_tinyqv.cpu.instr_data_start[18] ));
 sg13g2_nor3_1 _14193_ (.A(net2561),
    .B(_06065_),
    .C(_06066_),
    .Y(_06067_));
 sg13g2_a21oi_1 _14194_ (.A1(net2561),
    .A2(_05204_),
    .Y(_06068_),
    .B1(_06067_));
 sg13g2_a21oi_1 _14195_ (.A1(net1852),
    .A2(_06068_),
    .Y(_06069_),
    .B1(net1835));
 sg13g2_o21ai_1 _14196_ (.B1(_06069_),
    .Y(_06070_),
    .A1(net4301),
    .A2(net1852));
 sg13g2_a22oi_1 _14197_ (.Y(_06071_),
    .B1(net1807),
    .B2(net4839),
    .A2(net2281),
    .A1(\i_tinyqv.mem.q_ctrl.addr[14] ));
 sg13g2_nand2_1 _14198_ (.Y(_00789_),
    .A(_06070_),
    .B(net4840));
 sg13g2_o21ai_1 _14199_ (.B1(net2440),
    .Y(_06072_),
    .A1(net2565),
    .A2(_06065_));
 sg13g2_a21o_1 _14200_ (.A2(_06065_),
    .A1(net2565),
    .B1(_06072_),
    .X(_06073_));
 sg13g2_o21ai_1 _14201_ (.B1(_06073_),
    .Y(_06074_),
    .A1(net2440),
    .A2(_05215_));
 sg13g2_nand2_1 _14202_ (.Y(_06075_),
    .A(net3887),
    .B(net2281));
 sg13g2_nand2_1 _14203_ (.Y(_06076_),
    .A(net1852),
    .B(_06074_));
 sg13g2_a21oi_1 _14204_ (.A1(\addr[19] ),
    .A2(net1857),
    .Y(_06077_),
    .B1(net1835));
 sg13g2_a21oi_1 _14205_ (.A1(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .A2(net2221),
    .Y(_06078_),
    .B1(net1831));
 sg13g2_a22oi_1 _14206_ (.Y(_00790_),
    .B1(_06078_),
    .B2(_06075_),
    .A2(_06077_),
    .A1(_06076_));
 sg13g2_a21o_1 _14207_ (.A2(_06065_),
    .A1(net2565),
    .B1(\i_tinyqv.cpu.instr_data_start[20] ),
    .X(_06079_));
 sg13g2_nand3_1 _14208_ (.B(net2565),
    .C(_06065_),
    .A(\i_tinyqv.cpu.instr_data_start[20] ),
    .Y(_06080_));
 sg13g2_nand3_1 _14209_ (.B(_06079_),
    .C(_06080_),
    .A(net2440),
    .Y(_06081_));
 sg13g2_nand2_1 _14210_ (.Y(_06082_),
    .A(net1854),
    .B(_06081_));
 sg13g2_a21oi_1 _14211_ (.A1(net2560),
    .A2(_05227_),
    .Y(_06083_),
    .B1(_06082_));
 sg13g2_mux2_1 _14212_ (.A0(net5230),
    .A1(net4285),
    .S(net2281),
    .X(_06084_));
 sg13g2_o21ai_1 _14213_ (.B1(net1831),
    .Y(_06085_),
    .A1(net4779),
    .A2(net1852));
 sg13g2_nand2_1 _14214_ (.Y(_06086_),
    .A(net1835),
    .B(_06084_));
 sg13g2_o21ai_1 _14215_ (.B1(_06086_),
    .Y(_00791_),
    .A1(_06083_),
    .A2(_06085_));
 sg13g2_nor2_1 _14216_ (.A(_01969_),
    .B(_06080_),
    .Y(_06087_));
 sg13g2_nand2_1 _14217_ (.Y(_06088_),
    .A(net3814),
    .B(net2281));
 sg13g2_a21oi_1 _14218_ (.A1(\addr[21] ),
    .A2(net1858),
    .Y(_06089_),
    .B1(net1835));
 sg13g2_xnor2_1 _14219_ (.Y(_06090_),
    .A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(_06080_));
 sg13g2_o21ai_1 _14220_ (.B1(net1854),
    .Y(_06091_),
    .A1(net2560),
    .A2(_06090_));
 sg13g2_a21o_1 _14221_ (.A2(_05240_),
    .A1(net2560),
    .B1(_06091_),
    .X(_06092_));
 sg13g2_a21oi_1 _14222_ (.A1(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .A2(net2221),
    .Y(_06093_),
    .B1(net1831));
 sg13g2_a22oi_1 _14223_ (.Y(_00792_),
    .B1(_06093_),
    .B2(_06088_),
    .A2(_06092_),
    .A1(_06089_));
 sg13g2_nand2_1 _14224_ (.Y(_06094_),
    .A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(_06087_));
 sg13g2_nor2_1 _14225_ (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(_06087_),
    .Y(_06095_));
 sg13g2_nor2_1 _14226_ (.A(net2560),
    .B(_06095_),
    .Y(_06096_));
 sg13g2_a221oi_1 _14227_ (.B2(_06096_),
    .C1(net1857),
    .B1(_06094_),
    .A1(net2560),
    .Y(_06097_),
    .A2(_05252_));
 sg13g2_o21ai_1 _14228_ (.B1(net1831),
    .Y(_06098_),
    .A1(net4299),
    .A2(net1852));
 sg13g2_a22oi_1 _14229_ (.Y(_06099_),
    .B1(net1807),
    .B2(net4632),
    .A2(net2281),
    .A1(\i_tinyqv.mem.q_ctrl.addr[18] ));
 sg13g2_o21ai_1 _14230_ (.B1(net4633),
    .Y(_00793_),
    .A1(_06097_),
    .A2(_06098_));
 sg13g2_xor2_1 _14231_ (.B(_06094_),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .X(_06100_));
 sg13g2_o21ai_1 _14232_ (.B1(net1854),
    .Y(_06101_),
    .A1(net2560),
    .A2(_06100_));
 sg13g2_a21oi_1 _14233_ (.A1(net2560),
    .A2(_05264_),
    .Y(_06102_),
    .B1(_06101_));
 sg13g2_o21ai_1 _14234_ (.B1(net1832),
    .Y(_06103_),
    .A1(\addr[23] ),
    .A2(net1853));
 sg13g2_a22oi_1 _14235_ (.Y(_06104_),
    .B1(net1807),
    .B2(net4388),
    .A2(net2281),
    .A1(\i_tinyqv.mem.q_ctrl.addr[19] ));
 sg13g2_o21ai_1 _14236_ (.B1(net4389),
    .Y(_00794_),
    .A1(_06102_),
    .A2(_06103_));
 sg13g2_nor2_1 _14237_ (.A(net2441),
    .B(_04985_),
    .Y(_06105_));
 sg13g2_a21oi_1 _14238_ (.A1(net2441),
    .A2(\i_tinyqv.cpu.instr_write_offset[1] ),
    .Y(_06106_),
    .B1(_06105_));
 sg13g2_o21ai_1 _14239_ (.B1(net1833),
    .Y(_06107_),
    .A1(\addr[1] ),
    .A2(net1855));
 sg13g2_a21oi_1 _14240_ (.A1(net1855),
    .A2(_06106_),
    .Y(_06108_),
    .B1(_06107_));
 sg13g2_a21o_1 _14241_ (.A2(net1806),
    .A1(net3942),
    .B1(_06108_),
    .X(_00795_));
 sg13g2_mux2_1 _14242_ (.A0(\i_tinyqv.cpu.instr_write_offset[2] ),
    .A1(_05003_),
    .S(net2562),
    .X(_06109_));
 sg13g2_nor2_1 _14243_ (.A(net1860),
    .B(_06109_),
    .Y(_06110_));
 sg13g2_a221oi_1 _14244_ (.B2(_04738_),
    .C1(_06110_),
    .B1(_04737_),
    .A1(_02013_),
    .Y(_06111_),
    .A2(net1859));
 sg13g2_a21o_1 _14245_ (.A2(net1806),
    .A1(net3838),
    .B1(net4035),
    .X(_00796_));
 sg13g2_nand2_1 _14246_ (.Y(_06112_),
    .A(net3566),
    .B(net1806));
 sg13g2_or2_1 _14247_ (.X(_06113_),
    .B(\i_tinyqv.cpu.instr_write_offset[3] ),
    .A(net2574));
 sg13g2_a21oi_1 _14248_ (.A1(net2574),
    .A2(\i_tinyqv.cpu.instr_write_offset[3] ),
    .Y(_06114_),
    .B1(net2563));
 sg13g2_a221oi_1 _14249_ (.B2(_06114_),
    .C1(net1859),
    .B1(_06113_),
    .A1(net2563),
    .Y(_06115_),
    .A2(_05016_));
 sg13g2_o21ai_1 _14250_ (.B1(net1833),
    .Y(_06116_),
    .A1(net2466),
    .A2(net1855));
 sg13g2_o21ai_1 _14251_ (.B1(_06112_),
    .Y(_00797_),
    .A1(_06115_),
    .A2(_06116_));
 sg13g2_nand3_1 _14252_ (.B(_02002_),
    .C(_04652_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .Y(_06117_));
 sg13g2_nor2_1 _14253_ (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .B(net1805),
    .Y(_06118_));
 sg13g2_and2_1 _14254_ (.A(net2496),
    .B(net1805),
    .X(_06119_));
 sg13g2_a21oi_1 _14255_ (.A1(_02006_),
    .A2(_06119_),
    .Y(_00798_),
    .B1(_06118_));
 sg13g2_nor2_1 _14256_ (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .B(net1805),
    .Y(_06120_));
 sg13g2_a21oi_1 _14257_ (.A1(_02011_),
    .A2(_06119_),
    .Y(_00799_),
    .B1(_06120_));
 sg13g2_nor3_1 _14258_ (.A(net3481),
    .B(net2308),
    .C(net1956),
    .Y(_00800_));
 sg13g2_nor2b_1 _14259_ (.A(net3481),
    .B_N(net4280),
    .Y(_06121_));
 sg13g2_a21oi_1 _14260_ (.A1(_01958_),
    .A2(net2305),
    .Y(_06122_),
    .B1(net4280));
 sg13g2_nor3_1 _14261_ (.A(net1956),
    .B(_06121_),
    .C(_06122_),
    .Y(_00801_));
 sg13g2_nand2_1 _14262_ (.Y(_06123_),
    .A(net4170),
    .B(_03536_));
 sg13g2_o21ai_1 _14263_ (.B1(\i_crc16.bit_cnt[2] ),
    .Y(_06124_),
    .A1(\i_crc16.bit_cnt[1] ),
    .A2(net3481));
 sg13g2_a21oi_1 _14264_ (.A1(net4171),
    .A2(_06124_),
    .Y(_00802_),
    .B1(net1956));
 sg13g2_o21ai_1 _14265_ (.B1(net2643),
    .Y(_06125_),
    .A1(net4379),
    .A2(_04320_));
 sg13g2_inv_1 _14266_ (.Y(_00803_),
    .A(_06125_));
 sg13g2_nor2_1 _14267_ (.A(_04304_),
    .B(net2065),
    .Y(_06126_));
 sg13g2_nand2_2 _14268_ (.Y(_06127_),
    .A(net2645),
    .B(_04321_));
 sg13g2_a221oi_1 _14269_ (.B2(_06127_),
    .C1(net1872),
    .B1(_04425_),
    .A1(net5291),
    .Y(_06128_),
    .A2(_04321_));
 sg13g2_a21o_1 _14270_ (.A2(net1872),
    .A1(_04327_),
    .B1(_06128_),
    .X(_00804_));
 sg13g2_xnor2_1 _14271_ (.Y(_06129_),
    .A(net5143),
    .B(\i_wdt.counter[0] ));
 sg13g2_nand2_1 _14272_ (.Y(_06130_),
    .A(_04322_),
    .B(_06129_));
 sg13g2_a22oi_1 _14273_ (.Y(_06131_),
    .B1(net1872),
    .B2(net5143),
    .A2(net2064),
    .A1(net2557));
 sg13g2_a21oi_1 _14274_ (.A1(_06130_),
    .A2(_06131_),
    .Y(_00805_),
    .B1(net2422));
 sg13g2_o21ai_1 _14275_ (.B1(net5152),
    .Y(_06132_),
    .A1(net5143),
    .A2(\i_wdt.counter[0] ));
 sg13g2_a21oi_1 _14276_ (.A1(_04282_),
    .A2(_06132_),
    .Y(_06133_),
    .B1(net1885));
 sg13g2_a221oi_1 _14277_ (.B2(net5152),
    .C1(_06133_),
    .B1(net1871),
    .A1(net2556),
    .Y(_06134_),
    .A2(net2064));
 sg13g2_nor2_1 _14278_ (.A(net2424),
    .B(net5153),
    .Y(_00806_));
 sg13g2_nand2_1 _14279_ (.Y(_06135_),
    .A(net4628),
    .B(net1871));
 sg13g2_xnor2_1 _14280_ (.Y(_06136_),
    .A(net4628),
    .B(_04282_));
 sg13g2_a22oi_1 _14281_ (.Y(_06137_),
    .B1(_04322_),
    .B2(_06136_),
    .A2(net2064),
    .A1(net2555));
 sg13g2_a21oi_1 _14282_ (.A1(_06135_),
    .A2(_06137_),
    .Y(_00807_),
    .B1(net2422));
 sg13g2_o21ai_1 _14283_ (.B1(net5084),
    .Y(_06138_),
    .A1(net4628),
    .A2(_04282_));
 sg13g2_a21oi_1 _14284_ (.A1(_04283_),
    .A2(_06138_),
    .Y(_06139_),
    .B1(net1885));
 sg13g2_a221oi_1 _14285_ (.B2(net5084),
    .C1(_06139_),
    .B1(net1871),
    .A1(net2554),
    .Y(_06140_),
    .A2(net2064));
 sg13g2_nor2_1 _14286_ (.A(net2423),
    .B(net5085),
    .Y(_00808_));
 sg13g2_nand2_1 _14287_ (.Y(_06141_),
    .A(net4717),
    .B(net1871));
 sg13g2_xnor2_1 _14288_ (.Y(_06142_),
    .A(net4717),
    .B(_04283_));
 sg13g2_a22oi_1 _14289_ (.Y(_06143_),
    .B1(_04322_),
    .B2(_06142_),
    .A2(net2065),
    .A1(net2553));
 sg13g2_a21oi_1 _14290_ (.A1(_06141_),
    .A2(_06143_),
    .Y(_00809_),
    .B1(net2424));
 sg13g2_o21ai_1 _14291_ (.B1(net5317),
    .Y(_06144_),
    .A1(\i_wdt.counter[5] ),
    .A2(_04283_));
 sg13g2_nor2b_1 _14292_ (.A(_04284_),
    .B_N(_06144_),
    .Y(_06145_));
 sg13g2_a22oi_1 _14293_ (.Y(_06146_),
    .B1(net1871),
    .B2(net5317),
    .A2(net2064),
    .A1(net2552));
 sg13g2_o21ai_1 _14294_ (.B1(_06146_),
    .Y(_06147_),
    .A1(net1885),
    .A2(_06145_));
 sg13g2_and2_1 _14295_ (.A(net2637),
    .B(_06147_),
    .X(_00810_));
 sg13g2_nand2_1 _14296_ (.Y(_06148_),
    .A(net4395),
    .B(net1871));
 sg13g2_xor2_1 _14297_ (.B(_04284_),
    .A(net4395),
    .X(_06149_));
 sg13g2_a22oi_1 _14298_ (.Y(_06150_),
    .B1(_04322_),
    .B2(_06149_),
    .A2(net2064),
    .A1(net2551));
 sg13g2_a21oi_1 _14299_ (.A1(_06148_),
    .A2(_06150_),
    .Y(_00811_),
    .B1(net2423));
 sg13g2_nand2b_1 _14300_ (.Y(_06151_),
    .B(net5011),
    .A_N(_04285_));
 sg13g2_a21o_1 _14301_ (.A2(_06151_),
    .A1(_04286_),
    .B1(net1886),
    .X(_06152_));
 sg13g2_a22oi_1 _14302_ (.Y(_06153_),
    .B1(net1871),
    .B2(net5011),
    .A2(net2065),
    .A1(net2549));
 sg13g2_a21oi_1 _14303_ (.A1(_06152_),
    .A2(_06153_),
    .Y(_00812_),
    .B1(net2415));
 sg13g2_xnor2_1 _14304_ (.Y(_06154_),
    .A(net5173),
    .B(_04286_));
 sg13g2_nand2_1 _14305_ (.Y(_06155_),
    .A(_04322_),
    .B(_06154_));
 sg13g2_a22oi_1 _14306_ (.Y(_06156_),
    .B1(net1871),
    .B2(net5173),
    .A2(net2063),
    .A1(net2548));
 sg13g2_a21oi_1 _14307_ (.A1(_06155_),
    .A2(_06156_),
    .Y(_00813_),
    .B1(net2422));
 sg13g2_o21ai_1 _14308_ (.B1(net5105),
    .Y(_06157_),
    .A1(\i_wdt.counter[9] ),
    .A2(_04286_));
 sg13g2_a21oi_1 _14309_ (.A1(_04287_),
    .A2(_06157_),
    .Y(_06158_),
    .B1(net1886));
 sg13g2_a221oi_1 _14310_ (.B2(net5105),
    .C1(_06158_),
    .B1(net1872),
    .A1(net4958),
    .Y(_06159_),
    .A2(net2063));
 sg13g2_nor2_1 _14311_ (.A(net2423),
    .B(net5106),
    .Y(_00814_));
 sg13g2_nand2_1 _14312_ (.Y(_06160_),
    .A(net5136),
    .B(_04287_));
 sg13g2_a21oi_1 _14313_ (.A1(_04288_),
    .A2(_06160_),
    .Y(_06161_),
    .B1(net1885));
 sg13g2_a221oi_1 _14314_ (.B2(net5136),
    .C1(_06161_),
    .B1(net1872),
    .A1(net5104),
    .Y(_06162_),
    .A2(net2063));
 sg13g2_nor2_1 _14315_ (.A(net2415),
    .B(_06162_),
    .Y(_00815_));
 sg13g2_or3_1 _14316_ (.A(net5304),
    .B(_04288_),
    .C(net1885),
    .X(_06163_));
 sg13g2_nor2_1 _14317_ (.A(net5304),
    .B(net2063),
    .Y(_06164_));
 sg13g2_a21oi_1 _14318_ (.A1(_01780_),
    .A2(net2063),
    .Y(_06165_),
    .B1(_06164_));
 sg13g2_o21ai_1 _14319_ (.B1(_06165_),
    .Y(_06166_),
    .A1(_04288_),
    .A2(net1885));
 sg13g2_a21oi_1 _14320_ (.A1(_06163_),
    .A2(_06166_),
    .Y(_00816_),
    .B1(net2422));
 sg13g2_nand2_1 _14321_ (.Y(_06167_),
    .A(_01793_),
    .B(net2063));
 sg13g2_o21ai_1 _14322_ (.B1(_06167_),
    .Y(_06168_),
    .A1(net5102),
    .A2(net2063));
 sg13g2_mux2_1 _14323_ (.A0(net5102),
    .A1(_06168_),
    .S(_06163_),
    .X(_06169_));
 sg13g2_nor2_1 _14324_ (.A(net2422),
    .B(net5103),
    .Y(_00817_));
 sg13g2_nor2_1 _14325_ (.A(net5210),
    .B(net2063),
    .Y(_06170_));
 sg13g2_a21oi_1 _14326_ (.A1(_01792_),
    .A2(net2064),
    .Y(_06171_),
    .B1(_06170_));
 sg13g2_o21ai_1 _14327_ (.B1(_06171_),
    .Y(_06172_),
    .A1(net5102),
    .A2(_06163_));
 sg13g2_nand2_1 _14328_ (.Y(_06173_),
    .A(_04289_),
    .B(_04304_));
 sg13g2_nand2_1 _14329_ (.Y(_06174_),
    .A(net5211),
    .B(_04322_));
 sg13g2_a21oi_1 _14330_ (.A1(_06172_),
    .A2(_06174_),
    .Y(_00818_),
    .B1(net2422));
 sg13g2_xor2_1 _14331_ (.B(_06173_),
    .A(net5157),
    .X(_06175_));
 sg13g2_nand3_1 _14332_ (.B(net2638),
    .C(net2066),
    .A(net4979),
    .Y(_06176_));
 sg13g2_o21ai_1 _14333_ (.B1(_06176_),
    .Y(_00819_),
    .A1(_06127_),
    .A2(net5158));
 sg13g2_nand2_1 _14334_ (.Y(_06177_),
    .A(net5117),
    .B(_04290_));
 sg13g2_a21oi_1 _14335_ (.A1(_04291_),
    .A2(_06177_),
    .Y(_06178_),
    .B1(net1885));
 sg13g2_a221oi_1 _14336_ (.B2(net5117),
    .C1(_06178_),
    .B1(net1872),
    .A1(net4892),
    .Y(_06179_),
    .A2(net2066));
 sg13g2_nor2_1 _14337_ (.A(net2422),
    .B(_06179_),
    .Y(_00820_));
 sg13g2_o21ai_1 _14338_ (.B1(net4817),
    .Y(_06180_),
    .A1(_04291_),
    .A2(_04303_));
 sg13g2_nor3_1 _14339_ (.A(net4817),
    .B(_04291_),
    .C(_04303_),
    .Y(_06181_));
 sg13g2_nor2_1 _14340_ (.A(net2066),
    .B(_06181_),
    .Y(_06182_));
 sg13g2_a22oi_1 _14341_ (.Y(_00821_),
    .B1(net4818),
    .B2(_06182_),
    .A2(_06127_),
    .A1(_04476_));
 sg13g2_or3_1 _14342_ (.A(_04292_),
    .B(_04303_),
    .C(net2066),
    .X(_06183_));
 sg13g2_a22oi_1 _14343_ (.Y(_06184_),
    .B1(_06182_),
    .B2(net5027),
    .A2(net2066),
    .A1(net4877));
 sg13g2_a21oi_1 _14344_ (.A1(_06183_),
    .A2(_06184_),
    .Y(_00822_),
    .B1(net2423));
 sg13g2_o21ai_1 _14345_ (.B1(net4702),
    .Y(_06185_),
    .A1(_04292_),
    .A2(_04303_));
 sg13g2_nor3_2 _14346_ (.A(net4702),
    .B(_04292_),
    .C(_04303_),
    .Y(_06186_));
 sg13g2_nor2_1 _14347_ (.A(net2068),
    .B(_06186_),
    .Y(_06187_));
 sg13g2_a221oi_1 _14348_ (.B2(_06187_),
    .C1(net2420),
    .B1(_06185_),
    .A1(_01836_),
    .Y(_00823_),
    .A2(net2068));
 sg13g2_nand2b_1 _14349_ (.Y(_06188_),
    .B(_06186_),
    .A_N(net5006));
 sg13g2_nand2b_1 _14350_ (.Y(_06189_),
    .B(_04321_),
    .A_N(_06188_));
 sg13g2_a22oi_1 _14351_ (.Y(_06190_),
    .B1(_06187_),
    .B2(net5006),
    .A2(net2068),
    .A1(net4994));
 sg13g2_a21oi_1 _14352_ (.A1(_06189_),
    .A2(_06190_),
    .Y(_00824_),
    .B1(net2421));
 sg13g2_nand2_1 _14353_ (.Y(_06191_),
    .A(net4663),
    .B(_06188_));
 sg13g2_nor2_1 _14354_ (.A(net4663),
    .B(_06188_),
    .Y(_06192_));
 sg13g2_nor2_1 _14355_ (.A(net2067),
    .B(_06192_),
    .Y(_06193_));
 sg13g2_a221oi_1 _14356_ (.B2(_06193_),
    .C1(net2421),
    .B1(net4664),
    .A1(_01832_),
    .Y(_00825_),
    .A2(net2067));
 sg13g2_nor4_1 _14357_ (.A(net5123),
    .B(net4663),
    .C(net2068),
    .D(_06188_),
    .Y(_06194_));
 sg13g2_a221oi_1 _14358_ (.B2(net5123),
    .C1(_06194_),
    .B1(_06193_),
    .A1(net4905),
    .Y(_06195_),
    .A2(_04319_));
 sg13g2_nor2_1 _14359_ (.A(net2420),
    .B(_06195_),
    .Y(_00826_));
 sg13g2_nor4_1 _14360_ (.A(_01957_),
    .B(net5123),
    .C(net4663),
    .D(net5006),
    .Y(_06196_));
 sg13g2_a21oi_1 _14361_ (.A1(_06186_),
    .A2(_06196_),
    .Y(_06197_),
    .B1(net2068));
 sg13g2_o21ai_1 _14362_ (.B1(_06197_),
    .Y(_06198_),
    .A1(net5125),
    .A2(_06194_));
 sg13g2_nand2_1 _14363_ (.Y(_06199_),
    .A(net4928),
    .B(net2067));
 sg13g2_a21oi_1 _14364_ (.A1(_06198_),
    .A2(_06199_),
    .Y(_00827_),
    .B1(net2421));
 sg13g2_nand2_1 _14365_ (.Y(_06200_),
    .A(_04293_),
    .B(_06186_));
 sg13g2_nand2_1 _14366_ (.Y(_06201_),
    .A(net4236),
    .B(_06200_));
 sg13g2_or2_1 _14367_ (.X(_06202_),
    .B(_06200_),
    .A(net4236));
 sg13g2_and2_1 _14368_ (.A(_04321_),
    .B(_06202_),
    .X(_06203_));
 sg13g2_a221oi_1 _14369_ (.B2(_06203_),
    .C1(net2420),
    .B1(net4237),
    .A1(_01826_),
    .Y(_00828_),
    .A2(net2067));
 sg13g2_nand2_1 _14370_ (.Y(_06204_),
    .A(net4265),
    .B(_06202_));
 sg13g2_nor2_1 _14371_ (.A(net4265),
    .B(_06202_),
    .Y(_06205_));
 sg13g2_nor2_1 _14372_ (.A(net2067),
    .B(_06205_),
    .Y(_06206_));
 sg13g2_a22oi_1 _14373_ (.Y(_00829_),
    .B1(_06204_),
    .B2(_06206_),
    .A2(_06127_),
    .A1(_04505_));
 sg13g2_o21ai_1 _14374_ (.B1(net4432),
    .Y(_06207_),
    .A1(net4265),
    .A2(_06202_));
 sg13g2_a21oi_1 _14375_ (.A1(_01956_),
    .A2(_06205_),
    .Y(_06208_),
    .B1(net2067));
 sg13g2_a221oi_1 _14376_ (.B2(_06208_),
    .C1(net2420),
    .B1(_06207_),
    .A1(_01822_),
    .Y(_00830_),
    .A2(net2067));
 sg13g2_nand2_1 _14377_ (.Y(_06209_),
    .A(_01820_),
    .B(net2067));
 sg13g2_a21oi_1 _14378_ (.A1(net4869),
    .A2(_04321_),
    .Y(_06210_),
    .B1(_06208_));
 sg13g2_a22oi_1 _14379_ (.Y(_06211_),
    .B1(_06209_),
    .B2(_06210_),
    .A2(_06208_),
    .A1(net4869));
 sg13g2_nor2_1 _14380_ (.A(net2420),
    .B(net4870),
    .Y(_00831_));
 sg13g2_nand2b_1 _14381_ (.Y(_06212_),
    .B(net4893),
    .A_N(_06210_));
 sg13g2_nor2_1 _14382_ (.A(_04297_),
    .B(net1886),
    .Y(_06213_));
 sg13g2_a21oi_1 _14383_ (.A1(\data_to_write[28] ),
    .A2(net2069),
    .Y(_06214_),
    .B1(_06213_));
 sg13g2_a21oi_1 _14384_ (.A1(_06212_),
    .A2(_06214_),
    .Y(_00832_),
    .B1(net2420));
 sg13g2_mux2_1 _14385_ (.A0(net5215),
    .A1(net5055),
    .S(net2069),
    .X(_06215_));
 sg13g2_nand3b_1 _14386_ (.B(_06215_),
    .C(net2640),
    .Y(_06216_),
    .A_N(_06213_));
 sg13g2_or3_1 _14387_ (.A(net5215),
    .B(_04297_),
    .C(_04303_),
    .X(_06217_));
 sg13g2_o21ai_1 _14388_ (.B1(_06216_),
    .Y(_00833_),
    .A1(_06127_),
    .A2(_06217_));
 sg13g2_nand3_1 _14389_ (.B(_04321_),
    .C(_06217_),
    .A(net4346),
    .Y(_06218_));
 sg13g2_a22oi_1 _14390_ (.Y(_06219_),
    .B1(_04322_),
    .B2(_04299_),
    .A2(net2069),
    .A1(\data_to_write[30] ));
 sg13g2_a21oi_1 _14391_ (.A1(net4347),
    .A2(_06219_),
    .Y(_00834_),
    .B1(net2419));
 sg13g2_nand2_1 _14392_ (.Y(_06220_),
    .A(\data_to_write[31] ),
    .B(net2066));
 sg13g2_nand2_1 _14393_ (.Y(_06221_),
    .A(net4391),
    .B(_04321_));
 sg13g2_a221oi_1 _14394_ (.B2(_06221_),
    .C1(net2419),
    .B1(_06220_),
    .A1(_04299_),
    .Y(_00835_),
    .A2(_04322_));
 sg13g2_nand2_1 _14395_ (.Y(_06222_),
    .A(net4940),
    .B(_03448_));
 sg13g2_o21ai_1 _14396_ (.B1(net4715),
    .Y(_06223_),
    .A1(net4762),
    .A2(net4021));
 sg13g2_nand4_1 _14397_ (.B(_03449_),
    .C(_06222_),
    .A(net2632),
    .Y(_00836_),
    .D(_06223_));
 sg13g2_nand2_1 _14398_ (.Y(_06224_),
    .A(net2326),
    .B(net2087));
 sg13g2_a21oi_1 _14399_ (.A1(net2326),
    .A2(net2085),
    .Y(_06225_),
    .B1(net2415));
 sg13g2_nand2_2 _14400_ (.Y(_06226_),
    .A(net2638),
    .B(net2001));
 sg13g2_xnor2_1 _14401_ (.Y(_06227_),
    .A(net4534),
    .B(net2302));
 sg13g2_nor2_1 _14402_ (.A(net1953),
    .B(_06227_),
    .Y(_00837_));
 sg13g2_a21oi_1 _14403_ (.A1(\i_rtc.us_count[0] ),
    .A2(net2302),
    .Y(_06228_),
    .B1(net3767));
 sg13g2_nand2_1 _14404_ (.Y(_06229_),
    .A(\i_rtc.us_count[1] ),
    .B(\i_rtc.us_count[0] ));
 sg13g2_and3_2 _14405_ (.X(_06230_),
    .A(net3767),
    .B(\i_rtc.us_count[0] ),
    .C(net2302));
 sg13g2_nor3_1 _14406_ (.A(net1953),
    .B(net3768),
    .C(_06230_),
    .Y(_00838_));
 sg13g2_o21ai_1 _14407_ (.B1(net1999),
    .Y(_06231_),
    .A1(net3521),
    .A2(_06230_));
 sg13g2_a21oi_1 _14408_ (.A1(net3521),
    .A2(_06230_),
    .Y(_00839_),
    .B1(_06231_));
 sg13g2_and3_2 _14409_ (.X(_06232_),
    .A(net3605),
    .B(net3521),
    .C(_06230_));
 sg13g2_a21oi_1 _14410_ (.A1(net3521),
    .A2(_06230_),
    .Y(_06233_),
    .B1(net3605));
 sg13g2_nor3_1 _14411_ (.A(net1954),
    .B(_06232_),
    .C(net3606),
    .Y(_00840_));
 sg13g2_o21ai_1 _14412_ (.B1(net1999),
    .Y(_06234_),
    .A1(net4076),
    .A2(_06232_));
 sg13g2_a21oi_1 _14413_ (.A1(net4076),
    .A2(_06232_),
    .Y(_00841_),
    .B1(_06234_));
 sg13g2_a21oi_1 _14414_ (.A1(net4076),
    .A2(_06232_),
    .Y(_06235_),
    .B1(net4293));
 sg13g2_and3_1 _14415_ (.X(_06236_),
    .A(net4293),
    .B(net4076),
    .C(_06232_));
 sg13g2_nor3_1 _14416_ (.A(net1954),
    .B(_06235_),
    .C(_06236_),
    .Y(_00842_));
 sg13g2_nand2b_1 _14417_ (.Y(_06237_),
    .B(\i_rtc.us_count[14] ),
    .A_N(\i_rtc.us_count[15] ));
 sg13g2_nand2_1 _14418_ (.Y(_06238_),
    .A(\i_rtc.us_count[19] ),
    .B(\i_rtc.us_count[18] ));
 sg13g2_nand4_1 _14419_ (.B(\i_rtc.us_count[16] ),
    .C(\i_rtc.us_count[5] ),
    .A(\i_rtc.us_count[17] ),
    .Y(_06239_),
    .D(\i_rtc.us_count[4] ));
 sg13g2_nand2b_1 _14420_ (.Y(_06240_),
    .B(\i_rtc.us_count[9] ),
    .A_N(\i_rtc.us_count[8] ));
 sg13g2_nor2_1 _14421_ (.A(\i_rtc.us_count[7] ),
    .B(\i_rtc.us_count[6] ),
    .Y(_06241_));
 sg13g2_nor4_1 _14422_ (.A(\i_rtc.us_count[13] ),
    .B(\i_rtc.us_count[12] ),
    .C(\i_rtc.us_count[11] ),
    .D(\i_rtc.us_count[10] ),
    .Y(_06242_));
 sg13g2_nand3b_1 _14423_ (.B(_06241_),
    .C(_06242_),
    .Y(_06243_),
    .A_N(_06240_));
 sg13g2_nor4_1 _14424_ (.A(_06237_),
    .B(_06238_),
    .C(_06239_),
    .D(_06243_),
    .Y(_06244_));
 sg13g2_and4_1 _14425_ (.A(\i_rtc.us_count[19] ),
    .B(\i_rtc.us_count[18] ),
    .C(\i_rtc.us_count[17] ),
    .D(\i_rtc.us_count[16] ),
    .X(_06245_));
 sg13g2_and4_1 _14426_ (.A(\i_rtc.us_count[5] ),
    .B(\i_rtc.us_count[4] ),
    .C(_06241_),
    .D(_06245_),
    .X(_06246_));
 sg13g2_or3_1 _14427_ (.A(\i_rtc.us_count[11] ),
    .B(\i_rtc.us_count[10] ),
    .C(_06240_),
    .X(_06247_));
 sg13g2_nor4_1 _14428_ (.A(\i_rtc.us_count[13] ),
    .B(\i_rtc.us_count[12] ),
    .C(_06237_),
    .D(_06247_),
    .Y(_06248_));
 sg13g2_nor4_1 _14429_ (.A(\i_rtc.us_count[7] ),
    .B(\i_rtc.us_count[6] ),
    .C(_06229_),
    .D(_06247_),
    .Y(_06249_));
 sg13g2_nand4_1 _14430_ (.B(\i_rtc.us_count[4] ),
    .C(\i_rtc.us_count[3] ),
    .A(\i_rtc.us_count[5] ),
    .Y(_06250_),
    .D(\i_rtc.us_count[2] ));
 sg13g2_nor4_1 _14431_ (.A(\i_rtc.us_count[13] ),
    .B(\i_rtc.us_count[12] ),
    .C(_06237_),
    .D(_06250_),
    .Y(_06251_));
 sg13g2_nand4_1 _14432_ (.B(_06245_),
    .C(_06249_),
    .A(net2302),
    .Y(_06252_),
    .D(_06251_));
 sg13g2_nand2_2 _14433_ (.Y(_06253_),
    .A(net1999),
    .B(_06252_));
 sg13g2_inv_1 _14434_ (.Y(_06254_),
    .A(_06253_));
 sg13g2_and4_1 _14435_ (.A(net4415),
    .B(net4293),
    .C(net4076),
    .D(_06232_),
    .X(_06255_));
 sg13g2_nor2_1 _14436_ (.A(net4415),
    .B(_06236_),
    .Y(_06256_));
 sg13g2_nor3_1 _14437_ (.A(_06253_),
    .B(_06255_),
    .C(_06256_),
    .Y(_00843_));
 sg13g2_xnor2_1 _14438_ (.Y(_06257_),
    .A(net4861),
    .B(_06255_));
 sg13g2_nor2_1 _14439_ (.A(net1954),
    .B(_06257_),
    .Y(_00844_));
 sg13g2_a21oi_1 _14440_ (.A1(\i_rtc.us_count[7] ),
    .A2(_06255_),
    .Y(_06258_),
    .B1(net4012));
 sg13g2_and4_1 _14441_ (.A(net4012),
    .B(\i_rtc.us_count[7] ),
    .C(net4415),
    .D(_06236_),
    .X(_06259_));
 sg13g2_nor3_1 _14442_ (.A(net1953),
    .B(net4013),
    .C(_06259_),
    .Y(_00845_));
 sg13g2_nor2_1 _14443_ (.A(net4500),
    .B(_06259_),
    .Y(_06260_));
 sg13g2_and4_1 _14444_ (.A(net4500),
    .B(net4012),
    .C(\i_rtc.us_count[7] ),
    .D(_06255_),
    .X(_06261_));
 sg13g2_nor3_1 _14445_ (.A(_06253_),
    .B(net4501),
    .C(_06261_),
    .Y(_00846_));
 sg13g2_nor2_1 _14446_ (.A(net4580),
    .B(_06261_),
    .Y(_06262_));
 sg13g2_and2_1 _14447_ (.A(net4580),
    .B(_06261_),
    .X(_06263_));
 sg13g2_nor3_1 _14448_ (.A(net1953),
    .B(net4581),
    .C(_06263_),
    .Y(_00847_));
 sg13g2_xnor2_1 _14449_ (.Y(_06264_),
    .A(net4754),
    .B(_06263_));
 sg13g2_nor2_1 _14450_ (.A(net1953),
    .B(_06264_),
    .Y(_00848_));
 sg13g2_a21oi_1 _14451_ (.A1(\i_rtc.us_count[11] ),
    .A2(_06263_),
    .Y(_06265_),
    .B1(net4216));
 sg13g2_and3_1 _14452_ (.X(_06266_),
    .A(net4216),
    .B(net5386),
    .C(_06263_));
 sg13g2_nor3_1 _14453_ (.A(net1953),
    .B(net4217),
    .C(_06266_),
    .Y(_00849_));
 sg13g2_nor2_1 _14454_ (.A(net4704),
    .B(_06266_),
    .Y(_06267_));
 sg13g2_and2_1 _14455_ (.A(net4704),
    .B(_06266_),
    .X(_06268_));
 sg13g2_nor3_1 _14456_ (.A(net1953),
    .B(net4705),
    .C(_06268_),
    .Y(_00850_));
 sg13g2_and2_1 _14457_ (.A(net4863),
    .B(_06268_),
    .X(_06269_));
 sg13g2_o21ai_1 _14458_ (.B1(_06254_),
    .Y(_06270_),
    .A1(net4863),
    .A2(_06268_));
 sg13g2_nor2_1 _14459_ (.A(_06269_),
    .B(net4864),
    .Y(_00851_));
 sg13g2_nor2_1 _14460_ (.A(net4305),
    .B(_06269_),
    .Y(_06271_));
 sg13g2_and2_1 _14461_ (.A(net4305),
    .B(_06269_),
    .X(_06272_));
 sg13g2_nor3_1 _14462_ (.A(net1953),
    .B(net4306),
    .C(_06272_),
    .Y(_00852_));
 sg13g2_nor2_1 _14463_ (.A(net4803),
    .B(_06272_),
    .Y(_06273_));
 sg13g2_and2_1 _14464_ (.A(net4803),
    .B(_06272_),
    .X(_06274_));
 sg13g2_nor3_1 _14465_ (.A(_06253_),
    .B(net4804),
    .C(_06274_),
    .Y(_00853_));
 sg13g2_o21ai_1 _14466_ (.B1(_06254_),
    .Y(_06275_),
    .A1(net3607),
    .A2(_06274_));
 sg13g2_a21oi_1 _14467_ (.A1(net3607),
    .A2(_06274_),
    .Y(_00854_),
    .B1(_06275_));
 sg13g2_a21oi_1 _14468_ (.A1(net3607),
    .A2(_06274_),
    .Y(_06276_),
    .B1(net4092));
 sg13g2_and3_1 _14469_ (.X(_06277_),
    .A(net4092),
    .B(net3607),
    .C(_06274_));
 sg13g2_nor3_1 _14470_ (.A(_06253_),
    .B(net4093),
    .C(_06277_),
    .Y(_00855_));
 sg13g2_xnor2_1 _14471_ (.Y(_06278_),
    .A(net4680),
    .B(_06277_));
 sg13g2_nor2_1 _14472_ (.A(_06253_),
    .B(_06278_),
    .Y(_00856_));
 sg13g2_and4_1 _14473_ (.A(\i_rtc.seconds_out[0] ),
    .B(_06232_),
    .C(_06246_),
    .D(_06248_),
    .X(_06279_));
 sg13g2_xnor2_1 _14474_ (.Y(_06280_),
    .A(net5362),
    .B(_06252_));
 sg13g2_nand2_1 _14475_ (.Y(_06281_),
    .A(net2000),
    .B(_06280_));
 sg13g2_nor2_1 _14476_ (.A(net2415),
    .B(_06224_),
    .Y(_06282_));
 sg13g2_o21ai_1 _14477_ (.B1(_06281_),
    .Y(_00857_),
    .A1(_04425_),
    .A2(net2001));
 sg13g2_and4_1 _14478_ (.A(\i_rtc.seconds_out[1] ),
    .B(\i_rtc.seconds_out[0] ),
    .C(_06232_),
    .D(_06244_),
    .X(_06283_));
 sg13g2_nand2_1 _14479_ (.Y(_06284_),
    .A(\i_rtc.seconds_out[1] ),
    .B(\i_rtc.seconds_out[0] ));
 sg13g2_nor2_1 _14480_ (.A(_06252_),
    .B(_06284_),
    .Y(_06285_));
 sg13g2_xnor2_1 _14481_ (.Y(_06286_),
    .A(net5320),
    .B(_06279_));
 sg13g2_nand2_1 _14482_ (.Y(_06287_),
    .A(net2558),
    .B(net1946));
 sg13g2_o21ai_1 _14483_ (.B1(_06287_),
    .Y(_00858_),
    .A1(net1951),
    .A2(_06286_));
 sg13g2_and3_2 _14484_ (.X(_06288_),
    .A(net5076),
    .B(\i_rtc.seconds_out[1] ),
    .C(_06279_));
 sg13g2_xnor2_1 _14485_ (.Y(_06289_),
    .A(net5076),
    .B(_06285_));
 sg13g2_nand2_1 _14486_ (.Y(_06290_),
    .A(net2556),
    .B(net1945));
 sg13g2_o21ai_1 _14487_ (.B1(_06290_),
    .Y(_00859_),
    .A1(net1950),
    .A2(net5077));
 sg13g2_nand2_1 _14488_ (.Y(_06291_),
    .A(net5162),
    .B(_06288_));
 sg13g2_xnor2_1 _14489_ (.Y(_06292_),
    .A(net5162),
    .B(_06288_));
 sg13g2_nand2_1 _14490_ (.Y(_06293_),
    .A(net2555),
    .B(net1945));
 sg13g2_o21ai_1 _14491_ (.B1(_06293_),
    .Y(_00860_),
    .A1(net1950),
    .A2(net5163));
 sg13g2_and4_1 _14492_ (.A(net5179),
    .B(net5162),
    .C(net5076),
    .D(_06283_),
    .X(_06294_));
 sg13g2_and4_1 _14493_ (.A(net5179),
    .B(net5162),
    .C(net5076),
    .D(_06285_),
    .X(_06295_));
 sg13g2_xor2_1 _14494_ (.B(_06291_),
    .A(net5179),
    .X(_06296_));
 sg13g2_a22oi_1 _14495_ (.Y(_00861_),
    .B1(_06296_),
    .B2(net2001),
    .A2(net1950),
    .A1(_04434_));
 sg13g2_nand4_1 _14496_ (.B(net5179),
    .C(net5162),
    .A(net5258),
    .Y(_06297_),
    .D(_06288_));
 sg13g2_o21ai_1 _14497_ (.B1(_06297_),
    .Y(_06298_),
    .A1(net5258),
    .A2(_06294_));
 sg13g2_a22oi_1 _14498_ (.Y(_00862_),
    .B1(_06298_),
    .B2(net2001),
    .A2(net1950),
    .A1(_04438_));
 sg13g2_nand3_1 _14499_ (.B(net5258),
    .C(_06295_),
    .A(net5309),
    .Y(_06299_));
 sg13g2_xnor2_1 _14500_ (.Y(_06300_),
    .A(_01955_),
    .B(_06297_));
 sg13g2_a22oi_1 _14501_ (.Y(_00863_),
    .B1(_06300_),
    .B2(net2001),
    .A2(net1951),
    .A1(_04441_));
 sg13g2_and4_1 _14502_ (.A(\i_rtc.seconds_out[7] ),
    .B(\i_rtc.seconds_out[6] ),
    .C(net5258),
    .D(_06294_),
    .X(_06301_));
 sg13g2_nor3_1 _14503_ (.A(_01954_),
    .B(_01955_),
    .C(_06297_),
    .Y(_06302_));
 sg13g2_nor2_1 _14504_ (.A(_01954_),
    .B(_06299_),
    .Y(_06303_));
 sg13g2_xnor2_1 _14505_ (.Y(_06304_),
    .A(_01954_),
    .B(_06299_));
 sg13g2_a22oi_1 _14506_ (.Y(_00864_),
    .B1(_06304_),
    .B2(net2001),
    .A2(net1951),
    .A1(_04444_));
 sg13g2_o21ai_1 _14507_ (.B1(net2000),
    .Y(_06305_),
    .A1(net5197),
    .A2(_06301_));
 sg13g2_a21oi_1 _14508_ (.A1(net5197),
    .A2(_06302_),
    .Y(_06306_),
    .B1(_06305_));
 sg13g2_a21o_1 _14509_ (.A2(net1946),
    .A1(net2549),
    .B1(net5198),
    .X(_00865_));
 sg13g2_a21oi_1 _14510_ (.A1(net5197),
    .A2(_06301_),
    .Y(_06307_),
    .B1(net5288));
 sg13g2_nor2_1 _14511_ (.A(net1951),
    .B(_06307_),
    .Y(_06308_));
 sg13g2_nand3_1 _14512_ (.B(net5197),
    .C(_06301_),
    .A(net5288),
    .Y(_06309_));
 sg13g2_inv_1 _14513_ (.Y(_06310_),
    .A(_06309_));
 sg13g2_a22oi_1 _14514_ (.Y(_06311_),
    .B1(_06308_),
    .B2(net5289),
    .A2(net1946),
    .A1(net2548));
 sg13g2_inv_1 _14515_ (.Y(_00866_),
    .A(_06311_));
 sg13g2_o21ai_1 _14516_ (.B1(net2000),
    .Y(_06312_),
    .A1(net5231),
    .A2(_06310_));
 sg13g2_and4_1 _14517_ (.A(net5231),
    .B(\i_rtc.seconds_out[9] ),
    .C(net5197),
    .D(_06302_),
    .X(_06313_));
 sg13g2_or2_1 _14518_ (.X(_06314_),
    .B(net2001),
    .A(_04457_));
 sg13g2_and4_1 _14519_ (.A(\i_rtc.seconds_out[10] ),
    .B(\i_rtc.seconds_out[9] ),
    .C(\i_rtc.seconds_out[8] ),
    .D(_06303_),
    .X(_06315_));
 sg13g2_o21ai_1 _14520_ (.B1(_06314_),
    .Y(_00867_),
    .A1(net5232),
    .A2(_06313_));
 sg13g2_and2_1 _14521_ (.A(net5181),
    .B(_06313_),
    .X(_06316_));
 sg13g2_o21ai_1 _14522_ (.B1(net2000),
    .Y(_06317_),
    .A1(net5181),
    .A2(_06315_));
 sg13g2_nand2_1 _14523_ (.Y(_06318_),
    .A(net5104),
    .B(net1945));
 sg13g2_o21ai_1 _14524_ (.B1(_06318_),
    .Y(_00868_),
    .A1(_06316_),
    .A2(net5182));
 sg13g2_o21ai_1 _14525_ (.B1(net2000),
    .Y(_06319_),
    .A1(net5293),
    .A2(_06316_));
 sg13g2_nand4_1 _14526_ (.B(net5181),
    .C(net5231),
    .A(net5293),
    .Y(_06320_),
    .D(_06310_));
 sg13g2_nand2b_1 _14527_ (.Y(_06321_),
    .B(_06320_),
    .A_N(_06319_));
 sg13g2_nand2_1 _14528_ (.Y(_06322_),
    .A(net2547),
    .B(net1945));
 sg13g2_nand2_1 _14529_ (.Y(_00869_),
    .A(_06321_),
    .B(_06322_));
 sg13g2_and2_1 _14530_ (.A(_01953_),
    .B(_06320_),
    .X(_06323_));
 sg13g2_nor2_1 _14531_ (.A(_01953_),
    .B(_06320_),
    .Y(_06324_));
 sg13g2_and4_1 _14532_ (.A(net5239),
    .B(\i_rtc.seconds_out[12] ),
    .C(net5181),
    .D(_06315_),
    .X(_06325_));
 sg13g2_nor3_1 _14533_ (.A(net1950),
    .B(net5240),
    .C(_06325_),
    .Y(_06326_));
 sg13g2_a21o_1 _14534_ (.A2(net1945),
    .A1(net5053),
    .B1(net5241),
    .X(_00870_));
 sg13g2_nor2_1 _14535_ (.A(net5245),
    .B(_06324_),
    .Y(_06327_));
 sg13g2_and2_1 _14536_ (.A(net5245),
    .B(_06324_),
    .X(_06328_));
 sg13g2_nor3_1 _14537_ (.A(net1950),
    .B(net5246),
    .C(_06328_),
    .Y(_06329_));
 sg13g2_a21o_1 _14538_ (.A2(net1945),
    .A1(net4962),
    .B1(_06329_),
    .X(_00871_));
 sg13g2_a21oi_1 _14539_ (.A1(net5140),
    .A2(_06328_),
    .Y(_06330_),
    .B1(net1950));
 sg13g2_o21ai_1 _14540_ (.B1(_06330_),
    .Y(_06331_),
    .A1(net5140),
    .A2(_06328_));
 sg13g2_nand2_1 _14541_ (.Y(_06332_),
    .A(net4979),
    .B(net1945));
 sg13g2_nand2_1 _14542_ (.Y(_00872_),
    .A(net5141),
    .B(_06332_));
 sg13g2_a21oi_1 _14543_ (.A1(\i_rtc.seconds_out[15] ),
    .A2(_06328_),
    .Y(_06333_),
    .B1(net5114));
 sg13g2_and3_2 _14544_ (.X(_06334_),
    .A(net5114),
    .B(\i_rtc.seconds_out[15] ),
    .C(_06328_));
 sg13g2_and4_1 _14545_ (.A(\i_rtc.seconds_out[16] ),
    .B(\i_rtc.seconds_out[15] ),
    .C(\i_rtc.seconds_out[14] ),
    .D(_06325_),
    .X(_06335_));
 sg13g2_nor3_1 _14546_ (.A(net1950),
    .B(net5115),
    .C(_06334_),
    .Y(_06336_));
 sg13g2_a21o_1 _14547_ (.A2(net1945),
    .A1(net4892),
    .B1(net5116),
    .X(_00873_));
 sg13g2_and2_1 _14548_ (.A(net5030),
    .B(_06334_),
    .X(_06337_));
 sg13g2_xnor2_1 _14549_ (.Y(_06338_),
    .A(net5030),
    .B(_06335_));
 sg13g2_a22oi_1 _14550_ (.Y(_00874_),
    .B1(net5031),
    .B2(net2001),
    .A2(net1951),
    .A1(_04476_));
 sg13g2_nand2_1 _14551_ (.Y(_06339_),
    .A(net5180),
    .B(_06337_));
 sg13g2_o21ai_1 _14552_ (.B1(net1999),
    .Y(_06340_),
    .A1(net5180),
    .A2(_06337_));
 sg13g2_nor2b_1 _14553_ (.A(_06340_),
    .B_N(_06339_),
    .Y(_06341_));
 sg13g2_a21o_1 _14554_ (.A2(net1947),
    .A1(net4877),
    .B1(_06341_),
    .X(_00875_));
 sg13g2_nor2_1 _14555_ (.A(_01952_),
    .B(_06339_),
    .Y(_06342_));
 sg13g2_a21oi_1 _14556_ (.A1(_01952_),
    .A2(_06339_),
    .Y(_06343_),
    .B1(net1952));
 sg13g2_and4_1 _14557_ (.A(net5056),
    .B(net5180),
    .C(net5030),
    .D(_06335_),
    .X(_06344_));
 sg13g2_nor2b_1 _14558_ (.A(_06342_),
    .B_N(net5057),
    .Y(_06345_));
 sg13g2_a21o_1 _14559_ (.A2(net1947),
    .A1(net4912),
    .B1(net5058),
    .X(_00876_));
 sg13g2_and2_1 _14560_ (.A(net5213),
    .B(_06342_),
    .X(_06346_));
 sg13g2_o21ai_1 _14561_ (.B1(net2000),
    .Y(_06347_),
    .A1(net5213),
    .A2(_06344_));
 sg13g2_nand2_1 _14562_ (.Y(_06348_),
    .A(net4994),
    .B(net1948));
 sg13g2_o21ai_1 _14563_ (.B1(_06348_),
    .Y(_00877_),
    .A1(_06346_),
    .A2(_06347_));
 sg13g2_a21oi_1 _14564_ (.A1(net5100),
    .A2(_06346_),
    .Y(_06349_),
    .B1(net1955));
 sg13g2_o21ai_1 _14565_ (.B1(_06349_),
    .Y(_06350_),
    .A1(net5100),
    .A2(_06346_));
 sg13g2_nand2_1 _14566_ (.Y(_06351_),
    .A(net4933),
    .B(net1948));
 sg13g2_nand2_1 _14567_ (.Y(_00878_),
    .A(net5101),
    .B(_06351_));
 sg13g2_a21oi_1 _14568_ (.A1(net5100),
    .A2(_06346_),
    .Y(_06352_),
    .B1(net5193));
 sg13g2_and3_1 _14569_ (.X(_06353_),
    .A(\i_rtc.seconds_out[22] ),
    .B(\i_rtc.seconds_out[21] ),
    .C(_06346_));
 sg13g2_and4_1 _14570_ (.A(\i_rtc.seconds_out[22] ),
    .B(\i_rtc.seconds_out[21] ),
    .C(\i_rtc.seconds_out[20] ),
    .D(_06344_),
    .X(_06354_));
 sg13g2_nor3_1 _14571_ (.A(net1955),
    .B(net5194),
    .C(_06354_),
    .Y(_06355_));
 sg13g2_a21o_1 _14572_ (.A2(net1948),
    .A1(net4905),
    .B1(net5195),
    .X(_00879_));
 sg13g2_o21ai_1 _14573_ (.B1(net2000),
    .Y(_06356_),
    .A1(net5150),
    .A2(_06354_));
 sg13g2_a21oi_1 _14574_ (.A1(net5150),
    .A2(_06354_),
    .Y(_06357_),
    .B1(_06356_));
 sg13g2_a21o_1 _14575_ (.A2(net1947),
    .A1(net4928),
    .B1(net5151),
    .X(_00880_));
 sg13g2_a21oi_1 _14576_ (.A1(\i_rtc.seconds_out[23] ),
    .A2(_06354_),
    .Y(_06358_),
    .B1(net4733));
 sg13g2_nand3_1 _14577_ (.B(net5150),
    .C(_06353_),
    .A(net4733),
    .Y(_06359_));
 sg13g2_nand2_1 _14578_ (.Y(_06360_),
    .A(net1999),
    .B(_06359_));
 sg13g2_nand2_1 _14579_ (.Y(_06361_),
    .A(\data_to_write[24] ),
    .B(net1947));
 sg13g2_o21ai_1 _14580_ (.B1(_06361_),
    .Y(_00881_),
    .A1(net4734),
    .A2(_06360_));
 sg13g2_and2_1 _14581_ (.A(_01951_),
    .B(_06359_),
    .X(_06362_));
 sg13g2_and4_1 _14582_ (.A(net5176),
    .B(net4733),
    .C(\i_rtc.seconds_out[23] ),
    .D(_06354_),
    .X(_06363_));
 sg13g2_nor3_1 _14583_ (.A(net1955),
    .B(_06362_),
    .C(_06363_),
    .Y(_06364_));
 sg13g2_a21o_1 _14584_ (.A2(net1948),
    .A1(net5071),
    .B1(net5177),
    .X(_00882_));
 sg13g2_nor3_2 _14585_ (.A(_01950_),
    .B(_01951_),
    .C(_06359_),
    .Y(_06365_));
 sg13g2_o21ai_1 _14586_ (.B1(net1999),
    .Y(_06366_),
    .A1(net5087),
    .A2(_06363_));
 sg13g2_nand2_1 _14587_ (.Y(_06367_),
    .A(net5054),
    .B(net1947));
 sg13g2_o21ai_1 _14588_ (.B1(_06367_),
    .Y(_00883_),
    .A1(_06365_),
    .A2(net5088));
 sg13g2_o21ai_1 _14589_ (.B1(net1999),
    .Y(_06368_),
    .A1(\i_rtc.seconds_out[27] ),
    .A2(_06365_));
 sg13g2_a21oi_1 _14590_ (.A1(\i_rtc.seconds_out[27] ),
    .A2(_06365_),
    .Y(_06369_),
    .B1(_06368_));
 sg13g2_a21o_1 _14591_ (.A2(net1947),
    .A1(net5079),
    .B1(_06369_),
    .X(_00884_));
 sg13g2_nand3_1 _14592_ (.B(\i_rtc.seconds_out[27] ),
    .C(_06365_),
    .A(\i_rtc.seconds_out[28] ),
    .Y(_06370_));
 sg13g2_a21oi_1 _14593_ (.A1(\i_rtc.seconds_out[27] ),
    .A2(_06365_),
    .Y(_06371_),
    .B1(net5276));
 sg13g2_and4_1 _14594_ (.A(net5276),
    .B(\i_rtc.seconds_out[27] ),
    .C(net5087),
    .D(_06363_),
    .X(_06372_));
 sg13g2_nor2_1 _14595_ (.A(net5277),
    .B(_06372_),
    .Y(_06373_));
 sg13g2_a22oi_1 _14596_ (.Y(_06374_),
    .B1(net5278),
    .B2(net1999),
    .A2(net1947),
    .A1(net4927));
 sg13g2_inv_1 _14597_ (.Y(_00885_),
    .A(_06374_));
 sg13g2_a21oi_1 _14598_ (.A1(_01949_),
    .A2(_06370_),
    .Y(_06375_),
    .B1(net1952));
 sg13g2_nand2_1 _14599_ (.Y(_06376_),
    .A(net5222),
    .B(_06372_));
 sg13g2_a22oi_1 _14600_ (.Y(_06377_),
    .B1(_06375_),
    .B2(net5223),
    .A2(net1947),
    .A1(net5055));
 sg13g2_inv_1 _14601_ (.Y(_00886_),
    .A(net5224));
 sg13g2_nand3_1 _14602_ (.B(\i_rtc.seconds_out[29] ),
    .C(_06372_),
    .A(\i_rtc.seconds_out[30] ),
    .Y(_06378_));
 sg13g2_xor2_1 _14603_ (.B(_06376_),
    .A(net5046),
    .X(_06379_));
 sg13g2_nand2_1 _14604_ (.Y(_06380_),
    .A(net5005),
    .B(net1949));
 sg13g2_o21ai_1 _14605_ (.B1(_06380_),
    .Y(_00887_),
    .A1(net1952),
    .A2(net5047));
 sg13g2_xor2_1 _14606_ (.B(_06378_),
    .A(\i_rtc.seconds_out[31] ),
    .X(_06381_));
 sg13g2_nand2_1 _14607_ (.Y(_06382_),
    .A(net5020),
    .B(net1949));
 sg13g2_o21ai_1 _14608_ (.B1(_06382_),
    .Y(_00888_),
    .A1(net1952),
    .A2(_06381_));
 sg13g2_nor2_2 _14609_ (.A(net5201),
    .B(_01810_),
    .Y(_06383_));
 sg13g2_nand2b_1 _14610_ (.Y(_06384_),
    .B(net5345),
    .A_N(net5201));
 sg13g2_nor3_2 _14611_ (.A(net4363),
    .B(net2307),
    .C(_06384_),
    .Y(_06385_));
 sg13g2_nand2_2 _14612_ (.Y(_06386_),
    .A(net2663),
    .B(net2220));
 sg13g2_inv_1 _14613_ (.Y(_00889_),
    .A(_06386_));
 sg13g2_nor4_2 _14614_ (.A(_01947_),
    .B(\i_seal.byte_idx[2] ),
    .C(\i_seal.byte_idx[1] ),
    .Y(_06387_),
    .D(net2493));
 sg13g2_inv_1 _14615_ (.Y(_06388_),
    .A(net2280));
 sg13g2_nand2_1 _14616_ (.Y(_06389_),
    .A(net4363),
    .B(net2309));
 sg13g2_nor2_1 _14617_ (.A(net2280),
    .B(_06389_),
    .Y(_06390_));
 sg13g2_a21oi_1 _14618_ (.A1(_01948_),
    .A2(net2307),
    .Y(_06391_),
    .B1(_06390_));
 sg13g2_nand3_1 _14619_ (.B(net2326),
    .C(_03465_),
    .A(net2558),
    .Y(_06392_));
 sg13g2_a21o_1 _14620_ (.A2(_06392_),
    .A1(_01810_),
    .B1(\i_seal.state[1] ),
    .X(_06393_));
 sg13g2_a22oi_1 _14621_ (.Y(_06394_),
    .B1(_06393_),
    .B2(net4363),
    .A2(_06391_),
    .A1(_06383_));
 sg13g2_nor2_1 _14622_ (.A(net2424),
    .B(net4364),
    .Y(_00890_));
 sg13g2_nor2_2 _14623_ (.A(net2339),
    .B(_06392_),
    .Y(_06395_));
 sg13g2_o21ai_1 _14624_ (.B1(_06383_),
    .Y(_06396_),
    .A1(_06388_),
    .A2(_06389_));
 sg13g2_nand4_1 _14625_ (.B(_02472_),
    .C(_03463_),
    .A(net2558),
    .Y(_06397_),
    .D(_03465_));
 sg13g2_o21ai_1 _14626_ (.B1(net1997),
    .Y(_06398_),
    .A1(_06389_),
    .A2(_06396_));
 sg13g2_o21ai_1 _14627_ (.B1(_06398_),
    .Y(_06399_),
    .A1(_01810_),
    .A2(net2493));
 sg13g2_o21ai_1 _14628_ (.B1(net5346),
    .Y(_06400_),
    .A1(net2493),
    .A2(_06398_));
 sg13g2_nor2_1 _14629_ (.A(net2424),
    .B(net5347),
    .Y(_00891_));
 sg13g2_o21ai_1 _14630_ (.B1(_06383_),
    .Y(_06401_),
    .A1(net5299),
    .A2(net2493));
 sg13g2_nand2_2 _14631_ (.Y(_06402_),
    .A(net5299),
    .B(net2493));
 sg13g2_nand2_1 _14632_ (.Y(_06403_),
    .A(_06398_),
    .B(_06401_));
 sg13g2_o21ai_1 _14633_ (.B1(_06403_),
    .Y(_06404_),
    .A1(net5299),
    .A2(_06398_));
 sg13g2_nor2b_1 _14634_ (.A(_06402_),
    .B_N(_06398_),
    .Y(_06405_));
 sg13g2_nor3_1 _14635_ (.A(net2424),
    .B(net5300),
    .C(_06405_),
    .Y(_00892_));
 sg13g2_nor2_1 _14636_ (.A(net5190),
    .B(_06405_),
    .Y(_06406_));
 sg13g2_nor2_2 _14637_ (.A(net2424),
    .B(net1944),
    .Y(_06407_));
 sg13g2_nand2_2 _14638_ (.Y(_06408_),
    .A(net2638),
    .B(net1998));
 sg13g2_a21o_1 _14639_ (.A2(_06405_),
    .A1(net5190),
    .B1(_06408_),
    .X(_06409_));
 sg13g2_nor2_1 _14640_ (.A(net5191),
    .B(_06409_),
    .Y(_00893_));
 sg13g2_nand2_2 _14641_ (.Y(_06410_),
    .A(_01947_),
    .B(\i_seal.byte_idx[2] ));
 sg13g2_nor2_2 _14642_ (.A(_06402_),
    .B(_06410_),
    .Y(_06411_));
 sg13g2_nand4_1 _14643_ (.B(_06383_),
    .C(_06398_),
    .A(net2663),
    .Y(_06412_),
    .D(net2219));
 sg13g2_o21ai_1 _14644_ (.B1(_06412_),
    .Y(_00894_),
    .A1(_01947_),
    .A2(_06409_));
 sg13g2_nand2b_1 _14645_ (.Y(_06413_),
    .B(net5201),
    .A_N(\i_seal.state[0] ));
 sg13g2_nor2_1 _14646_ (.A(net2307),
    .B(_06413_),
    .Y(_06414_));
 sg13g2_or2_1 _14647_ (.X(_06415_),
    .B(_06413_),
    .A(net2307));
 sg13g2_o21ai_1 _14648_ (.B1(net2643),
    .Y(_06416_),
    .A1(net4682),
    .A2(net2195));
 sg13g2_a21oi_1 _14649_ (.A1(_01763_),
    .A2(net2195),
    .Y(_00895_),
    .B1(_06416_));
 sg13g2_o21ai_1 _14650_ (.B1(net2644),
    .Y(_06417_),
    .A1(net4687),
    .A2(net2195));
 sg13g2_a21oi_1 _14651_ (.A1(_01762_),
    .A2(net2195),
    .Y(_00896_),
    .B1(_06417_));
 sg13g2_o21ai_1 _14652_ (.B1(net2644),
    .Y(_06418_),
    .A1(net4747),
    .A2(net2201));
 sg13g2_a21oi_1 _14653_ (.A1(_01761_),
    .A2(net2197),
    .Y(_00897_),
    .B1(_06418_));
 sg13g2_o21ai_1 _14654_ (.B1(net2644),
    .Y(_06419_),
    .A1(net4843),
    .A2(net2198));
 sg13g2_a21oi_1 _14655_ (.A1(_01760_),
    .A2(net2198),
    .Y(_00898_),
    .B1(_06419_));
 sg13g2_o21ai_1 _14656_ (.B1(net2644),
    .Y(_06420_),
    .A1(\i_seal.sealed_crc[4] ),
    .A2(net2197));
 sg13g2_a21oi_1 _14657_ (.A1(_01759_),
    .A2(net2198),
    .Y(_00899_),
    .B1(_06420_));
 sg13g2_o21ai_1 _14658_ (.B1(net2644),
    .Y(_06421_),
    .A1(net4527),
    .A2(net2197));
 sg13g2_a21oi_1 _14659_ (.A1(_01758_),
    .A2(net2197),
    .Y(_00900_),
    .B1(_06421_));
 sg13g2_o21ai_1 _14660_ (.B1(net2643),
    .Y(_06422_),
    .A1(net4586),
    .A2(net2195));
 sg13g2_a21oi_1 _14661_ (.A1(_01757_),
    .A2(net2196),
    .Y(_00901_),
    .B1(_06422_));
 sg13g2_o21ai_1 _14662_ (.B1(net2643),
    .Y(_06423_),
    .A1(net4529),
    .A2(net2195));
 sg13g2_a21oi_1 _14663_ (.A1(_01756_),
    .A2(net2196),
    .Y(_00902_),
    .B1(_06423_));
 sg13g2_o21ai_1 _14664_ (.B1(net2646),
    .Y(_06424_),
    .A1(\crc16_read[8] ),
    .A2(net2191));
 sg13g2_a21oi_1 _14665_ (.A1(_01946_),
    .A2(net2191),
    .Y(_00903_),
    .B1(_06424_));
 sg13g2_o21ai_1 _14666_ (.B1(net2661),
    .Y(_06425_),
    .A1(\crc16_read[9] ),
    .A2(net2192));
 sg13g2_a21oi_1 _14667_ (.A1(_01945_),
    .A2(net2192),
    .Y(_00904_),
    .B1(_06425_));
 sg13g2_o21ai_1 _14668_ (.B1(net2661),
    .Y(_06426_),
    .A1(\crc16_read[10] ),
    .A2(net2192));
 sg13g2_a21oi_1 _14669_ (.A1(_01944_),
    .A2(net2192),
    .Y(_00905_),
    .B1(_06426_));
 sg13g2_o21ai_1 _14670_ (.B1(net2647),
    .Y(_06427_),
    .A1(\crc16_read[11] ),
    .A2(net2191));
 sg13g2_a21oi_1 _14671_ (.A1(_01943_),
    .A2(net2191),
    .Y(_00906_),
    .B1(_06427_));
 sg13g2_o21ai_1 _14672_ (.B1(net2652),
    .Y(_06428_),
    .A1(\crc16_read[12] ),
    .A2(net2192));
 sg13g2_a21oi_1 _14673_ (.A1(_01942_),
    .A2(net2192),
    .Y(_00907_),
    .B1(_06428_));
 sg13g2_o21ai_1 _14674_ (.B1(net2647),
    .Y(_06429_),
    .A1(net4653),
    .A2(net2202));
 sg13g2_a21oi_1 _14675_ (.A1(_01941_),
    .A2(net2202),
    .Y(_00908_),
    .B1(_06429_));
 sg13g2_o21ai_1 _14676_ (.B1(net2646),
    .Y(_06430_),
    .A1(\crc16_read[14] ),
    .A2(net2191));
 sg13g2_a21oi_1 _14677_ (.A1(_01940_),
    .A2(net2191),
    .Y(_00909_),
    .B1(_06430_));
 sg13g2_o21ai_1 _14678_ (.B1(net2646),
    .Y(_06431_),
    .A1(\crc16_read[15] ),
    .A2(net2191));
 sg13g2_a21oi_1 _14679_ (.A1(_01939_),
    .A2(net2191),
    .Y(_00910_),
    .B1(_06431_));
 sg13g2_o21ai_1 _14680_ (.B1(net2663),
    .Y(_06432_),
    .A1(\i_seal.sealed_mono[0] ),
    .A2(net2212));
 sg13g2_a21oi_1 _14681_ (.A1(_01920_),
    .A2(net2212),
    .Y(_00911_),
    .B1(_06432_));
 sg13g2_o21ai_1 _14682_ (.B1(net2664),
    .Y(_06433_),
    .A1(\i_seal.sealed_mono[1] ),
    .A2(net2212));
 sg13g2_a21oi_1 _14683_ (.A1(_01918_),
    .A2(net2212),
    .Y(_00912_),
    .B1(_06433_));
 sg13g2_o21ai_1 _14684_ (.B1(net2663),
    .Y(_06434_),
    .A1(\i_seal.sealed_mono[2] ),
    .A2(net2212));
 sg13g2_a21oi_1 _14685_ (.A1(_01916_),
    .A2(net2212),
    .Y(_00913_),
    .B1(_06434_));
 sg13g2_o21ai_1 _14686_ (.B1(net2648),
    .Y(_06435_),
    .A1(\i_seal.sealed_mono[3] ),
    .A2(net2199));
 sg13g2_a21oi_1 _14687_ (.A1(_01914_),
    .A2(net2199),
    .Y(_00914_),
    .B1(_06435_));
 sg13g2_o21ai_1 _14688_ (.B1(net2668),
    .Y(_06436_),
    .A1(\i_seal.sealed_mono[4] ),
    .A2(net2216));
 sg13g2_a21oi_1 _14689_ (.A1(_01912_),
    .A2(net2217),
    .Y(_00915_),
    .B1(_06436_));
 sg13g2_o21ai_1 _14690_ (.B1(net2667),
    .Y(_06437_),
    .A1(net4160),
    .A2(net2216));
 sg13g2_a21oi_1 _14691_ (.A1(_01910_),
    .A2(net2216),
    .Y(_00916_),
    .B1(_06437_));
 sg13g2_o21ai_1 _14692_ (.B1(net2665),
    .Y(_06438_),
    .A1(\i_seal.sealed_mono[6] ),
    .A2(net2214));
 sg13g2_a21oi_1 _14693_ (.A1(_01908_),
    .A2(net2214),
    .Y(_00917_),
    .B1(_06438_));
 sg13g2_o21ai_1 _14694_ (.B1(net2667),
    .Y(_06439_),
    .A1(\i_seal.sealed_mono[7] ),
    .A2(net2214));
 sg13g2_a21oi_1 _14695_ (.A1(_01906_),
    .A2(net2214),
    .Y(_00918_),
    .B1(_06439_));
 sg13g2_o21ai_1 _14696_ (.B1(net2666),
    .Y(_06440_),
    .A1(net4489),
    .A2(net2214));
 sg13g2_a21oi_1 _14697_ (.A1(_01904_),
    .A2(net2214),
    .Y(_00919_),
    .B1(_06440_));
 sg13g2_o21ai_1 _14698_ (.B1(net2648),
    .Y(_06441_),
    .A1(net4638),
    .A2(net2199));
 sg13g2_a21oi_1 _14699_ (.A1(_01902_),
    .A2(net2201),
    .Y(_00920_),
    .B1(_06441_));
 sg13g2_o21ai_1 _14700_ (.B1(net2661),
    .Y(_06442_),
    .A1(\i_seal.sealed_mono[10] ),
    .A2(net2211));
 sg13g2_a21oi_1 _14701_ (.A1(_01900_),
    .A2(net2211),
    .Y(_00921_),
    .B1(_06442_));
 sg13g2_o21ai_1 _14702_ (.B1(net2667),
    .Y(_06443_),
    .A1(\i_seal.cur_mono[11] ),
    .A2(net2193));
 sg13g2_a21oi_1 _14703_ (.A1(_01936_),
    .A2(net2194),
    .Y(_00922_),
    .B1(_06443_));
 sg13g2_o21ai_1 _14704_ (.B1(net2648),
    .Y(_06444_),
    .A1(\i_seal.cur_mono[12] ),
    .A2(net2193));
 sg13g2_a21oi_1 _14705_ (.A1(_01935_),
    .A2(net2193),
    .Y(_00923_),
    .B1(_06444_));
 sg13g2_o21ai_1 _14706_ (.B1(net2667),
    .Y(_06445_),
    .A1(net4429),
    .A2(net2216));
 sg13g2_a21oi_1 _14707_ (.A1(_01896_),
    .A2(net2216),
    .Y(_00924_),
    .B1(_06445_));
 sg13g2_o21ai_1 _14708_ (.B1(net2660),
    .Y(_06446_),
    .A1(\i_seal.sealed_mono[14] ),
    .A2(net2213));
 sg13g2_a21oi_1 _14709_ (.A1(_01894_),
    .A2(net2211),
    .Y(_00925_),
    .B1(_06446_));
 sg13g2_o21ai_1 _14710_ (.B1(net2660),
    .Y(_06447_),
    .A1(\i_seal.cur_mono[15] ),
    .A2(net2193));
 sg13g2_a21oi_1 _14711_ (.A1(_01932_),
    .A2(net2193),
    .Y(_00926_),
    .B1(_06447_));
 sg13g2_o21ai_1 _14712_ (.B1(net2646),
    .Y(_06448_),
    .A1(net4655),
    .A2(net2200));
 sg13g2_a21oi_1 _14713_ (.A1(_01891_),
    .A2(net2200),
    .Y(_00927_),
    .B1(_06448_));
 sg13g2_o21ai_1 _14714_ (.B1(net2665),
    .Y(_06449_),
    .A1(\i_seal.sealed_mono[17] ),
    .A2(net2215));
 sg13g2_a21oi_1 _14715_ (.A1(_01889_),
    .A2(net2215),
    .Y(_00928_),
    .B1(_06449_));
 sg13g2_o21ai_1 _14716_ (.B1(net2660),
    .Y(_06450_),
    .A1(net4326),
    .A2(net2211));
 sg13g2_a21oi_1 _14717_ (.A1(_01887_),
    .A2(net2215),
    .Y(_00929_),
    .B1(_06450_));
 sg13g2_o21ai_1 _14718_ (.B1(net2660),
    .Y(_06451_),
    .A1(net4561),
    .A2(net2211));
 sg13g2_a21oi_1 _14719_ (.A1(_01885_),
    .A2(net2211),
    .Y(_00930_),
    .B1(_06451_));
 sg13g2_o21ai_1 _14720_ (.B1(net2665),
    .Y(_06452_),
    .A1(\i_seal.sealed_mono[20] ),
    .A2(net2209));
 sg13g2_a21oi_1 _14721_ (.A1(_01883_),
    .A2(net2209),
    .Y(_00931_),
    .B1(_06452_));
 sg13g2_o21ai_1 _14722_ (.B1(net2661),
    .Y(_06453_),
    .A1(\i_seal.sealed_mono[21] ),
    .A2(net2211));
 sg13g2_a21oi_1 _14723_ (.A1(_01881_),
    .A2(net2211),
    .Y(_00932_),
    .B1(_06453_));
 sg13g2_o21ai_1 _14724_ (.B1(net2651),
    .Y(_06454_),
    .A1(\i_seal.sealed_mono[22] ),
    .A2(net2209));
 sg13g2_a21oi_1 _14725_ (.A1(_01879_),
    .A2(net2209),
    .Y(_00933_),
    .B1(_06454_));
 sg13g2_o21ai_1 _14726_ (.B1(net2661),
    .Y(_06455_),
    .A1(\i_seal.sealed_mono[23] ),
    .A2(net2204));
 sg13g2_a21oi_1 _14727_ (.A1(_01877_),
    .A2(net2204),
    .Y(_00934_),
    .B1(_06455_));
 sg13g2_o21ai_1 _14728_ (.B1(net2657),
    .Y(_06456_),
    .A1(\i_seal.sealed_mono[24] ),
    .A2(net2207));
 sg13g2_a21oi_1 _14729_ (.A1(_01875_),
    .A2(net2207),
    .Y(_00935_),
    .B1(_06456_));
 sg13g2_o21ai_1 _14730_ (.B1(net2657),
    .Y(_06457_),
    .A1(\i_seal.sealed_mono[25] ),
    .A2(net2207));
 sg13g2_a21oi_1 _14731_ (.A1(_01873_),
    .A2(net2207),
    .Y(_00936_),
    .B1(_06457_));
 sg13g2_o21ai_1 _14732_ (.B1(net2657),
    .Y(_06458_),
    .A1(\i_seal.sealed_mono[26] ),
    .A2(net2208));
 sg13g2_a21oi_1 _14733_ (.A1(_01871_),
    .A2(net2208),
    .Y(_00937_),
    .B1(_06458_));
 sg13g2_o21ai_1 _14734_ (.B1(net2658),
    .Y(_06459_),
    .A1(\i_seal.sealed_mono[27] ),
    .A2(net2206));
 sg13g2_a21oi_1 _14735_ (.A1(_01869_),
    .A2(net2206),
    .Y(_00938_),
    .B1(_06459_));
 sg13g2_o21ai_1 _14736_ (.B1(net2657),
    .Y(_06460_),
    .A1(\i_seal.sealed_mono[28] ),
    .A2(net2207));
 sg13g2_a21oi_1 _14737_ (.A1(_01867_),
    .A2(net2207),
    .Y(_00939_),
    .B1(_06460_));
 sg13g2_o21ai_1 _14738_ (.B1(net2656),
    .Y(_06461_),
    .A1(net4384),
    .A2(net2207));
 sg13g2_a21oi_1 _14739_ (.A1(_01865_),
    .A2(net2207),
    .Y(_00940_),
    .B1(_06461_));
 sg13g2_o21ai_1 _14740_ (.B1(net2658),
    .Y(_06462_),
    .A1(net4403),
    .A2(net2206));
 sg13g2_a21oi_1 _14741_ (.A1(_01863_),
    .A2(net2209),
    .Y(_00941_),
    .B1(_06462_));
 sg13g2_o21ai_1 _14742_ (.B1(net2658),
    .Y(_06463_),
    .A1(net4314),
    .A2(net2205));
 sg13g2_a21oi_1 _14743_ (.A1(_01861_),
    .A2(net2205),
    .Y(_00942_),
    .B1(_06463_));
 sg13g2_o21ai_1 _14744_ (.B1(net2648),
    .Y(_06464_),
    .A1(net4541),
    .A2(net2201));
 sg13g2_a21oi_1 _14745_ (.A1(_01858_),
    .A2(net2201),
    .Y(_00943_),
    .B1(_06464_));
 sg13g2_o21ai_1 _14746_ (.B1(net2664),
    .Y(_06465_),
    .A1(\i_seal.sealed_value[1] ),
    .A2(net2212));
 sg13g2_a21oi_1 _14747_ (.A1(_01857_),
    .A2(net2213),
    .Y(_00944_),
    .B1(_06465_));
 sg13g2_o21ai_1 _14748_ (.B1(net2663),
    .Y(_06466_),
    .A1(\i_seal.sealed_value[2] ),
    .A2(net2212));
 sg13g2_a21oi_1 _14749_ (.A1(_01856_),
    .A2(net2213),
    .Y(_00945_),
    .B1(_06466_));
 sg13g2_o21ai_1 _14750_ (.B1(net2644),
    .Y(_06467_),
    .A1(\i_seal.sealed_value[3] ),
    .A2(net2199));
 sg13g2_a21oi_1 _14751_ (.A1(_01855_),
    .A2(net2199),
    .Y(_00946_),
    .B1(_06467_));
 sg13g2_o21ai_1 _14752_ (.B1(net2667),
    .Y(_06468_),
    .A1(\i_seal.sealed_value[4] ),
    .A2(net2217));
 sg13g2_a21oi_1 _14753_ (.A1(_01854_),
    .A2(net2217),
    .Y(_00947_),
    .B1(_06468_));
 sg13g2_o21ai_1 _14754_ (.B1(net2668),
    .Y(_06469_),
    .A1(net4443),
    .A2(net2216));
 sg13g2_a21oi_1 _14755_ (.A1(_01853_),
    .A2(net2216),
    .Y(_00948_),
    .B1(_06469_));
 sg13g2_o21ai_1 _14756_ (.B1(net2666),
    .Y(_06470_),
    .A1(\i_seal.sealed_value[6] ),
    .A2(net2215));
 sg13g2_a21oi_1 _14757_ (.A1(_01852_),
    .A2(net2215),
    .Y(_00949_),
    .B1(_06470_));
 sg13g2_o21ai_1 _14758_ (.B1(net2667),
    .Y(_06471_),
    .A1(\i_seal.sealed_value[7] ),
    .A2(net2215));
 sg13g2_a21oi_1 _14759_ (.A1(_01851_),
    .A2(net2214),
    .Y(_00950_),
    .B1(_06471_));
 sg13g2_o21ai_1 _14760_ (.B1(net2665),
    .Y(_06472_),
    .A1(\i_seal.sealed_value[8] ),
    .A2(net2214));
 sg13g2_a21oi_1 _14761_ (.A1(_01850_),
    .A2(net2215),
    .Y(_00951_),
    .B1(_06472_));
 sg13g2_o21ai_1 _14762_ (.B1(net2643),
    .Y(_06473_),
    .A1(\i_seal.sealed_value[9] ),
    .A2(net2195));
 sg13g2_a21oi_1 _14763_ (.A1(_01849_),
    .A2(net2195),
    .Y(_00952_),
    .B1(_06473_));
 sg13g2_o21ai_1 _14764_ (.B1(net2646),
    .Y(_06474_),
    .A1(\i_seal.sealed_value[10] ),
    .A2(net2200));
 sg13g2_a21oi_1 _14765_ (.A1(_01848_),
    .A2(net2200),
    .Y(_00953_),
    .B1(_06474_));
 sg13g2_o21ai_1 _14766_ (.B1(net2645),
    .Y(_06475_),
    .A1(\i_seal.sealed_value[11] ),
    .A2(net2197));
 sg13g2_a21oi_1 _14767_ (.A1(_01847_),
    .A2(net2197),
    .Y(_00954_),
    .B1(_06475_));
 sg13g2_o21ai_1 _14768_ (.B1(net2645),
    .Y(_06476_),
    .A1(net4596),
    .A2(net2197));
 sg13g2_a21oi_1 _14769_ (.A1(_01846_),
    .A2(net2198),
    .Y(_00955_),
    .B1(_06476_));
 sg13g2_o21ai_1 _14770_ (.B1(net2645),
    .Y(_06477_),
    .A1(\i_seal.sealed_value[13] ),
    .A2(net2199));
 sg13g2_a21oi_1 _14771_ (.A1(_01845_),
    .A2(net2197),
    .Y(_00956_),
    .B1(_06477_));
 sg13g2_o21ai_1 _14772_ (.B1(net2646),
    .Y(_06478_),
    .A1(\i_seal.sealed_value[14] ),
    .A2(net2200));
 sg13g2_a21oi_1 _14773_ (.A1(_01844_),
    .A2(net2200),
    .Y(_00957_),
    .B1(_06478_));
 sg13g2_o21ai_1 _14774_ (.B1(net2643),
    .Y(_06479_),
    .A1(\i_seal.sealed_value[15] ),
    .A2(net2196));
 sg13g2_a21oi_1 _14775_ (.A1(_01843_),
    .A2(net2196),
    .Y(_00958_),
    .B1(_06479_));
 sg13g2_o21ai_1 _14776_ (.B1(net2647),
    .Y(_06480_),
    .A1(\i_seal.sealed_value[16] ),
    .A2(net2200));
 sg13g2_a21oi_1 _14777_ (.A1(_01841_),
    .A2(net2200),
    .Y(_00959_),
    .B1(_06480_));
 sg13g2_o21ai_1 _14778_ (.B1(net2660),
    .Y(_06481_),
    .A1(\i_seal.sealed_value[17] ),
    .A2(net2210));
 sg13g2_a21oi_1 _14779_ (.A1(_01839_),
    .A2(net2210),
    .Y(_00960_),
    .B1(_06481_));
 sg13g2_o21ai_1 _14780_ (.B1(net2660),
    .Y(_06482_),
    .A1(\i_seal.sealed_value[18] ),
    .A2(net2204));
 sg13g2_a21oi_1 _14781_ (.A1(_01837_),
    .A2(net2210),
    .Y(_00961_),
    .B1(_06482_));
 sg13g2_o21ai_1 _14782_ (.B1(net2653),
    .Y(_06483_),
    .A1(\i_seal.sealed_value[19] ),
    .A2(net2203));
 sg13g2_a21oi_1 _14783_ (.A1(_01835_),
    .A2(net2203),
    .Y(_00962_),
    .B1(_06483_));
 sg13g2_o21ai_1 _14784_ (.B1(net2665),
    .Y(_06484_),
    .A1(\i_seal.sealed_value[20] ),
    .A2(net2209));
 sg13g2_a21oi_1 _14785_ (.A1(_01833_),
    .A2(net2209),
    .Y(_00963_),
    .B1(_06484_));
 sg13g2_o21ai_1 _14786_ (.B1(net2642),
    .Y(_06485_),
    .A1(\i_seal.sealed_value[21] ),
    .A2(net2203));
 sg13g2_a21oi_1 _14787_ (.A1(_01831_),
    .A2(net2203),
    .Y(_00964_),
    .B1(_06485_));
 sg13g2_o21ai_1 _14788_ (.B1(net2651),
    .Y(_06486_),
    .A1(\i_seal.sealed_value[22] ),
    .A2(net2204));
 sg13g2_a21oi_1 _14789_ (.A1(_01829_),
    .A2(net2204),
    .Y(_00965_),
    .B1(_06486_));
 sg13g2_o21ai_1 _14790_ (.B1(net2642),
    .Y(_06487_),
    .A1(\i_seal.sealed_value[23] ),
    .A2(net2202));
 sg13g2_a21oi_1 _14791_ (.A1(_01827_),
    .A2(net2202),
    .Y(_00966_),
    .B1(_06487_));
 sg13g2_o21ai_1 _14792_ (.B1(net2651),
    .Y(_06488_),
    .A1(\i_seal.sealed_value[24] ),
    .A2(net2203));
 sg13g2_a21oi_1 _14793_ (.A1(_01825_),
    .A2(net2203),
    .Y(_00967_),
    .B1(_06488_));
 sg13g2_o21ai_1 _14794_ (.B1(net2651),
    .Y(_06489_),
    .A1(\i_seal.sealed_value[25] ),
    .A2(net2204));
 sg13g2_a21oi_1 _14795_ (.A1(_01823_),
    .A2(net2204),
    .Y(_00968_),
    .B1(_06489_));
 sg13g2_o21ai_1 _14796_ (.B1(net2655),
    .Y(_06490_),
    .A1(\i_seal.sealed_value[26] ),
    .A2(net2205));
 sg13g2_a21oi_1 _14797_ (.A1(_01821_),
    .A2(net2206),
    .Y(_00969_),
    .B1(_06490_));
 sg13g2_o21ai_1 _14798_ (.B1(net2655),
    .Y(_06491_),
    .A1(\i_seal.sealed_value[27] ),
    .A2(net2205));
 sg13g2_a21oi_1 _14799_ (.A1(_01819_),
    .A2(net2205),
    .Y(_00970_),
    .B1(_06491_));
 sg13g2_o21ai_1 _14800_ (.B1(net2651),
    .Y(_06492_),
    .A1(\i_seal.sealed_value[28] ),
    .A2(net2205));
 sg13g2_a21oi_1 _14801_ (.A1(_01817_),
    .A2(net2205),
    .Y(_00971_),
    .B1(_06492_));
 sg13g2_o21ai_1 _14802_ (.B1(net2653),
    .Y(_06493_),
    .A1(\i_seal.sealed_value[29] ),
    .A2(net2203));
 sg13g2_a21oi_1 _14803_ (.A1(_01815_),
    .A2(net2203),
    .Y(_00972_),
    .B1(_06493_));
 sg13g2_o21ai_1 _14804_ (.B1(net2651),
    .Y(_06494_),
    .A1(\i_seal.sealed_value[30] ),
    .A2(net2206));
 sg13g2_a21oi_1 _14805_ (.A1(_01813_),
    .A2(net2208),
    .Y(_00973_),
    .B1(_06494_));
 sg13g2_o21ai_1 _14806_ (.B1(net2656),
    .Y(_06495_),
    .A1(\i_seal.sealed_value[31] ),
    .A2(net2206));
 sg13g2_a21oi_1 _14807_ (.A1(_01811_),
    .A2(net2205),
    .Y(_00974_),
    .B1(_06495_));
 sg13g2_o21ai_1 _14808_ (.B1(net2658),
    .Y(_06496_),
    .A1(net4538),
    .A2(net2206));
 sg13g2_inv_1 _14809_ (.Y(_00975_),
    .A(_06496_));
 sg13g2_nor2_1 _14810_ (.A(\i_seal.session_locked ),
    .B(net2192),
    .Y(_06497_));
 sg13g2_o21ai_1 _14811_ (.B1(net2657),
    .Y(_06498_),
    .A1(net4084),
    .A2(net2158));
 sg13g2_a21oi_1 _14812_ (.A1(_01929_),
    .A2(net2158),
    .Y(_00976_),
    .B1(net4085));
 sg13g2_o21ai_1 _14813_ (.B1(net2657),
    .Y(_06499_),
    .A1(\i_seal.sealed_sid[1] ),
    .A2(net2158));
 sg13g2_a21oi_1 _14814_ (.A1(_01928_),
    .A2(net2158),
    .Y(_00977_),
    .B1(_06499_));
 sg13g2_o21ai_1 _14815_ (.B1(net2656),
    .Y(_06500_),
    .A1(\i_seal.sealed_sid[2] ),
    .A2(net2157));
 sg13g2_a21oi_1 _14816_ (.A1(_01927_),
    .A2(net2157),
    .Y(_00978_),
    .B1(_06500_));
 sg13g2_o21ai_1 _14817_ (.B1(net2655),
    .Y(_06501_),
    .A1(\i_seal.sealed_sid[3] ),
    .A2(net2156));
 sg13g2_a21oi_1 _14818_ (.A1(_01926_),
    .A2(net2156),
    .Y(_00979_),
    .B1(_06501_));
 sg13g2_o21ai_1 _14819_ (.B1(net2656),
    .Y(_06502_),
    .A1(net4020),
    .A2(net2157));
 sg13g2_a21oi_1 _14820_ (.A1(_01925_),
    .A2(net2157),
    .Y(_00980_),
    .B1(_06502_));
 sg13g2_o21ai_1 _14821_ (.B1(net2655),
    .Y(_06503_),
    .A1(\i_seal.sealed_sid[5] ),
    .A2(net2156));
 sg13g2_a21oi_1 _14822_ (.A1(_01924_),
    .A2(net2156),
    .Y(_00981_),
    .B1(_06503_));
 sg13g2_o21ai_1 _14823_ (.B1(net2655),
    .Y(_06504_),
    .A1(\i_seal.sealed_sid[6] ),
    .A2(net2156));
 sg13g2_a21oi_1 _14824_ (.A1(_01923_),
    .A2(net2156),
    .Y(_00982_),
    .B1(_06504_));
 sg13g2_o21ai_1 _14825_ (.B1(net2655),
    .Y(_06505_),
    .A1(net3992),
    .A2(net2156));
 sg13g2_a21oi_1 _14826_ (.A1(_01922_),
    .A2(net2156),
    .Y(_00983_),
    .B1(net3993));
 sg13g2_o21ai_1 _14827_ (.B1(net2662),
    .Y(_06506_),
    .A1(_01921_),
    .A2(net2193));
 sg13g2_a21oi_1 _14828_ (.A1(_01921_),
    .A2(net2193),
    .Y(_00984_),
    .B1(_06506_));
 sg13g2_o21ai_1 _14829_ (.B1(_01919_),
    .Y(_06507_),
    .A1(_01921_),
    .A2(net2193));
 sg13g2_nand3_1 _14830_ (.B(net4202),
    .C(net2216),
    .A(net4120),
    .Y(_06508_));
 sg13g2_and3_1 _14831_ (.X(_00985_),
    .A(net2662),
    .B(_06507_),
    .C(_06508_));
 sg13g2_or2_1 _14832_ (.X(_06509_),
    .B(_06508_),
    .A(_01917_));
 sg13g2_nand2_1 _14833_ (.Y(_06510_),
    .A(net2667),
    .B(_06509_));
 sg13g2_a21oi_1 _14834_ (.A1(_01917_),
    .A2(_06508_),
    .Y(_00986_),
    .B1(_06510_));
 sg13g2_and2_1 _14835_ (.A(_01915_),
    .B(_06509_),
    .X(_06511_));
 sg13g2_nor2_1 _14836_ (.A(_01915_),
    .B(_06509_),
    .Y(_06512_));
 sg13g2_nor3_1 _14837_ (.A(net2428),
    .B(_06511_),
    .C(_06512_),
    .Y(_00987_));
 sg13g2_nor3_2 _14838_ (.A(_01913_),
    .B(_01915_),
    .C(_06509_),
    .Y(_06513_));
 sg13g2_o21ai_1 _14839_ (.B1(net2668),
    .Y(_06514_),
    .A1(net4319),
    .A2(_06512_));
 sg13g2_nor2_1 _14840_ (.A(_06513_),
    .B(_06514_),
    .Y(_00988_));
 sg13g2_xnor2_1 _14841_ (.Y(_06515_),
    .A(net3889),
    .B(_06513_));
 sg13g2_nor2_1 _14842_ (.A(net2428),
    .B(_06515_),
    .Y(_00989_));
 sg13g2_a21oi_1 _14843_ (.A1(net3889),
    .A2(_06513_),
    .Y(_06516_),
    .B1(net3713));
 sg13g2_and3_2 _14844_ (.X(_06517_),
    .A(net3713),
    .B(net3889),
    .C(_06513_));
 sg13g2_nor3_1 _14845_ (.A(net2425),
    .B(net3890),
    .C(_06517_),
    .Y(_00990_));
 sg13g2_xnor2_1 _14846_ (.Y(_06518_),
    .A(net4308),
    .B(_06517_));
 sg13g2_nor2_1 _14847_ (.A(net2425),
    .B(_06518_),
    .Y(_00991_));
 sg13g2_a21oi_1 _14848_ (.A1(\i_seal.mono_count[7] ),
    .A2(_06517_),
    .Y(_06519_),
    .B1(net3931));
 sg13g2_and3_1 _14849_ (.X(_06520_),
    .A(net3931),
    .B(net4308),
    .C(_06517_));
 sg13g2_nor3_1 _14850_ (.A(net2425),
    .B(net3932),
    .C(_06520_),
    .Y(_00992_));
 sg13g2_nor2_1 _14851_ (.A(net3654),
    .B(_06520_),
    .Y(_06521_));
 sg13g2_and2_1 _14852_ (.A(net3654),
    .B(_06520_),
    .X(_06522_));
 sg13g2_nor3_1 _14853_ (.A(net2425),
    .B(_06521_),
    .C(_06522_),
    .Y(_00993_));
 sg13g2_and2_1 _14854_ (.A(net3727),
    .B(_06522_),
    .X(_06523_));
 sg13g2_o21ai_1 _14855_ (.B1(net2670),
    .Y(_06524_),
    .A1(net3727),
    .A2(_06522_));
 sg13g2_nor2_1 _14856_ (.A(_06523_),
    .B(_06524_),
    .Y(_00994_));
 sg13g2_xnor2_1 _14857_ (.Y(_06525_),
    .A(net4273),
    .B(_06523_));
 sg13g2_nor2_1 _14858_ (.A(net2425),
    .B(_06525_),
    .Y(_00995_));
 sg13g2_a21oi_1 _14859_ (.A1(\i_seal.mono_count[11] ),
    .A2(_06523_),
    .Y(_06526_),
    .B1(net3895));
 sg13g2_and3_2 _14860_ (.X(_06527_),
    .A(net3895),
    .B(net4273),
    .C(_06523_));
 sg13g2_nor3_1 _14861_ (.A(net2425),
    .B(net3896),
    .C(_06527_),
    .Y(_00996_));
 sg13g2_xnor2_1 _14862_ (.Y(_06528_),
    .A(net3901),
    .B(_06527_));
 sg13g2_nor2_1 _14863_ (.A(net2426),
    .B(_06528_),
    .Y(_00997_));
 sg13g2_a21oi_1 _14864_ (.A1(net3901),
    .A2(_06527_),
    .Y(_06529_),
    .B1(net3864));
 sg13g2_and3_1 _14865_ (.X(_06530_),
    .A(net3864),
    .B(net3901),
    .C(_06527_));
 sg13g2_nor3_1 _14866_ (.A(net2426),
    .B(net3902),
    .C(_06530_),
    .Y(_00998_));
 sg13g2_nor2_1 _14867_ (.A(net3870),
    .B(_06530_),
    .Y(_06531_));
 sg13g2_and2_1 _14868_ (.A(net3870),
    .B(_06530_),
    .X(_06532_));
 sg13g2_nor3_1 _14869_ (.A(net2426),
    .B(_06531_),
    .C(_06532_),
    .Y(_00999_));
 sg13g2_and2_1 _14870_ (.A(net3892),
    .B(_06532_),
    .X(_06533_));
 sg13g2_o21ai_1 _14871_ (.B1(net2670),
    .Y(_06534_),
    .A1(net3892),
    .A2(_06532_));
 sg13g2_nor2_1 _14872_ (.A(_06533_),
    .B(_06534_),
    .Y(_01000_));
 sg13g2_xnor2_1 _14873_ (.Y(_06535_),
    .A(net4039),
    .B(_06533_));
 sg13g2_nor2_1 _14874_ (.A(net2427),
    .B(_06535_),
    .Y(_01001_));
 sg13g2_a21oi_1 _14875_ (.A1(\i_seal.mono_count[17] ),
    .A2(_06533_),
    .Y(_06536_),
    .B1(net3971));
 sg13g2_and3_2 _14876_ (.X(_06537_),
    .A(net3971),
    .B(net4039),
    .C(_06533_));
 sg13g2_nor3_1 _14877_ (.A(net2427),
    .B(net3972),
    .C(_06537_),
    .Y(_01002_));
 sg13g2_xnor2_1 _14878_ (.Y(_06538_),
    .A(net3758),
    .B(_06537_));
 sg13g2_nor2_1 _14879_ (.A(net2427),
    .B(_06538_),
    .Y(_01003_));
 sg13g2_a21oi_1 _14880_ (.A1(net3758),
    .A2(_06537_),
    .Y(_06539_),
    .B1(net3665));
 sg13g2_and3_1 _14881_ (.X(_06540_),
    .A(net3665),
    .B(net3758),
    .C(_06537_));
 sg13g2_nor3_1 _14882_ (.A(net2427),
    .B(net3759),
    .C(_06540_),
    .Y(_01004_));
 sg13g2_nor2_1 _14883_ (.A(net3835),
    .B(_06540_),
    .Y(_06541_));
 sg13g2_and2_1 _14884_ (.A(net3835),
    .B(_06540_),
    .X(_06542_));
 sg13g2_nor3_1 _14885_ (.A(net2427),
    .B(_06541_),
    .C(_06542_),
    .Y(_01005_));
 sg13g2_xnor2_1 _14886_ (.Y(_06543_),
    .A(net4031),
    .B(_06542_));
 sg13g2_nor2_1 _14887_ (.A(net2427),
    .B(_06543_),
    .Y(_01006_));
 sg13g2_a21oi_1 _14888_ (.A1(net4031),
    .A2(_06542_),
    .Y(_06544_),
    .B1(net3999));
 sg13g2_and3_1 _14889_ (.X(_06545_),
    .A(net3999),
    .B(net4031),
    .C(_06542_));
 sg13g2_nor3_1 _14890_ (.A(net2428),
    .B(_06544_),
    .C(_06545_),
    .Y(_01007_));
 sg13g2_and2_1 _14891_ (.A(net3673),
    .B(_06545_),
    .X(_06546_));
 sg13g2_o21ai_1 _14892_ (.B1(net2666),
    .Y(_06547_),
    .A1(net3673),
    .A2(_06545_));
 sg13g2_nor2_1 _14893_ (.A(_06546_),
    .B(_06547_),
    .Y(_01008_));
 sg13g2_nand2_1 _14894_ (.Y(_06548_),
    .A(net3979),
    .B(_06546_));
 sg13g2_o21ai_1 _14895_ (.B1(net2666),
    .Y(_06549_),
    .A1(net3979),
    .A2(_06546_));
 sg13g2_nor2b_1 _14896_ (.A(_06549_),
    .B_N(_06548_),
    .Y(_01009_));
 sg13g2_a21oi_1 _14897_ (.A1(\i_seal.mono_count[25] ),
    .A2(_06546_),
    .Y(_06550_),
    .B1(net3550));
 sg13g2_nor2_1 _14898_ (.A(_01872_),
    .B(_06548_),
    .Y(_06551_));
 sg13g2_nor3_1 _14899_ (.A(net2428),
    .B(net3551),
    .C(_06551_),
    .Y(_01010_));
 sg13g2_nor3_1 _14900_ (.A(_01870_),
    .B(_01872_),
    .C(_06548_),
    .Y(_06552_));
 sg13g2_o21ai_1 _14901_ (.B1(net2657),
    .Y(_06553_),
    .A1(net3917),
    .A2(_06551_));
 sg13g2_nor2_1 _14902_ (.A(_06552_),
    .B(_06553_),
    .Y(_01011_));
 sg13g2_and2_1 _14903_ (.A(net3919),
    .B(_06552_),
    .X(_06554_));
 sg13g2_o21ai_1 _14904_ (.B1(net2657),
    .Y(_06555_),
    .A1(net3919),
    .A2(_06552_));
 sg13g2_nor2_1 _14905_ (.A(_06554_),
    .B(_06555_),
    .Y(_01012_));
 sg13g2_o21ai_1 _14906_ (.B1(net2673),
    .Y(_06556_),
    .A1(net3539),
    .A2(_06554_));
 sg13g2_a21oi_1 _14907_ (.A1(net3539),
    .A2(_06554_),
    .Y(_01013_),
    .B1(_06556_));
 sg13g2_a21oi_1 _14908_ (.A1(net3539),
    .A2(_06554_),
    .Y(_06557_),
    .B1(net3685));
 sg13g2_nand3_1 _14909_ (.B(net3539),
    .C(_06554_),
    .A(net3685),
    .Y(_06558_));
 sg13g2_nand2_1 _14910_ (.Y(_06559_),
    .A(net2673),
    .B(_06558_));
 sg13g2_nor2_1 _14911_ (.A(net3686),
    .B(_06559_),
    .Y(_01014_));
 sg13g2_o21ai_1 _14912_ (.B1(net2673),
    .Y(_06560_),
    .A1(_01862_),
    .A2(_06558_));
 sg13g2_a21oi_1 _14913_ (.A1(_01862_),
    .A2(_06558_),
    .Y(_01015_),
    .B1(_06560_));
 sg13g2_o21ai_1 _14914_ (.B1(net2663),
    .Y(_06561_),
    .A1(net4187),
    .A2(net1944));
 sg13g2_a21oi_1 _14915_ (.A1(_01921_),
    .A2(net1944),
    .Y(_01016_),
    .B1(_06561_));
 sg13g2_o21ai_1 _14916_ (.B1(net2662),
    .Y(_06562_),
    .A1(net4110),
    .A2(net1944));
 sg13g2_a21oi_1 _14917_ (.A1(_01919_),
    .A2(net1944),
    .Y(_01017_),
    .B1(_06562_));
 sg13g2_o21ai_1 _14918_ (.B1(net2662),
    .Y(_06563_),
    .A1(net4079),
    .A2(net1944));
 sg13g2_a21oi_1 _14919_ (.A1(_01917_),
    .A2(net1944),
    .Y(_01018_),
    .B1(_06563_));
 sg13g2_o21ai_1 _14920_ (.B1(net2667),
    .Y(_06564_),
    .A1(\i_seal.cur_mono[3] ),
    .A2(net1943));
 sg13g2_a21oi_1 _14921_ (.A1(_01915_),
    .A2(net1938),
    .Y(_01019_),
    .B1(_06564_));
 sg13g2_o21ai_1 _14922_ (.B1(net2668),
    .Y(_06565_),
    .A1(net4114),
    .A2(net1943));
 sg13g2_a21oi_1 _14923_ (.A1(_01913_),
    .A2(net1938),
    .Y(_01020_),
    .B1(_06565_));
 sg13g2_o21ai_1 _14924_ (.B1(net2668),
    .Y(_06566_),
    .A1(net4067),
    .A2(net1938));
 sg13g2_a21oi_1 _14925_ (.A1(_01911_),
    .A2(net1938),
    .Y(_01021_),
    .B1(_06566_));
 sg13g2_o21ai_1 _14926_ (.B1(net2668),
    .Y(_06567_),
    .A1(\i_seal.cur_mono[6] ),
    .A2(net1938));
 sg13g2_a21oi_1 _14927_ (.A1(_01909_),
    .A2(net1938),
    .Y(_01022_),
    .B1(_06567_));
 sg13g2_o21ai_1 _14928_ (.B1(net2668),
    .Y(_06568_),
    .A1(net4253),
    .A2(net1938));
 sg13g2_a21oi_1 _14929_ (.A1(_01907_),
    .A2(net1938),
    .Y(_01023_),
    .B1(_06568_));
 sg13g2_o21ai_1 _14930_ (.B1(net2670),
    .Y(_06569_),
    .A1(net3986),
    .A2(net1939));
 sg13g2_a21oi_1 _14931_ (.A1(_01905_),
    .A2(net1939),
    .Y(_01024_),
    .B1(_06569_));
 sg13g2_o21ai_1 _14932_ (.B1(net2670),
    .Y(_06570_),
    .A1(\i_seal.cur_mono[9] ),
    .A2(net1941));
 sg13g2_a21oi_1 _14933_ (.A1(_01903_),
    .A2(net1941),
    .Y(_01025_),
    .B1(_06570_));
 sg13g2_o21ai_1 _14934_ (.B1(net2670),
    .Y(_06571_),
    .A1(\i_seal.cur_mono[10] ),
    .A2(net1939));
 sg13g2_a21oi_1 _14935_ (.A1(_01901_),
    .A2(net1941),
    .Y(_01026_),
    .B1(_06571_));
 sg13g2_o21ai_1 _14936_ (.B1(net2671),
    .Y(_06572_),
    .A1(net4371),
    .A2(net1941));
 sg13g2_a21oi_1 _14937_ (.A1(_01899_),
    .A2(net1941),
    .Y(_01027_),
    .B1(_06572_));
 sg13g2_o21ai_1 _14938_ (.B1(net2671),
    .Y(_06573_),
    .A1(net4349),
    .A2(net1942));
 sg13g2_a21oi_1 _14939_ (.A1(_01898_),
    .A2(net1941),
    .Y(_01028_),
    .B1(_06573_));
 sg13g2_o21ai_1 _14940_ (.B1(net2670),
    .Y(_06574_),
    .A1(net4181),
    .A2(net1941));
 sg13g2_a21oi_1 _14941_ (.A1(_01897_),
    .A2(net1941),
    .Y(_01029_),
    .B1(_06574_));
 sg13g2_o21ai_1 _14942_ (.B1(net2670),
    .Y(_06575_),
    .A1(\i_seal.cur_mono[14] ),
    .A2(net1940));
 sg13g2_a21oi_1 _14943_ (.A1(_01895_),
    .A2(net1940),
    .Y(_01030_),
    .B1(_06575_));
 sg13g2_o21ai_1 _14944_ (.B1(net2670),
    .Y(_06576_),
    .A1(\i_seal.cur_mono[15] ),
    .A2(net1939));
 sg13g2_a21oi_1 _14945_ (.A1(_01893_),
    .A2(net1940),
    .Y(_01031_),
    .B1(_06576_));
 sg13g2_o21ai_1 _14946_ (.B1(net2672),
    .Y(_06577_),
    .A1(\i_seal.cur_mono[16] ),
    .A2(net1940));
 sg13g2_a21oi_1 _14947_ (.A1(_01892_),
    .A2(net1940),
    .Y(_01032_),
    .B1(_06577_));
 sg13g2_o21ai_1 _14948_ (.B1(net2671),
    .Y(_06578_),
    .A1(\i_seal.cur_mono[17] ),
    .A2(net1937));
 sg13g2_a21oi_1 _14949_ (.A1(_01890_),
    .A2(net1940),
    .Y(_01033_),
    .B1(_06578_));
 sg13g2_o21ai_1 _14950_ (.B1(net2671),
    .Y(_06579_),
    .A1(net4015),
    .A2(net1939));
 sg13g2_a21oi_1 _14951_ (.A1(_01888_),
    .A2(net1939),
    .Y(_01034_),
    .B1(_06579_));
 sg13g2_o21ai_1 _14952_ (.B1(net2671),
    .Y(_06580_),
    .A1(net4059),
    .A2(net1939));
 sg13g2_a21oi_1 _14953_ (.A1(_01886_),
    .A2(net1939),
    .Y(_01035_),
    .B1(_06580_));
 sg13g2_o21ai_1 _14954_ (.B1(net2671),
    .Y(_06581_),
    .A1(\i_seal.cur_mono[20] ),
    .A2(net1937));
 sg13g2_a21oi_1 _14955_ (.A1(_01884_),
    .A2(net1936),
    .Y(_01036_),
    .B1(_06581_));
 sg13g2_o21ai_1 _14956_ (.B1(net2666),
    .Y(_06582_),
    .A1(\i_seal.cur_mono[21] ),
    .A2(net1935));
 sg13g2_a21oi_1 _14957_ (.A1(_01882_),
    .A2(net1935),
    .Y(_01037_),
    .B1(_06582_));
 sg13g2_o21ai_1 _14958_ (.B1(net2671),
    .Y(_06583_),
    .A1(\i_seal.cur_mono[22] ),
    .A2(net1937));
 sg13g2_a21oi_1 _14959_ (.A1(_01880_),
    .A2(net1936),
    .Y(_01038_),
    .B1(_06583_));
 sg13g2_o21ai_1 _14960_ (.B1(net2665),
    .Y(_06584_),
    .A1(\i_seal.cur_mono[23] ),
    .A2(net1935));
 sg13g2_a21oi_1 _14961_ (.A1(_01878_),
    .A2(net1934),
    .Y(_01039_),
    .B1(_06584_));
 sg13g2_o21ai_1 _14962_ (.B1(net2665),
    .Y(_06585_),
    .A1(\i_seal.cur_mono[24] ),
    .A2(net1935));
 sg13g2_a21oi_1 _14963_ (.A1(_01876_),
    .A2(net1935),
    .Y(_01040_),
    .B1(_06585_));
 sg13g2_o21ai_1 _14964_ (.B1(net2665),
    .Y(_06586_),
    .A1(net3825),
    .A2(net1935));
 sg13g2_a21oi_1 _14965_ (.A1(_01874_),
    .A2(net1934),
    .Y(_01041_),
    .B1(_06586_));
 sg13g2_o21ai_1 _14966_ (.B1(net2658),
    .Y(_06587_),
    .A1(net3982),
    .A2(net1934));
 sg13g2_a21oi_1 _14967_ (.A1(_01872_),
    .A2(net1934),
    .Y(_01042_),
    .B1(_06587_));
 sg13g2_o21ai_1 _14968_ (.B1(net2659),
    .Y(_06588_),
    .A1(\i_seal.cur_mono[27] ),
    .A2(net1934));
 sg13g2_a21oi_1 _14969_ (.A1(_01870_),
    .A2(net1934),
    .Y(_01043_),
    .B1(_06588_));
 sg13g2_o21ai_1 _14970_ (.B1(net2658),
    .Y(_06589_),
    .A1(net3844),
    .A2(net1934));
 sg13g2_a21oi_1 _14971_ (.A1(_01868_),
    .A2(net1934),
    .Y(_01044_),
    .B1(_06589_));
 sg13g2_o21ai_1 _14972_ (.B1(net2658),
    .Y(_06590_),
    .A1(net4094),
    .A2(net1936));
 sg13g2_a21oi_1 _14973_ (.A1(_01866_),
    .A2(net1936),
    .Y(_01045_),
    .B1(_06590_));
 sg13g2_o21ai_1 _14974_ (.B1(net2673),
    .Y(_06591_),
    .A1(net3846),
    .A2(net1936));
 sg13g2_a21oi_1 _14975_ (.A1(_01864_),
    .A2(net1936),
    .Y(_01046_),
    .B1(net3847));
 sg13g2_o21ai_1 _14976_ (.B1(net2673),
    .Y(_06592_),
    .A1(net4047),
    .A2(net1936));
 sg13g2_a21oi_1 _14977_ (.A1(_01862_),
    .A2(net1936),
    .Y(_01047_),
    .B1(net4048));
 sg13g2_nand2_1 _14978_ (.Y(_06593_),
    .A(net3527),
    .B(_06407_));
 sg13g2_o21ai_1 _14979_ (.B1(_06593_),
    .Y(_01048_),
    .A1(_04429_),
    .A2(net1997));
 sg13g2_nand2_1 _14980_ (.Y(_06594_),
    .A(net3675),
    .B(_06407_));
 sg13g2_o21ai_1 _14981_ (.B1(_06594_),
    .Y(_01049_),
    .A1(_04433_),
    .A2(net1997));
 sg13g2_nand2_1 _14982_ (.Y(_06595_),
    .A(net3612),
    .B(_06407_));
 sg13g2_o21ai_1 _14983_ (.B1(_06595_),
    .Y(_01050_),
    .A1(_04434_),
    .A2(net1997));
 sg13g2_nand2_1 _14984_ (.Y(_06596_),
    .A(net3645),
    .B(_06407_));
 sg13g2_o21ai_1 _14985_ (.B1(_06596_),
    .Y(_01051_),
    .A1(_04438_),
    .A2(net1997));
 sg13g2_nand2_1 _14986_ (.Y(_06597_),
    .A(net3647),
    .B(_06407_));
 sg13g2_o21ai_1 _14987_ (.B1(_06597_),
    .Y(_01052_),
    .A1(_04441_),
    .A2(net1997));
 sg13g2_nand2_1 _14988_ (.Y(_06598_),
    .A(net3616),
    .B(_06407_));
 sg13g2_o21ai_1 _14989_ (.B1(_06598_),
    .Y(_01053_),
    .A1(_04444_),
    .A2(net1998));
 sg13g2_a22oi_1 _14990_ (.Y(_01054_),
    .B1(_06408_),
    .B2(_04450_),
    .A2(net1997),
    .A1(_01860_));
 sg13g2_a22oi_1 _14991_ (.Y(_01055_),
    .B1(_06408_),
    .B2(_04454_),
    .A2(net1998),
    .A1(_01859_));
 sg13g2_nor2b_2 _14992_ (.A(net2002),
    .B_N(_05849_),
    .Y(_06599_));
 sg13g2_o21ai_1 _14993_ (.B1(net2637),
    .Y(_06600_),
    .A1(net5045),
    .A2(net1924));
 sg13g2_a21oi_1 _14994_ (.A1(_01779_),
    .A2(net1924),
    .Y(_01056_),
    .B1(_06600_));
 sg13g2_o21ai_1 _14995_ (.B1(net2644),
    .Y(_06601_),
    .A1(net4572),
    .A2(net1925));
 sg13g2_a21oi_1 _14996_ (.A1(net2452),
    .A2(net1925),
    .Y(_01057_),
    .B1(_06601_));
 sg13g2_o21ai_1 _14997_ (.B1(net2648),
    .Y(_06602_),
    .A1(net4420),
    .A2(net1932));
 sg13g2_a21oi_1 _14998_ (.A1(_01777_),
    .A2(net1931),
    .Y(_01058_),
    .B1(_06602_));
 sg13g2_o21ai_1 _14999_ (.B1(net2644),
    .Y(_06603_),
    .A1(net4479),
    .A2(net1925));
 sg13g2_a21oi_1 _15000_ (.A1(net2453),
    .A2(net1924),
    .Y(_01059_),
    .B1(_06603_));
 sg13g2_o21ai_1 _15001_ (.B1(net2662),
    .Y(_06604_),
    .A1(net3956),
    .A2(net1933));
 sg13g2_a21oi_1 _15002_ (.A1(_01775_),
    .A2(net1932),
    .Y(_01060_),
    .B1(_06604_));
 sg13g2_o21ai_1 _15003_ (.B1(net2649),
    .Y(_06605_),
    .A1(net5083),
    .A2(net1931));
 sg13g2_a21oi_1 _15004_ (.A1(_01774_),
    .A2(net1932),
    .Y(_01061_),
    .B1(_06605_));
 sg13g2_o21ai_1 _15005_ (.B1(net2664),
    .Y(_06606_),
    .A1(net3950),
    .A2(net1932));
 sg13g2_a21oi_1 _15006_ (.A1(_01773_),
    .A2(net1933),
    .Y(_01062_),
    .B1(_06606_));
 sg13g2_o21ai_1 _15007_ (.B1(net2660),
    .Y(_06607_),
    .A1(net3926),
    .A2(net1932));
 sg13g2_a21oi_1 _15008_ (.A1(_01772_),
    .A2(net1933),
    .Y(_01063_),
    .B1(_06607_));
 sg13g2_nand2_1 _15009_ (.Y(_06608_),
    .A(net3785),
    .B(net2661));
 sg13g2_nand2b_1 _15010_ (.Y(_06609_),
    .B(net1932),
    .A_N(_04450_));
 sg13g2_o21ai_1 _15011_ (.B1(_06609_),
    .Y(_01064_),
    .A1(net1932),
    .A2(_06608_));
 sg13g2_o21ai_1 _15012_ (.B1(net2643),
    .Y(_06610_),
    .A1(net4197),
    .A2(net1925));
 sg13g2_a21oi_1 _15013_ (.A1(_01796_),
    .A2(net1925),
    .Y(_01065_),
    .B1(_06610_));
 sg13g2_o21ai_1 _15014_ (.B1(net2647),
    .Y(_06611_),
    .A1(net4267),
    .A2(net1931));
 sg13g2_a21oi_1 _15015_ (.A1(_01795_),
    .A2(net1931),
    .Y(_01066_),
    .B1(_06611_));
 sg13g2_o21ai_1 _15016_ (.B1(net2639),
    .Y(_06612_),
    .A1(net4430),
    .A2(net1924));
 sg13g2_a21oi_1 _15017_ (.A1(_01794_),
    .A2(net1924),
    .Y(_01067_),
    .B1(_06612_));
 sg13g2_o21ai_1 _15018_ (.B1(net2639),
    .Y(_06613_),
    .A1(net5095),
    .A2(net1924));
 sg13g2_a21oi_1 _15019_ (.A1(_01780_),
    .A2(net1924),
    .Y(_01068_),
    .B1(_06613_));
 sg13g2_o21ai_1 _15020_ (.B1(net2643),
    .Y(_06614_),
    .A1(net4221),
    .A2(net1925));
 sg13g2_a21oi_1 _15021_ (.A1(_01793_),
    .A2(net1924),
    .Y(_01069_),
    .B1(_06614_));
 sg13g2_o21ai_1 _15022_ (.B1(net2646),
    .Y(_06615_),
    .A1(net4029),
    .A2(net1931));
 sg13g2_a21oi_1 _15023_ (.A1(_01792_),
    .A2(net1931),
    .Y(_01070_),
    .B1(_06615_));
 sg13g2_o21ai_1 _15024_ (.B1(net2646),
    .Y(_06616_),
    .A1(net4118),
    .A2(net1931));
 sg13g2_a21oi_1 _15025_ (.A1(_01790_),
    .A2(net1931),
    .Y(_01071_),
    .B1(_06616_));
 sg13g2_o21ai_1 _15026_ (.B1(net2647),
    .Y(_06617_),
    .A1(net4005),
    .A2(net1930));
 sg13g2_a21oi_1 _15027_ (.A1(_01842_),
    .A2(net1930),
    .Y(_01072_),
    .B1(_06617_));
 sg13g2_o21ai_1 _15028_ (.B1(net2661),
    .Y(_06618_),
    .A1(net3962),
    .A2(net1929));
 sg13g2_a21oi_1 _15029_ (.A1(_01840_),
    .A2(net1929),
    .Y(_01073_),
    .B1(_06618_));
 sg13g2_o21ai_1 _15030_ (.B1(net2653),
    .Y(_06619_),
    .A1(net4016),
    .A2(net1928));
 sg13g2_a21oi_1 _15031_ (.A1(_01838_),
    .A2(net1929),
    .Y(_01074_),
    .B1(_06619_));
 sg13g2_o21ai_1 _15032_ (.B1(net2653),
    .Y(_06620_),
    .A1(net4317),
    .A2(net1927));
 sg13g2_a21oi_1 _15033_ (.A1(_01836_),
    .A2(net1927),
    .Y(_01075_),
    .B1(_06620_));
 sg13g2_o21ai_1 _15034_ (.B1(net2652),
    .Y(_06621_),
    .A1(net4007),
    .A2(net1928));
 sg13g2_a21oi_1 _15035_ (.A1(_01834_),
    .A2(net1929),
    .Y(_01076_),
    .B1(_06621_));
 sg13g2_o21ai_1 _15036_ (.B1(net2642),
    .Y(_06622_),
    .A1(net4155),
    .A2(net1930));
 sg13g2_a21oi_1 _15037_ (.A1(_01832_),
    .A2(net1930),
    .Y(_01077_),
    .B1(_06622_));
 sg13g2_o21ai_1 _15038_ (.B1(net2651),
    .Y(_06623_),
    .A1(net4098),
    .A2(net1926));
 sg13g2_a21oi_1 _15039_ (.A1(_01830_),
    .A2(net1926),
    .Y(_01078_),
    .B1(_06623_));
 sg13g2_o21ai_1 _15040_ (.B1(net2642),
    .Y(_06624_),
    .A1(net4134),
    .A2(net1930));
 sg13g2_a21oi_1 _15041_ (.A1(_01828_),
    .A2(net1930),
    .Y(_01079_),
    .B1(_06624_));
 sg13g2_o21ai_1 _15042_ (.B1(net2652),
    .Y(_06625_),
    .A1(net4189),
    .A2(net1926));
 sg13g2_a21oi_1 _15043_ (.A1(_01826_),
    .A2(net1926),
    .Y(_01080_),
    .B1(_06625_));
 sg13g2_o21ai_1 _15044_ (.B1(net2653),
    .Y(_06626_),
    .A1(net4393),
    .A2(net1926));
 sg13g2_a21oi_1 _15045_ (.A1(_01824_),
    .A2(net1927),
    .Y(_01081_),
    .B1(_06626_));
 sg13g2_o21ai_1 _15046_ (.B1(net2653),
    .Y(_06627_),
    .A1(net4324),
    .A2(net1927));
 sg13g2_a21oi_1 _15047_ (.A1(_01822_),
    .A2(net1927),
    .Y(_01082_),
    .B1(_06627_));
 sg13g2_o21ai_1 _15048_ (.B1(net2653),
    .Y(_06628_),
    .A1(net4327),
    .A2(net1926));
 sg13g2_a21oi_1 _15049_ (.A1(_01820_),
    .A2(net1927),
    .Y(_01083_),
    .B1(_06628_));
 sg13g2_o21ai_1 _15050_ (.B1(net2651),
    .Y(_06629_),
    .A1(net4071),
    .A2(net1928));
 sg13g2_a21oi_1 _15051_ (.A1(_01818_),
    .A2(net1928),
    .Y(_01084_),
    .B1(_06629_));
 sg13g2_o21ai_1 _15052_ (.B1(net2653),
    .Y(_06630_),
    .A1(net4382),
    .A2(net1927));
 sg13g2_a21oi_1 _15053_ (.A1(_01816_),
    .A2(net1927),
    .Y(_01085_),
    .B1(_06630_));
 sg13g2_o21ai_1 _15054_ (.B1(net2652),
    .Y(_06631_),
    .A1(net4077),
    .A2(net1928));
 sg13g2_a21oi_1 _15055_ (.A1(_01814_),
    .A2(net1928),
    .Y(_01086_),
    .B1(_06631_));
 sg13g2_o21ai_1 _15056_ (.B1(net2654),
    .Y(_06632_),
    .A1(net4227),
    .A2(net1926));
 sg13g2_a21oi_1 _15057_ (.A1(_01812_),
    .A2(net1926),
    .Y(_01087_),
    .B1(_06632_));
 sg13g2_a21oi_1 _15058_ (.A1(_06396_),
    .A2(net1997),
    .Y(_01088_),
    .B1(net2424));
 sg13g2_o21ai_1 _15059_ (.B1(_06384_),
    .Y(_06633_),
    .A1(net2309),
    .A2(net5202));
 sg13g2_and3_1 _15060_ (.X(_01089_),
    .A(net2649),
    .B(_06396_),
    .C(_06633_));
 sg13g2_and4_1 _15061_ (.A(net2637),
    .B(_03465_),
    .C(_04312_),
    .D(_05849_),
    .X(_01090_));
 sg13g2_nor4_2 _15062_ (.A(\i_seal.byte_idx[3] ),
    .B(\i_seal.byte_idx[2] ),
    .C(\i_seal.byte_idx[1] ),
    .Y(_06634_),
    .D(net2493));
 sg13g2_nand2b_2 _15063_ (.Y(_06635_),
    .B(\i_seal.byte_idx[1] ),
    .A_N(net2493));
 sg13g2_nor3_2 _15064_ (.A(\i_seal.byte_idx[3] ),
    .B(\i_seal.byte_idx[2] ),
    .C(_06635_),
    .Y(_06636_));
 sg13g2_nand2b_2 _15065_ (.Y(_06637_),
    .B(net2493),
    .A_N(\i_seal.byte_idx[1] ));
 sg13g2_nor2_2 _15066_ (.A(_06410_),
    .B(_06637_),
    .Y(_06638_));
 sg13g2_nor3_1 _15067_ (.A(_01920_),
    .B(_06410_),
    .C(_06637_),
    .Y(_06639_));
 sg13g2_nor3_2 _15068_ (.A(\i_seal.byte_idx[1] ),
    .B(\i_seal.byte_idx[0] ),
    .C(_06410_),
    .Y(_06640_));
 sg13g2_nor2_2 _15069_ (.A(_06410_),
    .B(_06635_),
    .Y(_06641_));
 sg13g2_nor3_2 _15070_ (.A(\i_seal.byte_idx[3] ),
    .B(\i_seal.byte_idx[2] ),
    .C(_06402_),
    .Y(_06642_));
 sg13g2_nor3_2 _15071_ (.A(\i_seal.byte_idx[3] ),
    .B(\i_seal.byte_idx[2] ),
    .C(_06637_),
    .Y(_06643_));
 sg13g2_a221oi_1 _15072_ (.B2(net3527),
    .C1(_06639_),
    .B1(_06634_),
    .A1(\i_seal.cur_mono[16] ),
    .Y(_06644_),
    .A2(net2219));
 sg13g2_a22oi_1 _15073_ (.Y(_06645_),
    .B1(_06643_),
    .B2(\i_seal.value_reg[0] ),
    .A2(_06387_),
    .A1(\i_seal.cur_mono[24] ));
 sg13g2_a22oi_1 _15074_ (.Y(_06646_),
    .B1(_06641_),
    .B2(\i_seal.cur_mono[8] ),
    .A2(_06640_),
    .A1(\i_seal.value_reg[24] ));
 sg13g2_nand3_1 _15075_ (.B(_06645_),
    .C(_06646_),
    .A(net2220),
    .Y(_06647_));
 sg13g2_a221oi_1 _15076_ (.B2(\i_seal.value_reg[16] ),
    .C1(_06647_),
    .B1(_06642_),
    .A1(net3785),
    .Y(_06648_),
    .A2(_06636_));
 sg13g2_nand2_1 _15077_ (.Y(_06649_),
    .A(net3958),
    .B(net2648));
 sg13g2_a22oi_1 _15078_ (.Y(_01091_),
    .B1(_06649_),
    .B2(_06386_),
    .A2(_06648_),
    .A1(_06644_));
 sg13g2_and2_1 _15079_ (.A(\i_seal.value_reg[9] ),
    .B(_06636_),
    .X(_06650_));
 sg13g2_a221oi_1 _15080_ (.B2(net4147),
    .C1(_06650_),
    .B1(net2219),
    .A1(net3825),
    .Y(_06651_),
    .A2(net2280));
 sg13g2_a22oi_1 _15081_ (.Y(_06652_),
    .B1(_06642_),
    .B2(net3962),
    .A2(_06634_),
    .A1(net3675));
 sg13g2_a22oi_1 _15082_ (.Y(_06653_),
    .B1(_06643_),
    .B2(\i_seal.value_reg[1] ),
    .A2(_06641_),
    .A1(\i_seal.cur_mono[9] ));
 sg13g2_nand3_1 _15083_ (.B(_06652_),
    .C(_06653_),
    .A(net2220),
    .Y(_06654_));
 sg13g2_a221oi_1 _15084_ (.B2(\i_seal.value_reg[25] ),
    .C1(_06654_),
    .B1(_06640_),
    .A1(net4110),
    .Y(_06655_),
    .A2(_06638_));
 sg13g2_nand2_1 _15085_ (.Y(_06656_),
    .A(net4191),
    .B(net2662));
 sg13g2_a22oi_1 _15086_ (.Y(_01092_),
    .B1(_06656_),
    .B2(_06386_),
    .A2(_06655_),
    .A1(_06651_));
 sg13g2_and2_1 _15087_ (.A(\i_seal.value_reg[2] ),
    .B(_06643_),
    .X(_06657_));
 sg13g2_a221oi_1 _15088_ (.B2(net4015),
    .C1(_06657_),
    .B1(net2219),
    .A1(net3982),
    .Y(_06658_),
    .A2(net2280));
 sg13g2_a22oi_1 _15089_ (.Y(_06659_),
    .B1(_06640_),
    .B2(\i_seal.value_reg[26] ),
    .A2(_06636_),
    .A1(net4267));
 sg13g2_a22oi_1 _15090_ (.Y(_06660_),
    .B1(_06642_),
    .B2(net4016),
    .A2(_06641_),
    .A1(\i_seal.cur_mono[10] ));
 sg13g2_nand3_1 _15091_ (.B(_06659_),
    .C(_06660_),
    .A(net2220),
    .Y(_06661_));
 sg13g2_a221oi_1 _15092_ (.B2(net4079),
    .C1(_06661_),
    .B1(_06638_),
    .A1(net3612),
    .Y(_06662_),
    .A2(_06634_));
 sg13g2_nand2_1 _15093_ (.Y(_06663_),
    .A(net4303),
    .B(net2662));
 sg13g2_a22oi_1 _15094_ (.Y(_01093_),
    .B1(_06663_),
    .B2(_06386_),
    .A2(_06662_),
    .A1(_06658_));
 sg13g2_and2_1 _15095_ (.A(\i_seal.value_reg[11] ),
    .B(_06636_),
    .X(_06664_));
 sg13g2_a221oi_1 _15096_ (.B2(\i_seal.value_reg[19] ),
    .C1(_06664_),
    .B1(_06642_),
    .A1(\i_seal.cur_mono[3] ),
    .Y(_06665_),
    .A2(_06638_));
 sg13g2_a22oi_1 _15097_ (.Y(_06666_),
    .B1(_06643_),
    .B2(\i_seal.value_reg[3] ),
    .A2(_06634_),
    .A1(net3645));
 sg13g2_a22oi_1 _15098_ (.Y(_06667_),
    .B1(_06641_),
    .B2(\i_seal.cur_mono[11] ),
    .A2(_06640_),
    .A1(\i_seal.value_reg[27] ));
 sg13g2_nand3_1 _15099_ (.B(_06666_),
    .C(_06667_),
    .A(net2220),
    .Y(_06668_));
 sg13g2_a221oi_1 _15100_ (.B2(net4059),
    .C1(_06668_),
    .B1(net2219),
    .A1(\i_seal.cur_mono[27] ),
    .Y(_06669_),
    .A2(net2280));
 sg13g2_nand2_1 _15101_ (.Y(_06670_),
    .A(net4140),
    .B(net2663));
 sg13g2_a22oi_1 _15102_ (.Y(_01094_),
    .B1(_06670_),
    .B2(_06386_),
    .A2(_06669_),
    .A1(_06665_));
 sg13g2_and2_1 _15103_ (.A(\i_seal.value_reg[12] ),
    .B(_06636_),
    .X(_06671_));
 sg13g2_a221oi_1 _15104_ (.B2(net4007),
    .C1(_06671_),
    .B1(_06642_),
    .A1(net4114),
    .Y(_06672_),
    .A2(_06638_));
 sg13g2_a22oi_1 _15105_ (.Y(_06673_),
    .B1(net2219),
    .B2(\i_seal.cur_mono[20] ),
    .A2(net2280),
    .A1(net3844));
 sg13g2_a22oi_1 _15106_ (.Y(_06674_),
    .B1(_06641_),
    .B2(\i_seal.cur_mono[12] ),
    .A2(_06634_),
    .A1(net3647));
 sg13g2_nand3_1 _15107_ (.B(_06673_),
    .C(_06674_),
    .A(net2220),
    .Y(_06675_));
 sg13g2_a221oi_1 _15108_ (.B2(net3956),
    .C1(_06675_),
    .B1(_06643_),
    .A1(net4071),
    .Y(_06676_),
    .A2(_06640_));
 sg13g2_nand2_1 _15109_ (.Y(_06677_),
    .A(net4213),
    .B(net2662));
 sg13g2_a22oi_1 _15110_ (.Y(_01095_),
    .B1(_06677_),
    .B2(_06386_),
    .A2(_06676_),
    .A1(_06672_));
 sg13g2_nor3_1 _15111_ (.A(_01896_),
    .B(_06410_),
    .C(_06635_),
    .Y(_06678_));
 sg13g2_a221oi_1 _15112_ (.B2(\i_seal.value_reg[29] ),
    .C1(_06678_),
    .B1(_06640_),
    .A1(net4067),
    .Y(_06679_),
    .A2(_06638_));
 sg13g2_a22oi_1 _15113_ (.Y(_06680_),
    .B1(_06634_),
    .B2(net3616),
    .A2(_06387_),
    .A1(net4094));
 sg13g2_a22oi_1 _15114_ (.Y(_06681_),
    .B1(_06643_),
    .B2(\i_seal.value_reg[5] ),
    .A2(net2219),
    .A1(\i_seal.cur_mono[21] ));
 sg13g2_nand3_1 _15115_ (.B(_06680_),
    .C(_06681_),
    .A(net2220),
    .Y(_06682_));
 sg13g2_a221oi_1 _15116_ (.B2(net4155),
    .C1(_06682_),
    .B1(_06642_),
    .A1(net4221),
    .Y(_06683_),
    .A2(_06636_));
 sg13g2_nand2_1 _15117_ (.Y(_06684_),
    .A(net4243),
    .B(net2663));
 sg13g2_a22oi_1 _15118_ (.Y(_01096_),
    .B1(_06684_),
    .B2(_06386_),
    .A2(_06683_),
    .A1(_06679_));
 sg13g2_and2_1 _15119_ (.A(net4029),
    .B(_06636_),
    .X(_06685_));
 sg13g2_a221oi_1 _15120_ (.B2(net4077),
    .C1(_06685_),
    .B1(_06640_),
    .A1(net4576),
    .Y(_06686_),
    .A2(_06638_));
 sg13g2_a22oi_1 _15121_ (.Y(_06687_),
    .B1(_06634_),
    .B2(net3912),
    .A2(net2280),
    .A1(net3846));
 sg13g2_a22oi_1 _15122_ (.Y(_06688_),
    .B1(_06642_),
    .B2(net4098),
    .A2(_06641_),
    .A1(net4777));
 sg13g2_nand3_1 _15123_ (.B(_06687_),
    .C(_06688_),
    .A(_06385_),
    .Y(_06689_));
 sg13g2_a221oi_1 _15124_ (.B2(net3950),
    .C1(_06689_),
    .B1(_06643_),
    .A1(net4559),
    .Y(_06690_),
    .A2(_06411_));
 sg13g2_o21ai_1 _15125_ (.B1(net2660),
    .Y(_06691_),
    .A1(net4907),
    .A2(_06385_));
 sg13g2_a21oi_1 _15126_ (.A1(_06686_),
    .A2(_06690_),
    .Y(_01097_),
    .B1(net4908));
 sg13g2_nor3_1 _15127_ (.A(_01906_),
    .B(_06410_),
    .C(_06637_),
    .Y(_06692_));
 sg13g2_a22oi_1 _15128_ (.Y(_06693_),
    .B1(_06643_),
    .B2(net3926),
    .A2(net2280),
    .A1(\i_seal.cur_mono[31] ));
 sg13g2_a22oi_1 _15129_ (.Y(_06694_),
    .B1(_06641_),
    .B2(\i_seal.cur_mono[15] ),
    .A2(_06640_),
    .A1(\i_seal.value_reg[31] ));
 sg13g2_a221oi_1 _15130_ (.B2(\i_seal.sensor_id_reg[7] ),
    .C1(_06692_),
    .B1(_06634_),
    .A1(\i_seal.cur_mono[23] ),
    .Y(_06695_),
    .A2(net2219));
 sg13g2_nand3_1 _15131_ (.B(_06693_),
    .C(_06694_),
    .A(net2220),
    .Y(_06696_));
 sg13g2_a221oi_1 _15132_ (.B2(\i_seal.value_reg[23] ),
    .C1(_06696_),
    .B1(_06642_),
    .A1(\i_seal.value_reg[15] ),
    .Y(_06697_),
    .A2(_06636_));
 sg13g2_nand2_1 _15133_ (.Y(_06698_),
    .A(net3968),
    .B(net2661));
 sg13g2_a22oi_1 _15134_ (.Y(_01098_),
    .B1(_06698_),
    .B2(_06386_),
    .A2(_06697_),
    .A1(_06695_));
 sg13g2_nand3_1 _15135_ (.B(net2387),
    .C(_02814_),
    .A(\i_tinyqv.cpu.is_load ),
    .Y(_06699_));
 sg13g2_nor2_1 _15136_ (.A(net2002),
    .B(_06699_),
    .Y(_06700_));
 sg13g2_nor2_1 _15137_ (.A(net4353),
    .B(_06700_),
    .Y(_06701_));
 sg13g2_nor3_1 _15138_ (.A(net2345),
    .B(net2002),
    .C(_06699_),
    .Y(_06702_));
 sg13g2_nor3_1 _15139_ (.A(_06408_),
    .B(_06701_),
    .C(_06702_),
    .Y(_01107_));
 sg13g2_o21ai_1 _15140_ (.B1(_06407_),
    .Y(_06703_),
    .A1(net2489),
    .A2(_06700_));
 sg13g2_a21oi_1 _15141_ (.A1(net2310),
    .A2(_06700_),
    .Y(_01108_),
    .B1(_06703_));
 sg13g2_mux2_1 _15142_ (.A0(net2487),
    .A1(_05843_),
    .S(_05870_),
    .X(_01109_));
 sg13g2_mux2_1 _15143_ (.A0(_02689_),
    .A1(_02683_),
    .S(_02791_),
    .X(_06704_));
 sg13g2_nand2_1 _15144_ (.Y(_06705_),
    .A(_05870_),
    .B(_06704_));
 sg13g2_o21ai_1 _15145_ (.B1(_06705_),
    .Y(_01110_),
    .A1(net2409),
    .A2(_05870_));
 sg13g2_nand2b_1 _15146_ (.Y(_06706_),
    .B(_02791_),
    .A_N(_02652_));
 sg13g2_o21ai_1 _15147_ (.B1(_06706_),
    .Y(_06707_),
    .A1(_02640_),
    .A2(_02791_));
 sg13g2_nor2_1 _15148_ (.A(net4568),
    .B(_05870_),
    .Y(_06708_));
 sg13g2_a21oi_1 _15149_ (.A1(_05870_),
    .A2(_06707_),
    .Y(_01111_),
    .B1(_06708_));
 sg13g2_nor2_1 _15150_ (.A(net4416),
    .B(_05870_),
    .Y(_06709_));
 sg13g2_o21ai_1 _15151_ (.B1(_05870_),
    .Y(_06710_),
    .A1(_02571_),
    .A2(_02791_));
 sg13g2_a21oi_1 _15152_ (.A1(_02604_),
    .A2(_02791_),
    .Y(_06711_),
    .B1(_06710_));
 sg13g2_nor2_1 _15153_ (.A(_06709_),
    .B(_06711_),
    .Y(_01112_));
 sg13g2_nand2_1 _15154_ (.Y(_06712_),
    .A(net3682),
    .B(net2355));
 sg13g2_o21ai_1 _15155_ (.B1(_06712_),
    .Y(_01113_),
    .A1(_02061_),
    .A2(net2355));
 sg13g2_mux2_1 _15156_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(net4438),
    .S(net2355),
    .X(_01114_));
 sg13g2_mux2_1 _15157_ (.A0(net4275),
    .A1(net4510),
    .S(net2356),
    .X(_01115_));
 sg13g2_mux2_1 _15158_ (.A0(net4512),
    .A1(net4412),
    .S(net2355),
    .X(_01116_));
 sg13g2_mux2_1 _15159_ (.A0(net3682),
    .A1(net4410),
    .S(net2356),
    .X(_01117_));
 sg13g2_mux2_1 _15160_ (.A0(net4438),
    .A1(net4469),
    .S(net2355),
    .X(_01118_));
 sg13g2_mux2_1 _15161_ (.A0(net4510),
    .A1(\i_tinyqv.cpu.i_core.mepc[10] ),
    .S(net2355),
    .X(_01119_));
 sg13g2_mux2_1 _15162_ (.A0(net4412),
    .A1(net4404),
    .S(net2354),
    .X(_01120_));
 sg13g2_mux2_1 _15163_ (.A0(net4410),
    .A1(\i_tinyqv.cpu.i_core.mepc[12] ),
    .S(net2356),
    .X(_01121_));
 sg13g2_mux2_1 _15164_ (.A0(net4469),
    .A1(net4509),
    .S(net2354),
    .X(_01122_));
 sg13g2_mux2_1 _15165_ (.A0(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A1(net4588),
    .S(net2354),
    .X(_01123_));
 sg13g2_mux2_1 _15166_ (.A0(net4404),
    .A1(\i_tinyqv.cpu.i_core.mepc[15] ),
    .S(net2353),
    .X(_01124_));
 sg13g2_mux2_1 _15167_ (.A0(net4642),
    .A1(\i_tinyqv.cpu.i_core.mepc[16] ),
    .S(net2355),
    .X(_01125_));
 sg13g2_mux2_1 _15168_ (.A0(net4509),
    .A1(net4551),
    .S(net2352),
    .X(_01126_));
 sg13g2_mux2_1 _15169_ (.A0(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A1(net4413),
    .S(net2353),
    .X(_01127_));
 sg13g2_mux2_1 _15170_ (.A0(net4598),
    .A1(net4296),
    .S(net2352),
    .X(_01128_));
 sg13g2_mux2_1 _15171_ (.A0(net4730),
    .A1(net4061),
    .S(net2354),
    .X(_01129_));
 sg13g2_nor2_1 _15172_ (.A(\i_tinyqv.cpu.i_core.mepc[17] ),
    .B(net2352),
    .Y(_06713_));
 sg13g2_a21oi_1 _15173_ (.A1(_02043_),
    .A2(net2352),
    .Y(_01130_),
    .B1(_06713_));
 sg13g2_nor2_1 _15174_ (.A(\i_tinyqv.cpu.i_core.mepc[18] ),
    .B(net2353),
    .Y(_06714_));
 sg13g2_a21oi_1 _15175_ (.A1(_02044_),
    .A2(net2353),
    .Y(_01131_),
    .B1(_06714_));
 sg13g2_nor2_1 _15176_ (.A(net4296),
    .B(net2352),
    .Y(_06715_));
 sg13g2_a21oi_1 _15177_ (.A1(_02045_),
    .A2(net2352),
    .Y(_01132_),
    .B1(_06715_));
 sg13g2_and2_1 _15178_ (.A(_02002_),
    .B(_04653_),
    .X(_06716_));
 sg13g2_mux2_1 _15179_ (.A0(net4584),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net1800),
    .X(_01133_));
 sg13g2_nor2_1 _15180_ (.A(net3984),
    .B(net1801),
    .Y(_06717_));
 sg13g2_a21oi_1 _15181_ (.A1(_02037_),
    .A2(net1801),
    .Y(_01134_),
    .B1(_06717_));
 sg13g2_mux2_1 _15182_ (.A0(net4557),
    .A1(\i_tinyqv.cpu.instr_data_in[4] ),
    .S(net1802),
    .X(_01135_));
 sg13g2_mux2_1 _15183_ (.A0(net4503),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(net1800),
    .X(_01136_));
 sg13g2_mux2_1 _15184_ (.A0(net4657),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net1802),
    .X(_01137_));
 sg13g2_mux2_1 _15185_ (.A0(net4498),
    .A1(\i_tinyqv.cpu.instr_data_in[7] ),
    .S(net1800),
    .X(_01138_));
 sg13g2_nor2_1 _15186_ (.A(net4209),
    .B(net1800),
    .Y(_06718_));
 sg13g2_a21oi_1 _15187_ (.A1(net2410),
    .A2(net1800),
    .Y(_01139_),
    .B1(_06718_));
 sg13g2_mux2_1 _15188_ (.A0(net4452),
    .A1(net2602),
    .S(net1800),
    .X(_01140_));
 sg13g2_mux2_1 _15189_ (.A0(net4582),
    .A1(net2600),
    .S(net1800),
    .X(_01141_));
 sg13g2_mux2_1 _15190_ (.A0(net4496),
    .A1(net2598),
    .S(net1800),
    .X(_01142_));
 sg13g2_mux2_1 _15191_ (.A0(net4454),
    .A1(net2596),
    .S(net1801),
    .X(_01143_));
 sg13g2_mux2_1 _15192_ (.A0(net4505),
    .A1(net2594),
    .S(net1801),
    .X(_01144_));
 sg13g2_mux2_1 _15193_ (.A0(net4570),
    .A1(net2592),
    .S(net1802),
    .X(_01145_));
 sg13g2_mux2_1 _15194_ (.A0(net4492),
    .A1(net2590),
    .S(net1801),
    .X(_01146_));
 sg13g2_nand2_1 _15195_ (.Y(_06719_),
    .A(net2496),
    .B(_04991_));
 sg13g2_o21ai_1 _15196_ (.B1(_06719_),
    .Y(_01147_),
    .A1(_04651_),
    .A2(_04768_));
 sg13g2_nand2_1 _15197_ (.Y(_06720_),
    .A(net2496),
    .B(_05007_));
 sg13g2_o21ai_1 _15198_ (.B1(_06720_),
    .Y(_01148_),
    .A1(_04651_),
    .A2(_04767_));
 sg13g2_nor2_1 _15199_ (.A(_01808_),
    .B(net2240),
    .Y(_06721_));
 sg13g2_and2_1 _15200_ (.A(net2242),
    .B(net2295),
    .X(_06722_));
 sg13g2_a21oi_1 _15201_ (.A1(net4963),
    .A2(_06722_),
    .Y(_06723_),
    .B1(_06721_));
 sg13g2_nor2_1 _15202_ (.A(net2444),
    .B(_06723_),
    .Y(_01149_));
 sg13g2_nor2b_1 _15203_ (.A(net2240),
    .B_N(net5113),
    .Y(_06724_));
 sg13g2_a21oi_1 _15204_ (.A1(net5042),
    .A2(_06722_),
    .Y(_06725_),
    .B1(_06724_));
 sg13g2_nor2_1 _15205_ (.A(net2444),
    .B(_06725_),
    .Y(_01150_));
 sg13g2_nor2b_1 _15206_ (.A(net2240),
    .B_N(net2472),
    .Y(_06726_));
 sg13g2_a21oi_1 _15207_ (.A1(net5004),
    .A2(_06722_),
    .Y(_06727_),
    .B1(_06726_));
 sg13g2_nor2_1 _15208_ (.A(net2449),
    .B(_06727_),
    .Y(_01151_));
 sg13g2_nor2b_1 _15209_ (.A(net2241),
    .B_N(net5172),
    .Y(_06728_));
 sg13g2_a21oi_1 _15210_ (.A1(net5146),
    .A2(_06722_),
    .Y(_06729_),
    .B1(_06728_));
 sg13g2_nor2_1 _15211_ (.A(net2445),
    .B(_06729_),
    .Y(_01152_));
 sg13g2_and2_1 _15212_ (.A(net2501),
    .B(net2240),
    .X(_06730_));
 sg13g2_nor2_1 _15213_ (.A(net5247),
    .B(net2154),
    .Y(_06731_));
 sg13g2_and2_1 _15214_ (.A(net2587),
    .B(_04571_),
    .X(_06732_));
 sg13g2_a21oi_1 _15215_ (.A1(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A2(net2298),
    .Y(_06733_),
    .B1(_06732_));
 sg13g2_a21oi_1 _15216_ (.A1(net2154),
    .A2(_06733_),
    .Y(_01153_),
    .B1(_06731_));
 sg13g2_nor2_1 _15217_ (.A(net5148),
    .B(net2153),
    .Y(_06734_));
 sg13g2_a21oi_1 _15218_ (.A1(_04988_),
    .A2(net2153),
    .Y(_01154_),
    .B1(_06734_));
 sg13g2_nor2_1 _15219_ (.A(net5316),
    .B(net2154),
    .Y(_06735_));
 sg13g2_a21oi_1 _15220_ (.A1(_04999_),
    .A2(net2154),
    .Y(_01155_),
    .B1(_06735_));
 sg13g2_nor2_1 _15221_ (.A(net2466),
    .B(net2155),
    .Y(_06736_));
 sg13g2_a21oi_1 _15222_ (.A1(_05012_),
    .A2(net2155),
    .Y(_01156_),
    .B1(_06736_));
 sg13g2_nor2_1 _15223_ (.A(net4402),
    .B(net2153),
    .Y(_06737_));
 sg13g2_a21oi_1 _15224_ (.A1(_05027_),
    .A2(net2154),
    .Y(_01157_),
    .B1(_06737_));
 sg13g2_mux2_1 _15225_ (.A0(net5263),
    .A1(_05039_),
    .S(net2154),
    .X(_01158_));
 sg13g2_nor2_1 _15226_ (.A(net5052),
    .B(net2153),
    .Y(_06738_));
 sg13g2_a21oi_1 _15227_ (.A1(_05050_),
    .A2(net2154),
    .Y(_01159_),
    .B1(_06738_));
 sg13g2_nor2_1 _15228_ (.A(net4232),
    .B(net2153),
    .Y(_06739_));
 sg13g2_a21oi_1 _15229_ (.A1(_05064_),
    .A2(net2153),
    .Y(_01160_),
    .B1(_06739_));
 sg13g2_nor2_1 _15230_ (.A(net4234),
    .B(net2153),
    .Y(_06740_));
 sg13g2_a21oi_1 _15231_ (.A1(_05077_),
    .A2(net2153),
    .Y(_01161_),
    .B1(_06740_));
 sg13g2_nor2_1 _15232_ (.A(net4342),
    .B(net2152),
    .Y(_06741_));
 sg13g2_a21oi_1 _15233_ (.A1(_05087_),
    .A2(net2152),
    .Y(_01162_),
    .B1(_06741_));
 sg13g2_nor2_1 _15234_ (.A(net4116),
    .B(net2152),
    .Y(_06742_));
 sg13g2_a21oi_1 _15235_ (.A1(_05098_),
    .A2(net2152),
    .Y(_01163_),
    .B1(_06742_));
 sg13g2_nor2_1 _15236_ (.A(net4225),
    .B(net2152),
    .Y(_06743_));
 sg13g2_a21oi_1 _15237_ (.A1(_05115_),
    .A2(net2152),
    .Y(_01164_),
    .B1(_06743_));
 sg13g2_mux2_1 _15238_ (.A0(net4630),
    .A1(_05122_),
    .S(net2155),
    .X(_01165_));
 sg13g2_nor2_1 _15239_ (.A(net4185),
    .B(net2151),
    .Y(_06744_));
 sg13g2_a21oi_1 _15240_ (.A1(_05143_),
    .A2(net2149),
    .Y(_01166_),
    .B1(_06744_));
 sg13g2_nor2_1 _15241_ (.A(net4400),
    .B(net2151),
    .Y(_06745_));
 sg13g2_a21oi_1 _15242_ (.A1(_05155_),
    .A2(net2151),
    .Y(_01167_),
    .B1(_06745_));
 sg13g2_mux2_1 _15243_ (.A0(net4531),
    .A1(_05166_),
    .S(net2149),
    .X(_01168_));
 sg13g2_nor2_1 _15244_ (.A(net4659),
    .B(net2151),
    .Y(_06746_));
 sg13g2_a21oi_1 _15245_ (.A1(_05179_),
    .A2(net2151),
    .Y(_01169_),
    .B1(_06746_));
 sg13g2_mux2_1 _15246_ (.A0(net4537),
    .A1(net4552),
    .S(net2149),
    .X(_01170_));
 sg13g2_nor2_1 _15247_ (.A(net4301),
    .B(net2149),
    .Y(_06747_));
 sg13g2_a21oi_1 _15248_ (.A1(_05207_),
    .A2(net2149),
    .Y(_01171_),
    .B1(_06747_));
 sg13g2_mux2_1 _15249_ (.A0(net4578),
    .A1(_05216_),
    .S(net2149),
    .X(_01172_));
 sg13g2_nor2_1 _15250_ (.A(net4779),
    .B(net2150),
    .Y(_06748_));
 sg13g2_a21oi_1 _15251_ (.A1(_05230_),
    .A2(net2149),
    .Y(_01173_),
    .B1(_06748_));
 sg13g2_mux2_1 _15252_ (.A0(net4766),
    .A1(_05242_),
    .S(net2150),
    .X(_01174_));
 sg13g2_nor2_1 _15253_ (.A(net4299),
    .B(net2149),
    .Y(_06749_));
 sg13g2_a21oi_1 _15254_ (.A1(_05254_),
    .A2(net2150),
    .Y(_01175_),
    .B1(_06749_));
 sg13g2_nor2_1 _15255_ (.A(net4599),
    .B(net2152),
    .Y(_06750_));
 sg13g2_a21oi_1 _15256_ (.A1(_05266_),
    .A2(net2150),
    .Y(_01176_),
    .B1(_06750_));
 sg13g2_nand2b_1 _15257_ (.Y(_06751_),
    .B(\i_spi.clock_count[0] ),
    .A_N(\i_spi.clock_divider[0] ));
 sg13g2_a22oi_1 _15258_ (.Y(_06752_),
    .B1(\i_spi.clock_divider[0] ),
    .B2(_01749_),
    .A2(_01978_),
    .A1(\i_spi.clock_count[3] ));
 sg13g2_xnor2_1 _15259_ (.Y(_06753_),
    .A(\i_spi.clock_count[2] ),
    .B(\i_spi.clock_divider[2] ));
 sg13g2_o21ai_1 _15260_ (.B1(net2454),
    .Y(_06754_),
    .A1(_01748_),
    .A2(\i_spi.clock_divider[1] ));
 sg13g2_a221oi_1 _15261_ (.B2(_01748_),
    .C1(_06754_),
    .B1(\i_spi.clock_divider[1] ),
    .A1(_01746_),
    .Y(_06755_),
    .A2(\i_spi.clock_divider[3] ));
 sg13g2_nand4_1 _15262_ (.B(_06752_),
    .C(_06753_),
    .A(_06751_),
    .Y(_06756_),
    .D(_06755_));
 sg13g2_nand2_1 _15263_ (.Y(_06757_),
    .A(net2326),
    .B(net2082));
 sg13g2_nor2_1 _15264_ (.A(net2458),
    .B(_06757_),
    .Y(_06758_));
 sg13g2_inv_2 _15265_ (.Y(_06759_),
    .A(_06758_));
 sg13g2_nand2_2 _15266_ (.Y(_06760_),
    .A(_06756_),
    .B(_06759_));
 sg13g2_o21ai_1 _15267_ (.B1(_06760_),
    .Y(_06761_),
    .A1(net5007),
    .A2(_01747_));
 sg13g2_inv_1 _15268_ (.Y(_06762_),
    .A(_06761_));
 sg13g2_nand2_2 _15269_ (.Y(_06763_),
    .A(net2628),
    .B(_06762_));
 sg13g2_nand2b_1 _15270_ (.Y(_06764_),
    .B(net2457),
    .A_N(\i_spi.data[0] ));
 sg13g2_o21ai_1 _15271_ (.B1(_06764_),
    .Y(_06765_),
    .A1(net2457),
    .A2(net2557));
 sg13g2_nand2_1 _15272_ (.Y(_06766_),
    .A(net3629),
    .B(net1888));
 sg13g2_o21ai_1 _15273_ (.B1(_06766_),
    .Y(_01177_),
    .A1(net1888),
    .A2(_06765_));
 sg13g2_nand2b_1 _15274_ (.Y(_06767_),
    .B(net2456),
    .A_N(net3629));
 sg13g2_o21ai_1 _15275_ (.B1(_06767_),
    .Y(_06768_),
    .A1(net2456),
    .A2(net2556));
 sg13g2_nand2_1 _15276_ (.Y(_06769_),
    .A(net3649),
    .B(net1887));
 sg13g2_o21ai_1 _15277_ (.B1(_06769_),
    .Y(_01178_),
    .A1(net1887),
    .A2(_06768_));
 sg13g2_nand2b_1 _15278_ (.Y(_06770_),
    .B(net2455),
    .A_N(net3649));
 sg13g2_o21ai_1 _15279_ (.B1(_06770_),
    .Y(_06771_),
    .A1(net2455),
    .A2(\crc_peri_data[3] ));
 sg13g2_nand2_1 _15280_ (.Y(_06772_),
    .A(net3670),
    .B(net1887));
 sg13g2_o21ai_1 _15281_ (.B1(_06772_),
    .Y(_01179_),
    .A1(net1887),
    .A2(_06771_));
 sg13g2_nand2b_1 _15282_ (.Y(_06773_),
    .B(net2455),
    .A_N(\i_spi.data[3] ));
 sg13g2_o21ai_1 _15283_ (.B1(_06773_),
    .Y(_06774_),
    .A1(net2456),
    .A2(\crc_peri_data[4] ));
 sg13g2_nand2_1 _15284_ (.Y(_06775_),
    .A(net3643),
    .B(net1887));
 sg13g2_o21ai_1 _15285_ (.B1(_06775_),
    .Y(_01180_),
    .A1(net1887),
    .A2(_06774_));
 sg13g2_nand2b_1 _15286_ (.Y(_06776_),
    .B(net2455),
    .A_N(net3643));
 sg13g2_o21ai_1 _15287_ (.B1(_06776_),
    .Y(_06777_),
    .A1(net2455),
    .A2(\crc_peri_data[5] ));
 sg13g2_nand2_1 _15288_ (.Y(_06778_),
    .A(net3659),
    .B(net1887));
 sg13g2_o21ai_1 _15289_ (.B1(_06778_),
    .Y(_01181_),
    .A1(net1888),
    .A2(_06777_));
 sg13g2_nand2b_1 _15290_ (.Y(_06779_),
    .B(net2455),
    .A_N(net3659));
 sg13g2_o21ai_1 _15291_ (.B1(_06779_),
    .Y(_06780_),
    .A1(net2456),
    .A2(net2552));
 sg13g2_nand2_1 _15292_ (.Y(_06781_),
    .A(net3850),
    .B(net1887));
 sg13g2_o21ai_1 _15293_ (.B1(_06781_),
    .Y(_01182_),
    .A1(net1888),
    .A2(_06780_));
 sg13g2_nand2b_1 _15294_ (.Y(_06782_),
    .B(net2455),
    .A_N(\i_spi.data[6] ));
 sg13g2_o21ai_1 _15295_ (.B1(_06782_),
    .Y(_06783_),
    .A1(net2455),
    .A2(\crc_peri_data[7] ));
 sg13g2_nand2_1 _15296_ (.Y(_06784_),
    .A(net3716),
    .B(_06763_));
 sg13g2_o21ai_1 _15297_ (.B1(_06784_),
    .Y(_01183_),
    .A1(_06763_),
    .A2(_06783_));
 sg13g2_nand2_2 _15298_ (.Y(_06785_),
    .A(net2467),
    .B(_02756_));
 sg13g2_inv_1 _15299_ (.Y(_06786_),
    .A(_06785_));
 sg13g2_nand4_1 _15300_ (.B(net4949),
    .C(net5122),
    .A(net2472),
    .Y(_06787_),
    .D(_02755_));
 sg13g2_o21ai_1 _15301_ (.B1(_06787_),
    .Y(_06788_),
    .A1(_02755_),
    .A2(_06785_));
 sg13g2_nand2_1 _15302_ (.Y(_06789_),
    .A(net2635),
    .B(_06788_));
 sg13g2_a21oi_2 _15303_ (.B1(_06789_),
    .Y(_01184_),
    .A2(_06785_),
    .A1(net2402));
 sg13g2_nand3_1 _15304_ (.B(net2081),
    .C(_05849_),
    .A(_01797_),
    .Y(_06790_));
 sg13g2_o21ai_1 _15305_ (.B1(_06790_),
    .Y(_06791_),
    .A1(_02025_),
    .A2(_03463_));
 sg13g2_nand2_1 _15306_ (.Y(_06792_),
    .A(net2308),
    .B(net1923));
 sg13g2_nand2b_1 _15307_ (.Y(_06793_),
    .B(net4170),
    .A_N(_03536_));
 sg13g2_a21oi_1 _15308_ (.A1(_06792_),
    .A2(_06793_),
    .Y(_01185_),
    .B1(net1956));
 sg13g2_mux2_1 _15309_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(net4545),
    .S(net1803),
    .X(_01186_));
 sg13g2_nand2_1 _15310_ (.Y(_06794_),
    .A(net3636),
    .B(net1803));
 sg13g2_o21ai_1 _15311_ (.B1(_06794_),
    .Y(_01187_),
    .A1(_02037_),
    .A2(net1803));
 sg13g2_mux2_1 _15312_ (.A0(\i_tinyqv.cpu.instr_data_in[4] ),
    .A1(net4590),
    .S(net1804),
    .X(_01188_));
 sg13g2_mux2_1 _15313_ (.A0(\i_tinyqv.cpu.instr_data_in[5] ),
    .A1(net4518),
    .S(net1803),
    .X(_01189_));
 sg13g2_mux2_1 _15314_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(net4621),
    .S(net1804),
    .X(_01190_));
 sg13g2_mux2_1 _15315_ (.A0(\i_tinyqv.cpu.instr_data_in[7] ),
    .A1(net4574),
    .S(net1803),
    .X(_01191_));
 sg13g2_nand2_1 _15316_ (.Y(_06795_),
    .A(net3693),
    .B(net1804));
 sg13g2_o21ai_1 _15317_ (.B1(_06795_),
    .Y(_01192_),
    .A1(net2410),
    .A2(net1804));
 sg13g2_mux2_1 _15318_ (.A0(net2602),
    .A1(net4473),
    .S(net1803),
    .X(_01193_));
 sg13g2_mux2_1 _15319_ (.A0(net2600),
    .A1(net4668),
    .S(net1804),
    .X(_01194_));
 sg13g2_mux2_1 _15320_ (.A0(net2598),
    .A1(net4523),
    .S(net1803),
    .X(_01195_));
 sg13g2_mux2_1 _15321_ (.A0(net2596),
    .A1(net4644),
    .S(net1803),
    .X(_01196_));
 sg13g2_mux2_1 _15322_ (.A0(net2594),
    .A1(net4601),
    .S(net1804),
    .X(_01197_));
 sg13g2_mux2_1 _15323_ (.A0(net2592),
    .A1(net4458),
    .S(net1805),
    .X(_01198_));
 sg13g2_mux2_1 _15324_ (.A0(net2590),
    .A1(net4525),
    .S(net1805),
    .X(_01199_));
 sg13g2_a21oi_1 _15325_ (.A1(_04649_),
    .A2(_04763_),
    .Y(_06796_),
    .B1(net2442));
 sg13g2_nand3_1 _15326_ (.B(_04649_),
    .C(_04763_),
    .A(net2496),
    .Y(_06797_));
 sg13g2_nor2_1 _15327_ (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .B(net1839),
    .Y(_06798_));
 sg13g2_a21oi_1 _15328_ (.A1(_02007_),
    .A2(_06796_),
    .Y(_01200_),
    .B1(_06798_));
 sg13g2_nor2_1 _15329_ (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .B(net1839),
    .Y(_06799_));
 sg13g2_a21oi_1 _15330_ (.A1(_02010_),
    .A2(_06796_),
    .Y(_01201_),
    .B1(_06799_));
 sg13g2_nand3_1 _15331_ (.B(_05354_),
    .C(net2332),
    .A(_05353_),
    .Y(_06800_));
 sg13g2_and2_1 _15332_ (.A(net2623),
    .B(_06800_),
    .X(_01202_));
 sg13g2_nand2_1 _15333_ (.Y(_06801_),
    .A(\i_i2c_peri.i_i2c.addr_reg[6] ),
    .B(_05381_));
 sg13g2_mux2_1 _15334_ (.A0(\i_i2c_peri.i_i2c.addr_reg[4] ),
    .A1(\i_i2c_peri.i_i2c.addr_reg[5] ),
    .S(net2507),
    .X(_06802_));
 sg13g2_and3_1 _15335_ (.X(_06803_),
    .A(net2506),
    .B(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .C(_06802_));
 sg13g2_nand2b_1 _15336_ (.Y(_06804_),
    .B(net2507),
    .A_N(\i_i2c_peri.i_i2c.addr_reg[1] ));
 sg13g2_o21ai_1 _15337_ (.B1(_06804_),
    .Y(_06805_),
    .A1(net2507),
    .A2(\i_i2c_peri.i_i2c.addr_reg[0] ));
 sg13g2_nand2_1 _15338_ (.Y(_06806_),
    .A(net2507),
    .B(\i_i2c_peri.i_i2c.addr_reg[3] ));
 sg13g2_a21oi_1 _15339_ (.A1(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .A2(_06806_),
    .Y(_06807_),
    .B1(net2506));
 sg13g2_a21oi_1 _15340_ (.A1(\i_i2c_peri.i_i2c.addr_reg[2] ),
    .A2(_05380_),
    .Y(_06808_),
    .B1(_06807_));
 sg13g2_o21ai_1 _15341_ (.B1(_06808_),
    .Y(_06809_),
    .A1(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .A2(_06805_));
 sg13g2_o21ai_1 _15342_ (.B1(_02023_),
    .Y(_06810_),
    .A1(_06803_),
    .A2(_06809_));
 sg13g2_a221oi_1 _15343_ (.B2(_06810_),
    .C1(_05392_),
    .B1(_06801_),
    .A1(_02016_),
    .Y(_06811_),
    .A2(_05382_));
 sg13g2_nand2b_1 _15344_ (.Y(_06812_),
    .B(\i_i2c_peri.i_i2c.data_reg[7] ),
    .A_N(_05382_));
 sg13g2_or2_1 _15345_ (.X(_06813_),
    .B(\i_i2c_peri.i_i2c.data_reg[5] ),
    .A(net2508));
 sg13g2_o21ai_1 _15346_ (.B1(_06813_),
    .Y(_06814_),
    .A1(\i_i2c_peri.i_i2c.bit_count_reg[1] ),
    .A2(\i_i2c_peri.i_i2c.data_reg[4] ));
 sg13g2_and3_1 _15347_ (.X(_06815_),
    .A(net2508),
    .B(net2506),
    .C(_02033_));
 sg13g2_a221oi_1 _15348_ (.B2(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .C1(_06815_),
    .B1(_06814_),
    .A1(_05380_),
    .Y(_06816_),
    .A2(_06812_));
 sg13g2_mux4_1 _15349_ (.S0(\i_i2c_peri.i_i2c.bit_count_reg[1] ),
    .A0(_02030_),
    .A1(_02028_),
    .A2(_02027_),
    .A3(_02029_),
    .S1(net2508),
    .X(_06817_));
 sg13g2_nand3_1 _15350_ (.B(_05386_),
    .C(_05890_),
    .A(_01966_),
    .Y(_06818_));
 sg13g2_a21oi_1 _15351_ (.A1(_05889_),
    .A2(_06817_),
    .Y(_06819_),
    .B1(_06818_));
 sg13g2_o21ai_1 _15352_ (.B1(_06819_),
    .Y(_06820_),
    .A1(_05889_),
    .A2(_06816_));
 sg13g2_or2_1 _15353_ (.X(_06821_),
    .B(_05418_),
    .A(_05358_));
 sg13g2_nand2_1 _15354_ (.Y(_06822_),
    .A(_05441_),
    .B(_06821_));
 sg13g2_a21oi_1 _15355_ (.A1(_05384_),
    .A2(net2222),
    .Y(_06823_),
    .B1(_05393_));
 sg13g2_and2_1 _15356_ (.A(_05424_),
    .B(_06823_),
    .X(_06824_));
 sg13g2_nand4_1 _15357_ (.B(_06820_),
    .C(_06822_),
    .A(_05389_),
    .Y(_06825_),
    .D(_06824_));
 sg13g2_nor3_1 _15358_ (.A(_05434_),
    .B(_06811_),
    .C(_06825_),
    .Y(_06826_));
 sg13g2_nor2_1 _15359_ (.A(_05365_),
    .B(_06826_),
    .Y(_06827_));
 sg13g2_nor3_1 _15360_ (.A(net4885),
    .B(\i_i2c_peri.i_i2c.delay_reg[1] ),
    .C(\i_i2c_peri.i_i2c.delay_reg[0] ),
    .Y(_06828_));
 sg13g2_nor2b_1 _15361_ (.A(net4760),
    .B_N(_06828_),
    .Y(_06829_));
 sg13g2_nor2b_1 _15362_ (.A(net4695),
    .B_N(_06829_),
    .Y(_06830_));
 sg13g2_nor2b_1 _15363_ (.A(net4871),
    .B_N(_06830_),
    .Y(_06831_));
 sg13g2_nor2b_2 _15364_ (.A(net4906),
    .B_N(_06831_),
    .Y(_06832_));
 sg13g2_nor4_1 _15365_ (.A(net4490),
    .B(net4618),
    .C(net4700),
    .D(net4245),
    .Y(_06833_));
 sg13g2_nand2_2 _15366_ (.Y(_06834_),
    .A(_06832_),
    .B(_06833_));
 sg13g2_nor3_1 _15367_ (.A(net4073),
    .B(\i_i2c_peri.i_i2c.delay_reg[11] ),
    .C(_06834_),
    .Y(_06835_));
 sg13g2_nand2b_1 _15368_ (.Y(_06836_),
    .B(_06835_),
    .A_N(net3722));
 sg13g2_nor2_2 _15369_ (.A(net4182),
    .B(\i_i2c_peri.i_i2c.delay_reg[15] ),
    .Y(_06837_));
 sg13g2_nor2_1 _15370_ (.A(net3876),
    .B(_06836_),
    .Y(_06838_));
 sg13g2_and2_1 _15371_ (.A(_06837_),
    .B(_06838_),
    .X(_06839_));
 sg13g2_nand2_1 _15372_ (.Y(_06840_),
    .A(_06837_),
    .B(_06838_));
 sg13g2_or2_1 _15373_ (.X(_06841_),
    .B(net5357),
    .A(net3409));
 sg13g2_nor2_2 _15374_ (.A(net1899),
    .B(_06841_),
    .Y(_06842_));
 sg13g2_or2_1 _15375_ (.X(_06843_),
    .B(_06841_),
    .A(net1899));
 sg13g2_nand2_1 _15376_ (.Y(_06844_),
    .A(net2464),
    .B(_01804_));
 sg13g2_nand2_1 _15377_ (.Y(_06845_),
    .A(net2461),
    .B(net2462));
 sg13g2_nand2_1 _15378_ (.Y(_06846_),
    .A(_05363_),
    .B(_06844_));
 sg13g2_o21ai_1 _15379_ (.B1(_06846_),
    .Y(_06847_),
    .A1(_06844_),
    .A2(_06845_));
 sg13g2_nor3_1 _15380_ (.A(net2545),
    .B(_05383_),
    .C(_05387_),
    .Y(_06848_));
 sg13g2_nor3_1 _15381_ (.A(_05391_),
    .B(_05441_),
    .C(_06848_),
    .Y(_06849_));
 sg13g2_nand2_1 _15382_ (.Y(_06850_),
    .A(_05389_),
    .B(_06849_));
 sg13g2_a21oi_1 _15383_ (.A1(_01966_),
    .A2(_05398_),
    .Y(_06851_),
    .B1(_05399_));
 sg13g2_a21oi_1 _15384_ (.A1(_05377_),
    .A2(_05379_),
    .Y(_06852_),
    .B1(_06851_));
 sg13g2_inv_1 _15385_ (.Y(_06853_),
    .A(_06852_));
 sg13g2_a21oi_1 _15386_ (.A1(_05364_),
    .A2(_06853_),
    .Y(_06854_),
    .B1(_06850_));
 sg13g2_nand2_1 _15387_ (.Y(_06855_),
    .A(net5159),
    .B(net2332));
 sg13g2_inv_1 _15388_ (.Y(_06856_),
    .A(_06855_));
 sg13g2_nand3_1 _15389_ (.B(_06854_),
    .C(_06856_),
    .A(_06824_),
    .Y(_06857_));
 sg13g2_nor2_1 _15390_ (.A(_05434_),
    .B(_06857_),
    .Y(_06858_));
 sg13g2_nor2_1 _15391_ (.A(_06841_),
    .B(_06858_),
    .Y(_06859_));
 sg13g2_nand3_1 _15392_ (.B(_06847_),
    .C(_06859_),
    .A(_06839_),
    .Y(_06860_));
 sg13g2_nand2_1 _15393_ (.Y(_06861_),
    .A(_01804_),
    .B(_05435_));
 sg13g2_inv_1 _15394_ (.Y(_06862_),
    .A(_06861_));
 sg13g2_o21ai_1 _15395_ (.B1(_06861_),
    .Y(_06863_),
    .A1(_01804_),
    .A2(_06827_));
 sg13g2_a21oi_1 _15396_ (.A1(net4823),
    .A2(_06860_),
    .Y(_06864_),
    .B1(net2412));
 sg13g2_o21ai_1 _15397_ (.B1(_06864_),
    .Y(_01203_),
    .A1(_06860_),
    .A2(_06863_));
 sg13g2_nor3_1 _15398_ (.A(net2461),
    .B(net2464),
    .C(\i_i2c_peri.i_i2c.phy_state_reg[0] ),
    .Y(_06865_));
 sg13g2_nand2_1 _15399_ (.Y(_06866_),
    .A(net2462),
    .B(_06865_));
 sg13g2_nand2_1 _15400_ (.Y(_06867_),
    .A(net2464),
    .B(net5372));
 sg13g2_nand2b_1 _15401_ (.Y(_06868_),
    .B(_06845_),
    .A_N(_06867_));
 sg13g2_nor2_1 _15402_ (.A(_05363_),
    .B(_06868_),
    .Y(_06869_));
 sg13g2_a21oi_1 _15403_ (.A1(net2462),
    .A2(_06865_),
    .Y(_06870_),
    .B1(_06869_));
 sg13g2_inv_1 _15404_ (.Y(_06871_),
    .A(_06870_));
 sg13g2_nand3b_1 _15405_ (.B(net5159),
    .C(net5349),
    .Y(_06872_),
    .A_N(net4377));
 sg13g2_inv_1 _15406_ (.Y(_06873_),
    .A(_06872_));
 sg13g2_nor2_1 _15407_ (.A(net2461),
    .B(_06844_),
    .Y(_06874_));
 sg13g2_nor2_1 _15408_ (.A(_06873_),
    .B(_06874_),
    .Y(_06875_));
 sg13g2_o21ai_1 _15409_ (.B1(_06875_),
    .Y(_06876_),
    .A1(\i_i2c_peri.i_i2c.phy_state_reg[0] ),
    .A2(_05365_));
 sg13g2_o21ai_1 _15410_ (.B1(_06842_),
    .Y(_06877_),
    .A1(_06871_),
    .A2(_06876_));
 sg13g2_a21oi_1 _15411_ (.A1(net4445),
    .A2(_06877_),
    .Y(_06878_),
    .B1(net2412));
 sg13g2_o21ai_1 _15412_ (.B1(_06878_),
    .Y(_01204_),
    .A1(_06871_),
    .A2(_06877_));
 sg13g2_nor4_2 _15413_ (.A(_01966_),
    .B(_05365_),
    .C(_05384_),
    .Y(_06879_),
    .D(_05387_));
 sg13g2_mux2_1 _15414_ (.A0(net4161),
    .A1(\i_i2c_peri.i_i2c.phy_rx_data_reg ),
    .S(_06879_),
    .X(_01205_));
 sg13g2_nor2_1 _15415_ (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[1] ),
    .B(net2189),
    .Y(_06880_));
 sg13g2_a21oi_1 _15416_ (.A1(_02027_),
    .A2(net2188),
    .Y(_01206_),
    .B1(_06880_));
 sg13g2_nor2_1 _15417_ (.A(net3948),
    .B(net2189),
    .Y(_06881_));
 sg13g2_a21oi_1 _15418_ (.A1(_02028_),
    .A2(net2188),
    .Y(_01207_),
    .B1(_06881_));
 sg13g2_nor2_1 _15419_ (.A(net4261),
    .B(net2188),
    .Y(_06882_));
 sg13g2_a21oi_1 _15420_ (.A1(_02029_),
    .A2(net2188),
    .Y(_01208_),
    .B1(_06882_));
 sg13g2_nor2_1 _15421_ (.A(net4207),
    .B(net2188),
    .Y(_06883_));
 sg13g2_a21oi_1 _15422_ (.A1(_02030_),
    .A2(net2188),
    .Y(_01209_),
    .B1(_06883_));
 sg13g2_nor2_1 _15423_ (.A(net4108),
    .B(net2188),
    .Y(_06884_));
 sg13g2_a21oi_1 _15424_ (.A1(_02031_),
    .A2(net2188),
    .Y(_01210_),
    .B1(_06884_));
 sg13g2_nor2_1 _15425_ (.A(net4057),
    .B(net2189),
    .Y(_06885_));
 sg13g2_a21oi_1 _15426_ (.A1(_02032_),
    .A2(net2189),
    .Y(_01211_),
    .B1(_06885_));
 sg13g2_nor2_1 _15427_ (.A(net3831),
    .B(net2190),
    .Y(_06886_));
 sg13g2_a21oi_1 _15428_ (.A1(_02033_),
    .A2(net2190),
    .Y(_01212_),
    .B1(_06886_));
 sg13g2_a21oi_1 _15429_ (.A1(\i_i2c_peri.i_i2c.sda_o_reg ),
    .A2(_02022_),
    .Y(_06887_),
    .B1(\i_i2c_peri.i_i2c.delay_scl_reg ));
 sg13g2_nor3_1 _15430_ (.A(_01806_),
    .B(net2412),
    .C(_06887_),
    .Y(_01213_));
 sg13g2_nand3_1 _15431_ (.B(net2464),
    .C(_01804_),
    .A(net2461),
    .Y(_06888_));
 sg13g2_nor3_1 _15432_ (.A(net2462),
    .B(_06843_),
    .C(net4378),
    .Y(_06889_));
 sg13g2_nor2_1 _15433_ (.A(net4329),
    .B(_06889_),
    .Y(_06890_));
 sg13g2_a21oi_1 _15434_ (.A1(_02022_),
    .A2(_06889_),
    .Y(_01214_),
    .B1(_06890_));
 sg13g2_nand2_1 _15435_ (.Y(_06891_),
    .A(\i_i2c_peri.i_i2c.bus_active_reg ),
    .B(net3631));
 sg13g2_o21ai_1 _15436_ (.B1(net2621),
    .Y(_06892_),
    .A1(\i_i2c_peri.i_i2c.bus_active_reg ),
    .A2(net3631));
 sg13g2_a21oi_1 _15437_ (.A1(net3397),
    .A2(net3632),
    .Y(_01215_),
    .B1(_06892_));
 sg13g2_nor2_1 _15438_ (.A(_05359_),
    .B(_06800_),
    .Y(_06893_));
 sg13g2_nor2_1 _15439_ (.A(\i_i2c_peri.i_i2c.mode_stop_reg ),
    .B(net2187),
    .Y(_06894_));
 sg13g2_a21oi_1 _15440_ (.A1(_01789_),
    .A2(net2187),
    .Y(_01216_),
    .B1(_06894_));
 sg13g2_nand2b_1 _15441_ (.Y(_01217_),
    .B(net2622),
    .A_N(net5));
 sg13g2_nand2b_1 _15442_ (.Y(_01218_),
    .B(net2622),
    .A_N(net3594));
 sg13g2_or2_1 _15443_ (.X(_06895_),
    .B(_05443_),
    .A(_05365_));
 sg13g2_mux2_1 _15444_ (.A0(\i_i2c_peri.i_i2c.s_axis_data_tlast ),
    .A1(net4165),
    .S(_06895_),
    .X(_01219_));
 sg13g2_o21ai_1 _15445_ (.B1(\i_i2c_peri.rx_has_data ),
    .Y(_06896_),
    .A1(_03444_),
    .A2(_06699_));
 sg13g2_inv_1 _15446_ (.Y(_06897_),
    .A(_06896_));
 sg13g2_a21oi_1 _15447_ (.A1(net4271),
    .A2(_06897_),
    .Y(_06898_),
    .B1(net4711));
 sg13g2_nor2_1 _15448_ (.A(net2413),
    .B(net4712),
    .Y(_01220_));
 sg13g2_nand2_1 _15449_ (.Y(_06899_),
    .A(_06844_),
    .B(_06872_));
 sg13g2_nor2_1 _15450_ (.A(_05363_),
    .B(_06899_),
    .Y(_06900_));
 sg13g2_a22oi_1 _15451_ (.Y(_06901_),
    .B1(_06870_),
    .B2(_06900_),
    .A2(net2332),
    .A1(_01804_));
 sg13g2_o21ai_1 _15452_ (.B1(_06859_),
    .Y(_06902_),
    .A1(_06862_),
    .A2(_06901_));
 sg13g2_o21ai_1 _15453_ (.B1(_06902_),
    .Y(_06903_),
    .A1(_06839_),
    .A2(_06841_));
 sg13g2_and2_1 _15454_ (.A(net2463),
    .B(_06874_),
    .X(_06904_));
 sg13g2_nand2_1 _15455_ (.Y(_06905_),
    .A(net2463),
    .B(_06874_));
 sg13g2_a21oi_1 _15456_ (.A1(net4651),
    .A2(net2144),
    .Y(_06906_),
    .B1(net1897));
 sg13g2_o21ai_1 _15457_ (.B1(net1894),
    .Y(_06907_),
    .A1(net4999),
    .A2(_06906_));
 sg13g2_o21ai_1 _15458_ (.B1(_06907_),
    .Y(_06908_),
    .A1(net4999),
    .A2(net1894));
 sg13g2_nor2_1 _15459_ (.A(net2414),
    .B(_06908_),
    .Y(_01221_));
 sg13g2_xnor2_1 _15460_ (.Y(_06909_),
    .A(net4935),
    .B(\i_i2c_peri.i_i2c.delay_reg[0] ));
 sg13g2_nand2_1 _15461_ (.Y(_06910_),
    .A(net4651),
    .B(net2148));
 sg13g2_o21ai_1 _15462_ (.B1(_06910_),
    .Y(_06911_),
    .A1(_01802_),
    .A2(net2147));
 sg13g2_o21ai_1 _15463_ (.B1(_06909_),
    .Y(_06912_),
    .A1(net1897),
    .A2(_06911_));
 sg13g2_o21ai_1 _15464_ (.B1(net2627),
    .Y(_06913_),
    .A1(net4935),
    .A2(net1894));
 sg13g2_a21oi_1 _15465_ (.A1(net1894),
    .A2(_06912_),
    .Y(_01222_),
    .B1(_06913_));
 sg13g2_o21ai_1 _15466_ (.B1(net4885),
    .Y(_06914_),
    .A1(\i_i2c_peri.i_i2c.delay_reg[1] ),
    .A2(\i_i2c_peri.i_i2c.delay_reg[0] ));
 sg13g2_nand2b_1 _15467_ (.Y(_06915_),
    .B(_06914_),
    .A_N(_06828_));
 sg13g2_a21oi_1 _15468_ (.A1(\i2c_config_out[2] ),
    .A2(net2144),
    .Y(_06916_),
    .B1(net1897));
 sg13g2_o21ai_1 _15469_ (.B1(_06916_),
    .Y(_06917_),
    .A1(_01802_),
    .A2(net2144));
 sg13g2_nand2_1 _15470_ (.Y(_06918_),
    .A(_06915_),
    .B(_06917_));
 sg13g2_o21ai_1 _15471_ (.B1(net2628),
    .Y(_06919_),
    .A1(net4885),
    .A2(net1894));
 sg13g2_a21oi_1 _15472_ (.A1(net1894),
    .A2(_06918_),
    .Y(_01223_),
    .B1(_06919_));
 sg13g2_nor2b_1 _15473_ (.A(_06828_),
    .B_N(net4760),
    .Y(_06920_));
 sg13g2_a21oi_1 _15474_ (.A1(\i2c_config_out[3] ),
    .A2(net2145),
    .Y(_06921_),
    .B1(net1897));
 sg13g2_o21ai_1 _15475_ (.B1(_06921_),
    .Y(_06922_),
    .A1(_01801_),
    .A2(net2145));
 sg13g2_o21ai_1 _15476_ (.B1(_06922_),
    .Y(_06923_),
    .A1(_06829_),
    .A2(_06920_));
 sg13g2_o21ai_1 _15477_ (.B1(net2627),
    .Y(_06924_),
    .A1(net4760),
    .A2(net1895));
 sg13g2_a21oi_1 _15478_ (.A1(net1895),
    .A2(_06923_),
    .Y(_01224_),
    .B1(_06924_));
 sg13g2_nor2b_1 _15479_ (.A(_06829_),
    .B_N(net4695),
    .Y(_06925_));
 sg13g2_a21oi_1 _15480_ (.A1(\i2c_config_out[4] ),
    .A2(net2145),
    .Y(_06926_),
    .B1(net1897));
 sg13g2_o21ai_1 _15481_ (.B1(_06926_),
    .Y(_06927_),
    .A1(_01800_),
    .A2(net2145));
 sg13g2_o21ai_1 _15482_ (.B1(_06927_),
    .Y(_06928_),
    .A1(_06830_),
    .A2(_06925_));
 sg13g2_o21ai_1 _15483_ (.B1(net2627),
    .Y(_06929_),
    .A1(net4695),
    .A2(net1895));
 sg13g2_a21oi_1 _15484_ (.A1(net1895),
    .A2(_06928_),
    .Y(_01225_),
    .B1(_06929_));
 sg13g2_nor2b_1 _15485_ (.A(_06830_),
    .B_N(net4871),
    .Y(_06930_));
 sg13g2_a21oi_1 _15486_ (.A1(\i2c_config_out[5] ),
    .A2(net2145),
    .Y(_06931_),
    .B1(net1898));
 sg13g2_o21ai_1 _15487_ (.B1(_06931_),
    .Y(_06932_),
    .A1(_01799_),
    .A2(net2145));
 sg13g2_o21ai_1 _15488_ (.B1(_06932_),
    .Y(_06933_),
    .A1(_06831_),
    .A2(_06930_));
 sg13g2_o21ai_1 _15489_ (.B1(net2627),
    .Y(_06934_),
    .A1(net4871),
    .A2(net1896));
 sg13g2_a21oi_1 _15490_ (.A1(net1896),
    .A2(_06933_),
    .Y(_01226_),
    .B1(_06934_));
 sg13g2_nor2b_1 _15491_ (.A(_06831_),
    .B_N(net4906),
    .Y(_06935_));
 sg13g2_a21oi_1 _15492_ (.A1(net4898),
    .A2(net2146),
    .Y(_06936_),
    .B1(net1898));
 sg13g2_o21ai_1 _15493_ (.B1(_06936_),
    .Y(_06937_),
    .A1(_01798_),
    .A2(net2146));
 sg13g2_o21ai_1 _15494_ (.B1(_06937_),
    .Y(_06938_),
    .A1(_06832_),
    .A2(_06935_));
 sg13g2_o21ai_1 _15495_ (.B1(net2627),
    .Y(_06939_),
    .A1(net4906),
    .A2(net1893));
 sg13g2_a21oi_1 _15496_ (.A1(net1896),
    .A2(_06938_),
    .Y(_01227_),
    .B1(_06939_));
 sg13g2_nand2_1 _15497_ (.Y(_06940_),
    .A(_06832_),
    .B(net1893));
 sg13g2_or2_1 _15498_ (.X(_06941_),
    .B(_06940_),
    .A(net4245));
 sg13g2_nand2_1 _15499_ (.Y(_06942_),
    .A(net4245),
    .B(_06940_));
 sg13g2_a21o_1 _15500_ (.A2(net2146),
    .A1(\i2c_config_out[7] ),
    .B1(net1898),
    .X(_06943_));
 sg13g2_a21oi_1 _15501_ (.A1(\i2c_config_out[6] ),
    .A2(net2147),
    .Y(_06944_),
    .B1(_06943_));
 sg13g2_a221oi_1 _15502_ (.B2(net1893),
    .C1(net2411),
    .B1(_06944_),
    .A1(_06941_),
    .Y(_01228_),
    .A2(net4246));
 sg13g2_or2_1 _15503_ (.X(_06945_),
    .B(_06941_),
    .A(net4700));
 sg13g2_nand2_1 _15504_ (.Y(_06946_),
    .A(net4700),
    .B(_06941_));
 sg13g2_and2_1 _15505_ (.A(\i2c_config_out[8] ),
    .B(net2146),
    .X(_06947_));
 sg13g2_a21oi_1 _15506_ (.A1(\i2c_config_out[7] ),
    .A2(net2147),
    .Y(_06948_),
    .B1(_06947_));
 sg13g2_nor2_2 _15507_ (.A(net1899),
    .B(_06902_),
    .Y(_06949_));
 sg13g2_a221oi_1 _15508_ (.B2(_06949_),
    .C1(net2412),
    .B1(_06948_),
    .A1(_06945_),
    .Y(_01229_),
    .A2(_06946_));
 sg13g2_or3_1 _15509_ (.A(net4618),
    .B(\i_i2c_peri.i_i2c.delay_reg[8] ),
    .C(_06941_),
    .X(_06950_));
 sg13g2_o21ai_1 _15510_ (.B1(net4618),
    .Y(_06951_),
    .A1(\i_i2c_peri.i_i2c.delay_reg[8] ),
    .A2(_06941_));
 sg13g2_nand2b_1 _15511_ (.Y(_06952_),
    .B(net2144),
    .A_N(\i2c_config_out[9] ));
 sg13g2_o21ai_1 _15512_ (.B1(_06952_),
    .Y(_06953_),
    .A1(\i2c_config_out[8] ),
    .A2(net2144));
 sg13g2_a221oi_1 _15513_ (.B2(_06949_),
    .C1(net2411),
    .B1(_06953_),
    .A1(_06950_),
    .Y(_01230_),
    .A2(net4619));
 sg13g2_nand2_1 _15514_ (.Y(_06954_),
    .A(\i2c_config_out[10] ),
    .B(net2144));
 sg13g2_a21oi_1 _15515_ (.A1(\i2c_config_out[9] ),
    .A2(net2147),
    .Y(_06955_),
    .B1(net1897));
 sg13g2_a21oi_1 _15516_ (.A1(_06954_),
    .A2(_06955_),
    .Y(_06956_),
    .B1(_06834_));
 sg13g2_a22oi_1 _15517_ (.Y(_06957_),
    .B1(_06956_),
    .B2(net1893),
    .A2(_06950_),
    .A1(net4490));
 sg13g2_nor2_1 _15518_ (.A(net2411),
    .B(net4491),
    .Y(_01231_));
 sg13g2_mux2_1 _15519_ (.A0(\i2c_config_out[11] ),
    .A1(\i2c_config_out[10] ),
    .S(net2147),
    .X(_06958_));
 sg13g2_xnor2_1 _15520_ (.Y(_06959_),
    .A(net4899),
    .B(_06834_));
 sg13g2_o21ai_1 _15521_ (.B1(_06959_),
    .Y(_06960_),
    .A1(net1897),
    .A2(_06958_));
 sg13g2_o21ai_1 _15522_ (.B1(net2627),
    .Y(_06961_),
    .A1(net4899),
    .A2(net1894));
 sg13g2_a21oi_1 _15523_ (.A1(net1894),
    .A2(_06960_),
    .Y(_01232_),
    .B1(_06961_));
 sg13g2_nand2_1 _15524_ (.Y(_06962_),
    .A(_06835_),
    .B(net1893));
 sg13g2_nor3_1 _15525_ (.A(_01805_),
    .B(\i_i2c_peri.i_i2c.delay_reg[11] ),
    .C(_06834_),
    .Y(_06963_));
 sg13g2_nand2_1 _15526_ (.Y(_06964_),
    .A(\i2c_config_out[11] ),
    .B(net2147));
 sg13g2_a21oi_1 _15527_ (.A1(\i2c_config_out[12] ),
    .A2(net2144),
    .Y(_06965_),
    .B1(net1897));
 sg13g2_a21o_1 _15528_ (.A2(_06965_),
    .A1(_06964_),
    .B1(_06963_),
    .X(_06966_));
 sg13g2_a221oi_1 _15529_ (.B2(net1893),
    .C1(net2411),
    .B1(_06966_),
    .A1(_01805_),
    .Y(_01233_),
    .A2(_06962_));
 sg13g2_and2_1 _15530_ (.A(\i2c_config_out[12] ),
    .B(net2148),
    .X(_06967_));
 sg13g2_a21oi_1 _15531_ (.A1(\i2c_config_out[13] ),
    .A2(net2144),
    .Y(_06968_),
    .B1(_06967_));
 sg13g2_nand2b_1 _15532_ (.Y(_06969_),
    .B(net1893),
    .A_N(_06836_));
 sg13g2_a21oi_1 _15533_ (.A1(_06839_),
    .A2(_06968_),
    .Y(_06970_),
    .B1(_06969_));
 sg13g2_a21oi_1 _15534_ (.A1(net3722),
    .A2(_06962_),
    .Y(_06971_),
    .B1(_06970_));
 sg13g2_nor2_1 _15535_ (.A(net2411),
    .B(net3723),
    .Y(_01234_));
 sg13g2_o21ai_1 _15536_ (.B1(_06837_),
    .Y(_06972_),
    .A1(_01791_),
    .A2(net2147));
 sg13g2_a21oi_1 _15537_ (.A1(\i2c_config_out[13] ),
    .A2(net2147),
    .Y(_06973_),
    .B1(_06972_));
 sg13g2_nand2_1 _15538_ (.Y(_06974_),
    .A(_06838_),
    .B(net1893));
 sg13g2_nor2_1 _15539_ (.A(_06973_),
    .B(_06974_),
    .Y(_06975_));
 sg13g2_a21oi_1 _15540_ (.A1(net3876),
    .A2(_06969_),
    .Y(_06976_),
    .B1(_06975_));
 sg13g2_nor2_1 _15541_ (.A(net2411),
    .B(net3877),
    .Y(_01235_));
 sg13g2_xor2_1 _15542_ (.B(_06974_),
    .A(\i_i2c_peri.i_i2c.delay_reg[15] ),
    .X(_06977_));
 sg13g2_o21ai_1 _15543_ (.B1(_06837_),
    .Y(_06978_),
    .A1(_01791_),
    .A2(net2146));
 sg13g2_a21oi_1 _15544_ (.A1(net4923),
    .A2(net2146),
    .Y(_06979_),
    .B1(_06978_));
 sg13g2_nor3_1 _15545_ (.A(net2411),
    .B(_06977_),
    .C(net4924),
    .Y(_01236_));
 sg13g2_o21ai_1 _15546_ (.B1(net4182),
    .Y(_06980_),
    .A1(\i_i2c_peri.i_i2c.delay_reg[15] ),
    .A2(_06974_));
 sg13g2_nand3_1 _15547_ (.B(net2148),
    .C(_06949_),
    .A(\i2c_config_out[15] ),
    .Y(_06981_));
 sg13g2_a21oi_1 _15548_ (.A1(net4183),
    .A2(_06981_),
    .Y(_01237_),
    .B1(net2411));
 sg13g2_o21ai_1 _15549_ (.B1(net5159),
    .Y(_06982_),
    .A1(net2461),
    .A2(net2464));
 sg13g2_o21ai_1 _15550_ (.B1(_05364_),
    .Y(_06983_),
    .A1(_05434_),
    .A2(_06850_));
 sg13g2_a22oi_1 _15551_ (.Y(_06984_),
    .B1(_06983_),
    .B2(_06856_),
    .A2(_06982_),
    .A1(_05365_));
 sg13g2_o21ai_1 _15552_ (.B1(net2624),
    .Y(_06985_),
    .A1(net5159),
    .A2(_06842_));
 sg13g2_a21oi_1 _15553_ (.A1(_06842_),
    .A2(_06984_),
    .Y(_01238_),
    .B1(net5160));
 sg13g2_nor2_1 _15554_ (.A(_06855_),
    .B(_06983_),
    .Y(_06986_));
 sg13g2_nor3_1 _15555_ (.A(_06843_),
    .B(_06899_),
    .C(_06986_),
    .Y(_06987_));
 sg13g2_o21ai_1 _15556_ (.B1(net2624),
    .Y(_06988_),
    .A1(net2464),
    .A2(_06842_));
 sg13g2_nor2_1 _15557_ (.A(_06987_),
    .B(_06988_),
    .Y(_01239_));
 sg13g2_nand2_1 _15558_ (.Y(_06989_),
    .A(_06872_),
    .B(_06888_));
 sg13g2_nand2_1 _15559_ (.Y(_06990_),
    .A(net2463),
    .B(_06989_));
 sg13g2_o21ai_1 _15560_ (.B1(_06866_),
    .Y(_06991_),
    .A1(net2462),
    .A2(_06867_));
 sg13g2_o21ai_1 _15561_ (.B1(_06990_),
    .Y(_06992_),
    .A1(_06854_),
    .A2(_06855_));
 sg13g2_nor4_1 _15562_ (.A(_06862_),
    .B(net2148),
    .C(_06991_),
    .D(_06992_),
    .Y(_06993_));
 sg13g2_o21ai_1 _15563_ (.B1(net2624),
    .Y(_06994_),
    .A1(net2462),
    .A2(_06842_));
 sg13g2_a21oi_1 _15564_ (.A1(_06842_),
    .A2(_06993_),
    .Y(_01240_),
    .B1(_06994_));
 sg13g2_a21oi_1 _15565_ (.A1(_06824_),
    .A2(_06852_),
    .Y(_06995_),
    .B1(_06855_));
 sg13g2_nor3_1 _15566_ (.A(_06869_),
    .B(_06989_),
    .C(_06995_),
    .Y(_06996_));
 sg13g2_o21ai_1 _15567_ (.B1(net2624),
    .Y(_06997_),
    .A1(net2461),
    .A2(_06842_));
 sg13g2_a21oi_1 _15568_ (.A1(_06842_),
    .A2(_06996_),
    .Y(_01241_),
    .B1(net5350));
 sg13g2_nor2_1 _15569_ (.A(net3650),
    .B(net2187),
    .Y(_06998_));
 sg13g2_a21oi_1 _15570_ (.A1(\i_i2c_peri.cmd_read_reg ),
    .A2(net2187),
    .Y(_01242_),
    .B1(_06998_));
 sg13g2_nor2_1 _15571_ (.A(net3770),
    .B(net2185),
    .Y(_06999_));
 sg13g2_a21oi_1 _15572_ (.A1(_01788_),
    .A2(net2185),
    .Y(_01243_),
    .B1(_06999_));
 sg13g2_nor2_1 _15573_ (.A(net4255),
    .B(net2185),
    .Y(_07000_));
 sg13g2_a21oi_1 _15574_ (.A1(_01787_),
    .A2(net2185),
    .Y(_01244_),
    .B1(_07000_));
 sg13g2_nor2_1 _15575_ (.A(net4241),
    .B(net2186),
    .Y(_07001_));
 sg13g2_a21oi_1 _15576_ (.A1(_01786_),
    .A2(net2186),
    .Y(_01245_),
    .B1(_07001_));
 sg13g2_nor2_1 _15577_ (.A(net4127),
    .B(net2185),
    .Y(_07002_));
 sg13g2_a21oi_1 _15578_ (.A1(_01785_),
    .A2(net2186),
    .Y(_01246_),
    .B1(_07002_));
 sg13g2_nor2_1 _15579_ (.A(\i_i2c_peri.i_i2c.addr_reg[4] ),
    .B(net2185),
    .Y(_07003_));
 sg13g2_a21oi_1 _15580_ (.A1(_01784_),
    .A2(net2186),
    .Y(_01247_),
    .B1(_07003_));
 sg13g2_nor2_1 _15581_ (.A(net4248),
    .B(net2186),
    .Y(_07004_));
 sg13g2_a21oi_1 _15582_ (.A1(_01783_),
    .A2(net2186),
    .Y(_01248_),
    .B1(_07004_));
 sg13g2_nor2_1 _15583_ (.A(net3805),
    .B(net2185),
    .Y(_07005_));
 sg13g2_a21oi_1 _15584_ (.A1(_01782_),
    .A2(net2185),
    .Y(_01249_),
    .B1(_07005_));
 sg13g2_mux2_1 _15585_ (.A0(net4566),
    .A1(\i_i2c_peri.cmd_read_reg ),
    .S(net2187),
    .X(_01250_));
 sg13g2_nor3_1 _15586_ (.A(net2413),
    .B(_06843_),
    .C(_06875_),
    .Y(_01251_));
 sg13g2_nand2_1 _15587_ (.Y(_07006_),
    .A(net3479),
    .B(_05974_));
 sg13g2_nand3_1 _15588_ (.B(net1860),
    .C(net1834),
    .A(\addr[0] ),
    .Y(_07007_));
 sg13g2_nand2_1 _15589_ (.Y(_01252_),
    .A(_07006_),
    .B(_07007_));
 sg13g2_mux2_1 _15590_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(net4549),
    .S(net1837),
    .X(_01253_));
 sg13g2_nand2_1 _15591_ (.Y(_07008_),
    .A(net3729),
    .B(net1837));
 sg13g2_o21ai_1 _15592_ (.B1(_07008_),
    .Y(_01254_),
    .A1(_02037_),
    .A2(net1837));
 sg13g2_mux2_1 _15593_ (.A0(\i_tinyqv.cpu.instr_data_in[4] ),
    .A1(net4666),
    .S(net1838),
    .X(_01255_));
 sg13g2_mux2_1 _15594_ (.A0(\i_tinyqv.cpu.instr_data_in[5] ),
    .A1(net4448),
    .S(net1837),
    .X(_01256_));
 sg13g2_mux2_1 _15595_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(net4494),
    .S(net1838),
    .X(_01257_));
 sg13g2_mux2_1 _15596_ (.A0(\i_tinyqv.cpu.instr_data_in[7] ),
    .A1(net4427),
    .S(net1837),
    .X(_01258_));
 sg13g2_nand2_1 _15597_ (.Y(_07009_),
    .A(net3802),
    .B(net1838));
 sg13g2_o21ai_1 _15598_ (.B1(_07009_),
    .Y(_01259_),
    .A1(net2410),
    .A2(net1838));
 sg13g2_mux2_1 _15599_ (.A0(net2602),
    .A1(net4407),
    .S(net1837),
    .X(_01260_));
 sg13g2_mux2_1 _15600_ (.A0(net2600),
    .A1(net4661),
    .S(net1838),
    .X(_01261_));
 sg13g2_mux2_1 _15601_ (.A0(net2598),
    .A1(net4424),
    .S(net1837),
    .X(_01262_));
 sg13g2_mux2_1 _15602_ (.A0(net2596),
    .A1(net4487),
    .S(net1837),
    .X(_01263_));
 sg13g2_mux2_1 _15603_ (.A0(net2594),
    .A1(net4616),
    .S(net1838),
    .X(_01264_));
 sg13g2_mux2_1 _15604_ (.A0(net2592),
    .A1(net4547),
    .S(net1839),
    .X(_01265_));
 sg13g2_mux2_1 _15605_ (.A0(net2590),
    .A1(net4634),
    .S(net1839),
    .X(_01266_));
 sg13g2_nor3_1 _15606_ (.A(net2325),
    .B(_03442_),
    .C(_03452_),
    .Y(_07010_));
 sg13g2_nand2_2 _15607_ (.Y(_07011_),
    .A(net2326),
    .B(net2079));
 sg13g2_a21oi_1 _15608_ (.A1(net2559),
    .A2(net2048),
    .Y(_07012_),
    .B1(net2414));
 sg13g2_o21ai_1 _15609_ (.B1(_07012_),
    .Y(_01267_),
    .A1(_01803_),
    .A2(net2049));
 sg13g2_a21oi_1 _15610_ (.A1(net2557),
    .A2(net2047),
    .Y(_07013_),
    .B1(net2414));
 sg13g2_o21ai_1 _15611_ (.B1(_07013_),
    .Y(_01268_),
    .A1(_01802_),
    .A2(net2047));
 sg13g2_a21oi_1 _15612_ (.A1(net4954),
    .A2(_07011_),
    .Y(_07014_),
    .B1(net2414));
 sg13g2_o21ai_1 _15613_ (.B1(_07014_),
    .Y(_01269_),
    .A1(_01777_),
    .A2(_07011_));
 sg13g2_a21oi_1 _15614_ (.A1(net4805),
    .A2(_07011_),
    .Y(_07015_),
    .B1(net2414));
 sg13g2_o21ai_1 _15615_ (.B1(_07015_),
    .Y(_01270_),
    .A1(_01776_),
    .A2(_07011_));
 sg13g2_a21oi_1 _15616_ (.A1(net4862),
    .A2(_07011_),
    .Y(_07016_),
    .B1(net2412));
 sg13g2_o21ai_1 _15617_ (.B1(_07016_),
    .Y(_01271_),
    .A1(_01775_),
    .A2(_07011_));
 sg13g2_a21oi_1 _15618_ (.A1(net4897),
    .A2(_07011_),
    .Y(_07017_),
    .B1(net2412));
 sg13g2_o21ai_1 _15619_ (.B1(_07017_),
    .Y(_01272_),
    .A1(_01774_),
    .A2(_07011_));
 sg13g2_o21ai_1 _15620_ (.B1(net2626),
    .Y(_07018_),
    .A1(net4898),
    .A2(net2050));
 sg13g2_a21oi_1 _15621_ (.A1(_01773_),
    .A2(net2050),
    .Y(_01273_),
    .B1(_07018_));
 sg13g2_o21ai_1 _15622_ (.B1(net2626),
    .Y(_07019_),
    .A1(net4931),
    .A2(net2050));
 sg13g2_a21oi_1 _15623_ (.A1(_01772_),
    .A2(net2050),
    .Y(_01274_),
    .B1(_07019_));
 sg13g2_o21ai_1 _15624_ (.B1(net2627),
    .Y(_07020_),
    .A1(net5110),
    .A2(net2050));
 sg13g2_a21oi_1 _15625_ (.A1(_01797_),
    .A2(net2050),
    .Y(_01275_),
    .B1(_07020_));
 sg13g2_o21ai_1 _15626_ (.B1(net2631),
    .Y(_07021_),
    .A1(net5078),
    .A2(net2047));
 sg13g2_a21oi_1 _15627_ (.A1(_01796_),
    .A2(net2047),
    .Y(_01276_),
    .B1(_07021_));
 sg13g2_o21ai_1 _15628_ (.B1(net2631),
    .Y(_07022_),
    .A1(net5081),
    .A2(net2049));
 sg13g2_a21oi_1 _15629_ (.A1(_01795_),
    .A2(net2048),
    .Y(_01277_),
    .B1(_07022_));
 sg13g2_o21ai_1 _15630_ (.B1(net2631),
    .Y(_07023_),
    .A1(net5002),
    .A2(net2048));
 sg13g2_a21oi_1 _15631_ (.A1(_01794_),
    .A2(net2048),
    .Y(_01278_),
    .B1(_07023_));
 sg13g2_o21ai_1 _15632_ (.B1(net2627),
    .Y(_07024_),
    .A1(net5126),
    .A2(net2047));
 sg13g2_a21oi_1 _15633_ (.A1(_01780_),
    .A2(net2047),
    .Y(_01279_),
    .B1(_07024_));
 sg13g2_o21ai_1 _15634_ (.B1(net2631),
    .Y(_07025_),
    .A1(net5118),
    .A2(net2048));
 sg13g2_a21oi_1 _15635_ (.A1(_01793_),
    .A2(net2048),
    .Y(_01280_),
    .B1(_07025_));
 sg13g2_o21ai_1 _15636_ (.B1(net2631),
    .Y(_07026_),
    .A1(net5086),
    .A2(net2047));
 sg13g2_a21oi_1 _15637_ (.A1(_01792_),
    .A2(net2047),
    .Y(_01281_),
    .B1(_07026_));
 sg13g2_o21ai_1 _15638_ (.B1(net2631),
    .Y(_07027_),
    .A1(net4923),
    .A2(net2048));
 sg13g2_a21oi_1 _15639_ (.A1(_01790_),
    .A2(net2048),
    .Y(_01282_),
    .B1(_07027_));
 sg13g2_nor2_2 _15640_ (.A(net2325),
    .B(_03444_),
    .Y(_07028_));
 sg13g2_nand2_2 _15641_ (.Y(_07029_),
    .A(net2550),
    .B(_07028_));
 sg13g2_nand2_1 _15642_ (.Y(_07030_),
    .A(net5188),
    .B(net1904));
 sg13g2_nor4_2 _15643_ (.A(_02014_),
    .B(net2325),
    .C(_03474_),
    .Y(_07031_),
    .D(_03475_));
 sg13g2_o21ai_1 _15644_ (.B1(_07030_),
    .Y(_07032_),
    .A1(_01779_),
    .A2(net1904));
 sg13g2_and2_1 _15645_ (.A(net2618),
    .B(_07032_),
    .X(_01283_));
 sg13g2_nand2_1 _15646_ (.Y(_07033_),
    .A(net5169),
    .B(net1904));
 sg13g2_o21ai_1 _15647_ (.B1(_07033_),
    .Y(_07034_),
    .A1(net2452),
    .A2(net1904));
 sg13g2_and2_1 _15648_ (.A(net2618),
    .B(_07034_),
    .X(_01284_));
 sg13g2_nand2_1 _15649_ (.Y(_07035_),
    .A(net5206),
    .B(net1905));
 sg13g2_o21ai_1 _15650_ (.B1(_07035_),
    .Y(_07036_),
    .A1(_01777_),
    .A2(net1905));
 sg13g2_and2_1 _15651_ (.A(net2615),
    .B(_07036_),
    .X(_01285_));
 sg13g2_nand2_1 _15652_ (.Y(_07037_),
    .A(net5200),
    .B(net1904));
 sg13g2_o21ai_1 _15653_ (.B1(_07037_),
    .Y(_07038_),
    .A1(net2453),
    .A2(net1905));
 sg13g2_and2_1 _15654_ (.A(net2615),
    .B(_07038_),
    .X(_01286_));
 sg13g2_nand2_1 _15655_ (.Y(_07039_),
    .A(net4292),
    .B(net1905));
 sg13g2_o21ai_1 _15656_ (.B1(_07039_),
    .Y(_07040_),
    .A1(_01775_),
    .A2(net1905));
 sg13g2_and2_1 _15657_ (.A(net2615),
    .B(_07040_),
    .X(_01287_));
 sg13g2_nand2_1 _15658_ (.Y(_07041_),
    .A(net5147),
    .B(net1904));
 sg13g2_o21ai_1 _15659_ (.B1(_07041_),
    .Y(_07042_),
    .A1(_01774_),
    .A2(net1905));
 sg13g2_and2_1 _15660_ (.A(net2615),
    .B(_07042_),
    .X(_01288_));
 sg13g2_nand2_1 _15661_ (.Y(_07043_),
    .A(net5139),
    .B(net1904));
 sg13g2_o21ai_1 _15662_ (.B1(_07043_),
    .Y(_07044_),
    .A1(_01773_),
    .A2(net1904));
 sg13g2_and2_1 _15663_ (.A(net2618),
    .B(_07044_),
    .X(_01289_));
 sg13g2_nor2_1 _15664_ (.A(_04309_),
    .B(_07029_),
    .Y(_07045_));
 sg13g2_a21o_1 _15665_ (.A2(_04310_),
    .A1(net2547),
    .B1(net2548),
    .X(_07046_));
 sg13g2_a21oi_1 _15666_ (.A1(_07028_),
    .A2(_07046_),
    .Y(_07047_),
    .B1(_07045_));
 sg13g2_or2_1 _15667_ (.X(_07048_),
    .B(_07047_),
    .A(net4055));
 sg13g2_nand3b_1 _15668_ (.B(_07031_),
    .C(net2550),
    .Y(_07049_),
    .A_N(_04309_));
 sg13g2_and2_1 _15669_ (.A(net2547),
    .B(_07031_),
    .X(_07050_));
 sg13g2_a22oi_1 _15670_ (.Y(_07051_),
    .B1(_07050_),
    .B2(_04310_),
    .A2(_07031_),
    .A1(net2548));
 sg13g2_a21oi_2 _15671_ (.B1(net4055),
    .Y(_07052_),
    .A2(_07051_),
    .A1(_07049_));
 sg13g2_nand4_1 _15672_ (.B(_07031_),
    .C(_07049_),
    .A(net2548),
    .Y(_07053_),
    .D(_07052_));
 sg13g2_o21ai_1 _15673_ (.B1(net2623),
    .Y(_07054_),
    .A1(net2547),
    .A2(_07053_));
 sg13g2_a21oi_1 _15674_ (.A1(_01789_),
    .A2(net1892),
    .Y(_01290_),
    .B1(_07054_));
 sg13g2_o21ai_1 _15675_ (.B1(net2623),
    .Y(_07055_),
    .A1(net4903),
    .A2(_07052_));
 sg13g2_a21oi_1 _15676_ (.A1(_07049_),
    .A2(_07052_),
    .Y(_01291_),
    .B1(_07055_));
 sg13g2_nand2_1 _15677_ (.Y(_07056_),
    .A(net4723),
    .B(net1892));
 sg13g2_a21oi_1 _15678_ (.A1(_07053_),
    .A2(_07056_),
    .Y(_01292_),
    .B1(net2413));
 sg13g2_o21ai_1 _15679_ (.B1(net2619),
    .Y(_07057_),
    .A1(net4975),
    .A2(_07052_));
 sg13g2_a21oi_1 _15680_ (.A1(_01797_),
    .A2(_07052_),
    .Y(_01293_),
    .B1(_07057_));
 sg13g2_o21ai_1 _15681_ (.B1(net2618),
    .Y(_07058_),
    .A1(_07032_),
    .A2(net1890));
 sg13g2_a21oi_1 _15682_ (.A1(_01788_),
    .A2(net1890),
    .Y(_01294_),
    .B1(_07058_));
 sg13g2_o21ai_1 _15683_ (.B1(net2618),
    .Y(_07059_),
    .A1(_07034_),
    .A2(net1890));
 sg13g2_a21oi_1 _15684_ (.A1(_01787_),
    .A2(net1890),
    .Y(_01295_),
    .B1(_07059_));
 sg13g2_o21ai_1 _15685_ (.B1(net2615),
    .Y(_07060_),
    .A1(_07036_),
    .A2(net1891));
 sg13g2_a21oi_1 _15686_ (.A1(_01786_),
    .A2(net1890),
    .Y(_01296_),
    .B1(_07060_));
 sg13g2_o21ai_1 _15687_ (.B1(net2615),
    .Y(_07061_),
    .A1(_07038_),
    .A2(net1890));
 sg13g2_a21oi_1 _15688_ (.A1(_01785_),
    .A2(net1891),
    .Y(_01297_),
    .B1(_07061_));
 sg13g2_o21ai_1 _15689_ (.B1(net2615),
    .Y(_07062_),
    .A1(_07040_),
    .A2(net1891));
 sg13g2_a21oi_1 _15690_ (.A1(_01784_),
    .A2(net1891),
    .Y(_01298_),
    .B1(_07062_));
 sg13g2_o21ai_1 _15691_ (.B1(net2615),
    .Y(_07063_),
    .A1(_07042_),
    .A2(net1891));
 sg13g2_a21oi_1 _15692_ (.A1(_01783_),
    .A2(net1891),
    .Y(_01299_),
    .B1(_07063_));
 sg13g2_o21ai_1 _15693_ (.B1(net2618),
    .Y(_07064_),
    .A1(_07044_),
    .A2(net1890));
 sg13g2_a21oi_1 _15694_ (.A1(_01782_),
    .A2(net1890),
    .Y(_01300_),
    .B1(_07064_));
 sg13g2_nand2_1 _15695_ (.Y(_07065_),
    .A(net2623),
    .B(_05357_));
 sg13g2_a21oi_1 _15696_ (.A1(_01781_),
    .A2(_07047_),
    .Y(_01301_),
    .B1(_07065_));
 sg13g2_nor3_1 _15697_ (.A(\i_i2c_peri.tx_pending ),
    .B(net2550),
    .C(_04309_),
    .Y(_07066_));
 sg13g2_and2_1 _15698_ (.A(_07028_),
    .B(_07066_),
    .X(_07067_));
 sg13g2_o21ai_1 _15699_ (.B1(net2619),
    .Y(_07068_),
    .A1(net4612),
    .A2(net1903));
 sg13g2_a21oi_1 _15700_ (.A1(_01780_),
    .A2(net1903),
    .Y(_01302_),
    .B1(_07068_));
 sg13g2_o21ai_1 _15701_ (.B1(net2616),
    .Y(_07069_),
    .A1(net4470),
    .A2(net1901));
 sg13g2_a21oi_1 _15702_ (.A1(_01779_),
    .A2(net1901),
    .Y(_01303_),
    .B1(_07069_));
 sg13g2_o21ai_1 _15703_ (.B1(net2616),
    .Y(_07070_),
    .A1(net4729),
    .A2(net1900));
 sg13g2_a21oi_1 _15704_ (.A1(net2452),
    .A2(net1901),
    .Y(_01304_),
    .B1(_07070_));
 sg13g2_o21ai_1 _15705_ (.B1(net2616),
    .Y(_07071_),
    .A1(net4725),
    .A2(net1900));
 sg13g2_a21oi_1 _15706_ (.A1(_01777_),
    .A2(net1900),
    .Y(_01305_),
    .B1(_07071_));
 sg13g2_o21ai_1 _15707_ (.B1(net2616),
    .Y(_07072_),
    .A1(net4767),
    .A2(net1900));
 sg13g2_a21oi_1 _15708_ (.A1(net2453),
    .A2(net1900),
    .Y(_01306_),
    .B1(_07072_));
 sg13g2_o21ai_1 _15709_ (.B1(net2616),
    .Y(_07073_),
    .A1(net4749),
    .A2(net1900));
 sg13g2_a21oi_1 _15710_ (.A1(_01775_),
    .A2(net1901),
    .Y(_01307_),
    .B1(_07073_));
 sg13g2_o21ai_1 _15711_ (.B1(net2616),
    .Y(_07074_),
    .A1(net4812),
    .A2(net1900));
 sg13g2_a21oi_1 _15712_ (.A1(_01774_),
    .A2(net1900),
    .Y(_01308_),
    .B1(_07074_));
 sg13g2_o21ai_1 _15713_ (.B1(net2616),
    .Y(_07075_),
    .A1(net4507),
    .A2(net1902));
 sg13g2_a21oi_1 _15714_ (.A1(_01773_),
    .A2(net1902),
    .Y(_01309_),
    .B1(_07075_));
 sg13g2_o21ai_1 _15715_ (.B1(net2619),
    .Y(_07076_),
    .A1(net4460),
    .A2(net1902));
 sg13g2_a21oi_1 _15716_ (.A1(_01772_),
    .A2(net1902),
    .Y(_01310_),
    .B1(_07076_));
 sg13g2_a21oi_1 _15717_ (.A1(net5093),
    .A2(_05371_),
    .Y(_07077_),
    .B1(net1903));
 sg13g2_nor2_1 _15718_ (.A(net2413),
    .B(net5094),
    .Y(_01311_));
 sg13g2_a21oi_1 _15719_ (.A1(_02024_),
    .A2(_06896_),
    .Y(_01312_),
    .B1(net2412));
 sg13g2_nand2_2 _15720_ (.Y(_07078_),
    .A(net4271),
    .B(_06896_));
 sg13g2_o21ai_1 _15721_ (.B1(net2621),
    .Y(_07079_),
    .A1(net4161),
    .A2(net1863));
 sg13g2_a21oi_1 _15722_ (.A1(_01771_),
    .A2(net1863),
    .Y(_01313_),
    .B1(_07079_));
 sg13g2_o21ai_1 _15723_ (.B1(net2621),
    .Y(_07080_),
    .A1(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[1] ),
    .A2(net1863));
 sg13g2_a21oi_1 _15724_ (.A1(_01770_),
    .A2(net1862),
    .Y(_01314_),
    .B1(_07080_));
 sg13g2_o21ai_1 _15725_ (.B1(net2621),
    .Y(_07081_),
    .A1(net3948),
    .A2(net1862));
 sg13g2_a21oi_1 _15726_ (.A1(_01769_),
    .A2(net1862),
    .Y(_01315_),
    .B1(_07081_));
 sg13g2_o21ai_1 _15727_ (.B1(net2622),
    .Y(_07082_),
    .A1(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[3] ),
    .A2(net1863));
 sg13g2_a21oi_1 _15728_ (.A1(_01768_),
    .A2(net1863),
    .Y(_01316_),
    .B1(_07082_));
 sg13g2_o21ai_1 _15729_ (.B1(net2621),
    .Y(_07083_),
    .A1(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[4] ),
    .A2(net1862));
 sg13g2_a21oi_1 _15730_ (.A1(_01767_),
    .A2(net1862),
    .Y(_01317_),
    .B1(_07083_));
 sg13g2_o21ai_1 _15731_ (.B1(net2622),
    .Y(_07084_),
    .A1(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[5] ),
    .A2(_07078_));
 sg13g2_a21oi_1 _15732_ (.A1(_01766_),
    .A2(net1863),
    .Y(_01318_),
    .B1(_07084_));
 sg13g2_o21ai_1 _15733_ (.B1(net2621),
    .Y(_07085_),
    .A1(net4057),
    .A2(net1863));
 sg13g2_a21oi_1 _15734_ (.A1(_01765_),
    .A2(net1862),
    .Y(_01319_),
    .B1(_07085_));
 sg13g2_o21ai_1 _15735_ (.B1(net2621),
    .Y(_07086_),
    .A1(net3831),
    .A2(net1862));
 sg13g2_a21oi_1 _15736_ (.A1(_01764_),
    .A2(net1862),
    .Y(_01320_),
    .B1(_07086_));
 sg13g2_o21ai_1 _15737_ (.B1(_07031_),
    .Y(_07087_),
    .A1(\data_to_write[12] ),
    .A2(_04311_));
 sg13g2_a21oi_1 _15738_ (.A1(\i2c_data_out[8] ),
    .A2(_07087_),
    .Y(_07088_),
    .B1(net4289));
 sg13g2_nor2_1 _15739_ (.A(net2414),
    .B(net4290),
    .Y(_01321_));
 sg13g2_nor2_1 _15740_ (.A(net2559),
    .B(net2340),
    .Y(_07089_));
 sg13g2_nor2_1 _15741_ (.A(net3958),
    .B(_03463_),
    .Y(_07090_));
 sg13g2_nor3_1 _15742_ (.A(_06792_),
    .B(_07089_),
    .C(_07090_),
    .Y(_07091_));
 sg13g2_a21oi_1 _15743_ (.A1(\crc16_read[1] ),
    .A2(net2305),
    .Y(_07092_),
    .B1(_07091_));
 sg13g2_a21oi_1 _15744_ (.A1(net4832),
    .A2(_07092_),
    .Y(_07093_),
    .B1(net1957));
 sg13g2_o21ai_1 _15745_ (.B1(_07093_),
    .Y(_01322_),
    .A1(net4832),
    .A2(_07092_));
 sg13g2_nand2_1 _15746_ (.Y(_07094_),
    .A(net4191),
    .B(net2338));
 sg13g2_o21ai_1 _15747_ (.B1(_07094_),
    .Y(_07095_),
    .A1(net2452),
    .A2(net2340));
 sg13g2_nand2_1 _15748_ (.Y(_07096_),
    .A(net1923),
    .B(_07095_));
 sg13g2_xnor2_1 _15749_ (.Y(_07097_),
    .A(_01762_),
    .B(_07096_));
 sg13g2_a21oi_1 _15750_ (.A1(net4874),
    .A2(net2304),
    .Y(_07098_),
    .B1(net1956));
 sg13g2_o21ai_1 _15751_ (.B1(_07098_),
    .Y(_01323_),
    .A1(net2304),
    .A2(_07097_));
 sg13g2_nand2_1 _15752_ (.Y(_07099_),
    .A(net4303),
    .B(net2338));
 sg13g2_o21ai_1 _15753_ (.B1(_07099_),
    .Y(_07100_),
    .A1(_01777_),
    .A2(net2339));
 sg13g2_nand2_1 _15754_ (.Y(_07101_),
    .A(net1923),
    .B(_07100_));
 sg13g2_xnor2_1 _15755_ (.Y(_07102_),
    .A(_01761_),
    .B(_07101_));
 sg13g2_a21oi_1 _15756_ (.A1(net4964),
    .A2(net2305),
    .Y(_07103_),
    .B1(net1957));
 sg13g2_o21ai_1 _15757_ (.B1(_07103_),
    .Y(_01324_),
    .A1(net2304),
    .A2(_07102_));
 sg13g2_nand2_1 _15758_ (.Y(_07104_),
    .A(net4140),
    .B(net2338));
 sg13g2_o21ai_1 _15759_ (.B1(_07104_),
    .Y(_07105_),
    .A1(net2453),
    .A2(net2340));
 sg13g2_nand2_1 _15760_ (.Y(_07106_),
    .A(net1923),
    .B(_07105_));
 sg13g2_xnor2_1 _15761_ (.Y(_07107_),
    .A(_01760_),
    .B(_07106_));
 sg13g2_a21oi_1 _15762_ (.A1(net4719),
    .A2(net2304),
    .Y(_07108_),
    .B1(net1957));
 sg13g2_o21ai_1 _15763_ (.B1(_07108_),
    .Y(_01325_),
    .A1(net2304),
    .A2(_07107_));
 sg13g2_nand2_1 _15764_ (.Y(_07109_),
    .A(net4213),
    .B(net2338));
 sg13g2_o21ai_1 _15765_ (.B1(_07109_),
    .Y(_07110_),
    .A1(_01775_),
    .A2(net2339));
 sg13g2_nand3_1 _15766_ (.B(net1923),
    .C(_07110_),
    .A(net4719),
    .Y(_07111_));
 sg13g2_a21oi_1 _15767_ (.A1(_06791_),
    .A2(_07110_),
    .Y(_07112_),
    .B1(net4719));
 sg13g2_nand2_1 _15768_ (.Y(_07113_),
    .A(net2308),
    .B(_07111_));
 sg13g2_a21oi_1 _15769_ (.A1(net5013),
    .A2(net2304),
    .Y(_07114_),
    .B1(net1957));
 sg13g2_o21ai_1 _15770_ (.B1(_07114_),
    .Y(_01326_),
    .A1(_07112_),
    .A2(_07113_));
 sg13g2_nand2_1 _15771_ (.Y(_07115_),
    .A(net4243),
    .B(net2339));
 sg13g2_o21ai_1 _15772_ (.B1(_07115_),
    .Y(_07116_),
    .A1(_01774_),
    .A2(net2340));
 sg13g2_nand2_1 _15773_ (.Y(_07117_),
    .A(net1923),
    .B(_07116_));
 sg13g2_xnor2_1 _15774_ (.Y(_07118_),
    .A(_01758_),
    .B(_07117_));
 sg13g2_a21oi_1 _15775_ (.A1(net4992),
    .A2(net2304),
    .Y(_07119_),
    .B1(net1956));
 sg13g2_o21ai_1 _15776_ (.B1(_07119_),
    .Y(_01327_),
    .A1(net2304),
    .A2(_07118_));
 sg13g2_nand2_1 _15777_ (.Y(_07120_),
    .A(net4907),
    .B(net2338));
 sg13g2_o21ai_1 _15778_ (.B1(_07120_),
    .Y(_07121_),
    .A1(_01773_),
    .A2(net2338));
 sg13g2_nand2_1 _15779_ (.Y(_07122_),
    .A(net1923),
    .B(_07121_));
 sg13g2_xnor2_1 _15780_ (.Y(_07123_),
    .A(_01757_),
    .B(_07122_));
 sg13g2_a21oi_1 _15781_ (.A1(net4990),
    .A2(net2306),
    .Y(_07124_),
    .B1(net1956));
 sg13g2_o21ai_1 _15782_ (.B1(_07124_),
    .Y(_01328_),
    .A1(net2306),
    .A2(_07123_));
 sg13g2_nand2_1 _15783_ (.Y(_07125_),
    .A(net3968),
    .B(net2338));
 sg13g2_o21ai_1 _15784_ (.B1(_07125_),
    .Y(_07126_),
    .A1(_01772_),
    .A2(net2338));
 sg13g2_nand2_1 _15785_ (.Y(_07127_),
    .A(net1923),
    .B(_07126_));
 sg13g2_xnor2_1 _15786_ (.Y(_07128_),
    .A(_01756_),
    .B(_07127_));
 sg13g2_a21oi_1 _15787_ (.A1(net4943),
    .A2(net2306),
    .Y(_07129_),
    .B1(net1956));
 sg13g2_o21ai_1 _15788_ (.B1(_07129_),
    .Y(_01329_),
    .A1(net2306),
    .A2(_07128_));
 sg13g2_nand4_1 _15789_ (.B(net2326),
    .C(_03447_),
    .A(_01754_),
    .Y(_07130_),
    .D(net2076));
 sg13g2_nor2_1 _15790_ (.A(net2559),
    .B(net1996),
    .Y(_07131_));
 sg13g2_nor2_1 _15791_ (.A(net3906),
    .B(\i_uart_tx.cycle_counter[1] ),
    .Y(_07132_));
 sg13g2_nand2_1 _15792_ (.Y(_07133_),
    .A(net4354),
    .B(_07132_));
 sg13g2_nand2_1 _15793_ (.Y(_07134_),
    .A(net3995),
    .B(net4466));
 sg13g2_nand2_1 _15794_ (.Y(_07135_),
    .A(net4646),
    .B(net4675));
 sg13g2_nor4_1 _15795_ (.A(net4606),
    .B(net4691),
    .C(_07134_),
    .D(_07135_),
    .Y(_07136_));
 sg13g2_nand2b_2 _15796_ (.Y(_07137_),
    .B(_07136_),
    .A_N(_07133_));
 sg13g2_nor2b_1 _15797_ (.A(net4606),
    .B_N(net4675),
    .Y(_07138_));
 sg13g2_nor4_1 _15798_ (.A(net4691),
    .B(_01755_),
    .C(_07133_),
    .D(_07134_),
    .Y(_07139_));
 sg13g2_nand4_1 _15799_ (.B(_06223_),
    .C(_07138_),
    .A(_03448_),
    .Y(_07140_),
    .D(_07139_));
 sg13g2_mux2_1 _15800_ (.A0(net5295),
    .A1(net4940),
    .S(_07140_),
    .X(_07141_));
 sg13g2_nor2b_1 _15801_ (.A(_07141_),
    .B_N(net1996),
    .Y(_07142_));
 sg13g2_nor3_1 _15802_ (.A(net2415),
    .B(_07131_),
    .C(_07142_),
    .Y(_01330_));
 sg13g2_nor2_1 _15803_ (.A(net2557),
    .B(net1996),
    .Y(_07143_));
 sg13g2_mux2_1 _15804_ (.A0(net5305),
    .A1(net5295),
    .S(_07140_),
    .X(_07144_));
 sg13g2_nor2b_1 _15805_ (.A(_07144_),
    .B_N(net1995),
    .Y(_07145_));
 sg13g2_nor3_1 _15806_ (.A(net2415),
    .B(_07143_),
    .C(_07145_),
    .Y(_01331_));
 sg13g2_nor2_1 _15807_ (.A(net2556),
    .B(net1995),
    .Y(_07146_));
 sg13g2_mux2_1 _15808_ (.A0(net5301),
    .A1(\i_uart_tx.data_to_send[2] ),
    .S(_07140_),
    .X(_07147_));
 sg13g2_nor2b_1 _15809_ (.A(net5302),
    .B_N(net1995),
    .Y(_07148_));
 sg13g2_nor3_1 _15810_ (.A(net2415),
    .B(_07146_),
    .C(_07148_),
    .Y(_01332_));
 sg13g2_nor2_1 _15811_ (.A(net4848),
    .B(net1994),
    .Y(_07149_));
 sg13g2_mux2_1 _15812_ (.A0(\i_uart_tx.data_to_send[4] ),
    .A1(\i_uart_tx.data_to_send[3] ),
    .S(_07140_),
    .X(_07150_));
 sg13g2_nor2b_1 _15813_ (.A(_07150_),
    .B_N(net1994),
    .Y(_07151_));
 sg13g2_nor3_1 _15814_ (.A(net2416),
    .B(_07149_),
    .C(_07151_),
    .Y(_01333_));
 sg13g2_nor2_1 _15815_ (.A(net4793),
    .B(net1994),
    .Y(_07152_));
 sg13g2_mux2_1 _15816_ (.A0(\i_uart_tx.data_to_send[5] ),
    .A1(\i_uart_tx.data_to_send[4] ),
    .S(_07140_),
    .X(_07153_));
 sg13g2_nor2b_1 _15817_ (.A(_07153_),
    .B_N(net1994),
    .Y(_07154_));
 sg13g2_nor3_1 _15818_ (.A(net2416),
    .B(_07152_),
    .C(_07154_),
    .Y(_01334_));
 sg13g2_nor2_1 _15819_ (.A(net4814),
    .B(net1994),
    .Y(_07155_));
 sg13g2_mux2_1 _15820_ (.A0(\i_uart_tx.data_to_send[6] ),
    .A1(\i_uart_tx.data_to_send[5] ),
    .S(_07140_),
    .X(_07156_));
 sg13g2_nor2b_1 _15821_ (.A(_07156_),
    .B_N(net1995),
    .Y(_07157_));
 sg13g2_nor3_1 _15822_ (.A(net2416),
    .B(_07155_),
    .C(_07157_),
    .Y(_01335_));
 sg13g2_nor2_1 _15823_ (.A(net4708),
    .B(net1994),
    .Y(_07158_));
 sg13g2_mux2_1 _15824_ (.A0(net3591),
    .A1(\i_uart_tx.data_to_send[6] ),
    .S(_07140_),
    .X(_07159_));
 sg13g2_nor2b_1 _15825_ (.A(_07159_),
    .B_N(net1995),
    .Y(_07160_));
 sg13g2_nor3_1 _15826_ (.A(net2416),
    .B(_07158_),
    .C(_07160_),
    .Y(_01336_));
 sg13g2_nand4_1 _15827_ (.B(net2637),
    .C(net1994),
    .A(net3591),
    .Y(_07161_),
    .D(_07140_));
 sg13g2_o21ai_1 _15828_ (.B1(_07161_),
    .Y(_01337_),
    .A1(_04444_),
    .A2(net1994));
 sg13g2_nand2_1 _15829_ (.Y(_07162_),
    .A(net2632),
    .B(_07137_));
 sg13g2_nor2_1 _15830_ (.A(net4354),
    .B(_03449_),
    .Y(_07163_));
 sg13g2_and2_1 _15831_ (.A(net4354),
    .B(_03449_),
    .X(_07164_));
 sg13g2_nor3_1 _15832_ (.A(net2143),
    .B(net4355),
    .C(_07164_),
    .Y(_01338_));
 sg13g2_a21oi_1 _15833_ (.A1(net4891),
    .A2(_07164_),
    .Y(_07165_),
    .B1(net2142));
 sg13g2_o21ai_1 _15834_ (.B1(_07165_),
    .Y(_07166_),
    .A1(net4891),
    .A2(_07164_));
 sg13g2_inv_1 _15835_ (.Y(_01339_),
    .A(_07166_));
 sg13g2_a21oi_1 _15836_ (.A1(\i_uart_tx.cycle_counter[1] ),
    .A2(_07164_),
    .Y(_07167_),
    .B1(net3906));
 sg13g2_and3_1 _15837_ (.X(_07168_),
    .A(net3906),
    .B(\i_uart_tx.cycle_counter[1] ),
    .C(_07164_));
 sg13g2_nor3_1 _15838_ (.A(net2142),
    .B(net3907),
    .C(_07168_),
    .Y(_01340_));
 sg13g2_nor2_1 _15839_ (.A(net4675),
    .B(_07168_),
    .Y(_07169_));
 sg13g2_and2_1 _15840_ (.A(net4675),
    .B(_07168_),
    .X(_07170_));
 sg13g2_nor3_1 _15841_ (.A(net2142),
    .B(net4676),
    .C(_07170_),
    .Y(_01341_));
 sg13g2_nor2_1 _15842_ (.A(net4646),
    .B(_07170_),
    .Y(_07171_));
 sg13g2_and2_1 _15843_ (.A(net4646),
    .B(_07170_),
    .X(_07172_));
 sg13g2_nor3_1 _15844_ (.A(net2142),
    .B(net4647),
    .C(_07172_),
    .Y(_01342_));
 sg13g2_nor2_1 _15845_ (.A(net4691),
    .B(_07172_),
    .Y(_07173_));
 sg13g2_and2_1 _15846_ (.A(net4691),
    .B(_07172_),
    .X(_07174_));
 sg13g2_nor3_1 _15847_ (.A(net2142),
    .B(_07173_),
    .C(_07174_),
    .Y(_01343_));
 sg13g2_nor2_1 _15848_ (.A(net4466),
    .B(_07174_),
    .Y(_07175_));
 sg13g2_and2_1 _15849_ (.A(net4466),
    .B(_07174_),
    .X(_07176_));
 sg13g2_nor3_1 _15850_ (.A(net2142),
    .B(net4467),
    .C(_07176_),
    .Y(_01344_));
 sg13g2_nor2_1 _15851_ (.A(net3995),
    .B(_07176_),
    .Y(_07177_));
 sg13g2_nor2b_1 _15852_ (.A(_07134_),
    .B_N(_07174_),
    .Y(_07178_));
 sg13g2_nor3_1 _15853_ (.A(net2142),
    .B(net3996),
    .C(_07178_),
    .Y(_01345_));
 sg13g2_xnor2_1 _15854_ (.Y(_07179_),
    .A(net4606),
    .B(_07178_));
 sg13g2_nor2_1 _15855_ (.A(net2142),
    .B(net4607),
    .Y(_01346_));
 sg13g2_and4_1 _15856_ (.A(net4715),
    .B(_01753_),
    .C(\i_uart_tx.fsm_state[1] ),
    .D(_01754_),
    .X(_07180_));
 sg13g2_inv_1 _15857_ (.Y(_07181_),
    .A(_07180_));
 sg13g2_nor4_1 _15858_ (.A(net5040),
    .B(_03447_),
    .C(_07137_),
    .D(_07180_),
    .Y(_07182_));
 sg13g2_a21oi_1 _15859_ (.A1(net5040),
    .A2(_07137_),
    .Y(_07183_),
    .B1(_07182_));
 sg13g2_a21oi_1 _15860_ (.A1(net1996),
    .A2(net5041),
    .Y(_01347_),
    .B1(net2414));
 sg13g2_nand2_1 _15861_ (.Y(_07184_),
    .A(_03449_),
    .B(_07137_));
 sg13g2_a22oi_1 _15862_ (.Y(_07185_),
    .B1(_07181_),
    .B2(_01754_),
    .A2(_07137_),
    .A1(_03449_));
 sg13g2_o21ai_1 _15863_ (.B1(net2632),
    .Y(_07186_),
    .A1(net4021),
    .A2(_07185_));
 sg13g2_a21oi_1 _15864_ (.A1(net4021),
    .A2(_07185_),
    .Y(_01348_),
    .B1(_07186_));
 sg13g2_nand4_1 _15865_ (.B(\i_uart_tx.fsm_state[0] ),
    .C(_07138_),
    .A(net4021),
    .Y(_07187_),
    .D(_07139_));
 sg13g2_nand3_1 _15866_ (.B(net4021),
    .C(\i_uart_tx.fsm_state[0] ),
    .A(net4762),
    .Y(_07188_));
 sg13g2_nand2_1 _15867_ (.Y(_07189_),
    .A(net2632),
    .B(_07188_));
 sg13g2_a22oi_1 _15868_ (.Y(_01349_),
    .B1(_07189_),
    .B2(net2143),
    .A2(_07187_),
    .A1(_01753_));
 sg13g2_xnor2_1 _15869_ (.Y(_07190_),
    .A(net4715),
    .B(_07188_));
 sg13g2_nand4_1 _15870_ (.B(_07181_),
    .C(_07184_),
    .A(net2632),
    .Y(_07191_),
    .D(_07190_));
 sg13g2_o21ai_1 _15871_ (.B1(_07191_),
    .Y(_01350_),
    .A1(_01752_),
    .A2(net2143));
 sg13g2_nand3b_1 _15872_ (.B(net3818),
    .C(net3811),
    .Y(_07192_),
    .A_N(net4713));
 sg13g2_nor2_1 _15873_ (.A(\i_uart_rx.cycle_counter[2] ),
    .B(net4820),
    .Y(_07193_));
 sg13g2_nand3_1 _15874_ (.B(net4764),
    .C(_07193_),
    .A(net4539),
    .Y(_07194_));
 sg13g2_nor4_2 _15875_ (.A(_01988_),
    .B(net4953),
    .C(_07192_),
    .Y(_07195_),
    .D(_07194_));
 sg13g2_or3_1 _15876_ (.A(\i_uart_rx.fsm_state[3] ),
    .B(net4787),
    .C(net2459),
    .X(_07196_));
 sg13g2_o21ai_1 _15877_ (.B1(\i_uart_rx.fsm_state[3] ),
    .Y(_07197_),
    .A1(\i_uart_rx.fsm_state[2] ),
    .A2(\i_uart_rx.fsm_state[1] ));
 sg13g2_nand3_1 _15878_ (.B(_07196_),
    .C(_07197_),
    .A(_07195_),
    .Y(_07198_));
 sg13g2_mux2_1 _15879_ (.A0(\i_uart_rx.recieved_data[1] ),
    .A1(net4193),
    .S(_07198_),
    .X(_01351_));
 sg13g2_mux2_1 _15880_ (.A0(net4697),
    .A1(\i_uart_rx.recieved_data[1] ),
    .S(_07198_),
    .X(_01352_));
 sg13g2_mux2_1 _15881_ (.A0(net4699),
    .A1(net4697),
    .S(_07198_),
    .X(_01353_));
 sg13g2_mux2_1 _15882_ (.A0(net4738),
    .A1(net4699),
    .S(_07198_),
    .X(_01354_));
 sg13g2_mux2_1 _15883_ (.A0(net4731),
    .A1(net4738),
    .S(_07198_),
    .X(_01355_));
 sg13g2_mux2_1 _15884_ (.A0(\i_uart_rx.recieved_data[6] ),
    .A1(net4731),
    .S(_07198_),
    .X(_01356_));
 sg13g2_mux2_1 _15885_ (.A0(net4295),
    .A1(net4775),
    .S(_07198_),
    .X(_01357_));
 sg13g2_mux2_1 _15886_ (.A0(net4044),
    .A1(net4295),
    .S(_07198_),
    .X(_01358_));
 sg13g2_nor2_1 _15887_ (.A(\i_uart_rx.fsm_state[0] ),
    .B(_07196_),
    .Y(_07199_));
 sg13g2_nor2_1 _15888_ (.A(_07195_),
    .B(_07199_),
    .Y(_07200_));
 sg13g2_nand3b_1 _15889_ (.B(_07200_),
    .C(net2641),
    .Y(_07201_),
    .A_N(_03671_));
 sg13g2_nor2_1 _15890_ (.A(net3408),
    .B(net2102),
    .Y(_01359_));
 sg13g2_and2_1 _15891_ (.A(net3408),
    .B(net4953),
    .X(_07202_));
 sg13g2_nor2_1 _15892_ (.A(net3408),
    .B(net4953),
    .Y(_07203_));
 sg13g2_nor3_1 _15893_ (.A(net2102),
    .B(_07202_),
    .C(_07203_),
    .Y(_01360_));
 sg13g2_xnor2_1 _15894_ (.Y(_07204_),
    .A(net4821),
    .B(_07202_));
 sg13g2_nor2_1 _15895_ (.A(net2102),
    .B(net4822),
    .Y(_01361_));
 sg13g2_a21oi_1 _15896_ (.A1(\i_uart_rx.cycle_counter[2] ),
    .A2(_07202_),
    .Y(_07205_),
    .B1(net3811));
 sg13g2_and3_1 _15897_ (.X(_07206_),
    .A(\i_uart_rx.cycle_counter[2] ),
    .B(net3811),
    .C(_07202_));
 sg13g2_nor3_1 _15898_ (.A(net2102),
    .B(net3812),
    .C(_07206_),
    .Y(_01362_));
 sg13g2_nor2_1 _15899_ (.A(net4539),
    .B(_07206_),
    .Y(_07207_));
 sg13g2_and2_1 _15900_ (.A(net4539),
    .B(_07206_),
    .X(_07208_));
 sg13g2_nor3_1 _15901_ (.A(net2102),
    .B(net4540),
    .C(_07208_),
    .Y(_01363_));
 sg13g2_xnor2_1 _15902_ (.Y(_07209_),
    .A(net4820),
    .B(_07208_));
 sg13g2_nor2_1 _15903_ (.A(net2102),
    .B(_07209_),
    .Y(_01364_));
 sg13g2_a21oi_1 _15904_ (.A1(\i_uart_rx.cycle_counter[5] ),
    .A2(_07208_),
    .Y(_07210_),
    .B1(net3818));
 sg13g2_and3_1 _15905_ (.X(_07211_),
    .A(net5385),
    .B(net3818),
    .C(_07208_));
 sg13g2_nor3_1 _15906_ (.A(net2102),
    .B(net3819),
    .C(_07211_),
    .Y(_01365_));
 sg13g2_nor2_1 _15907_ (.A(net4764),
    .B(_07211_),
    .Y(_07212_));
 sg13g2_and2_1 _15908_ (.A(net4764),
    .B(_07211_),
    .X(_07213_));
 sg13g2_nor3_1 _15909_ (.A(net2102),
    .B(net4765),
    .C(_07213_),
    .Y(_01366_));
 sg13g2_a21oi_1 _15910_ (.A1(net4713),
    .A2(_07213_),
    .Y(_07214_),
    .B1(_07201_));
 sg13g2_o21ai_1 _15911_ (.B1(_07214_),
    .Y(_07215_),
    .A1(net4713),
    .A2(_07213_));
 sg13g2_inv_1 _15912_ (.Y(_01367_),
    .A(net4714));
 sg13g2_nor2_1 _15913_ (.A(\i_uart_rx.cycle_counter[4] ),
    .B(\i_uart_rx.cycle_counter[7] ),
    .Y(_07216_));
 sg13g2_nand4_1 _15914_ (.B(\i_uart_rx.cycle_counter[5] ),
    .C(_07203_),
    .A(\i_uart_rx.cycle_counter[2] ),
    .Y(_07217_),
    .D(_07216_));
 sg13g2_nor2_1 _15915_ (.A(_07192_),
    .B(_07217_),
    .Y(_07218_));
 sg13g2_nor2_1 _15916_ (.A(net4044),
    .B(_07218_),
    .Y(_07219_));
 sg13g2_and2_1 _15917_ (.A(_01751_),
    .B(_07218_),
    .X(_07220_));
 sg13g2_nor3_1 _15918_ (.A(net2418),
    .B(net4045),
    .C(_07220_),
    .Y(_01368_));
 sg13g2_nand2b_1 _15919_ (.Y(_01369_),
    .B(net2635),
    .A_N(net3407));
 sg13g2_nand2b_2 _15920_ (.Y(_01370_),
    .B(net2634),
    .A_N(net9));
 sg13g2_nor2_1 _15921_ (.A(_03669_),
    .B(_07199_),
    .Y(_07221_));
 sg13g2_nand2_1 _15922_ (.Y(_07222_),
    .A(_03670_),
    .B(_07200_));
 sg13g2_o21ai_1 _15923_ (.B1(_03671_),
    .Y(_07223_),
    .A1(_03469_),
    .A2(_06699_));
 sg13g2_a21oi_1 _15924_ (.A1(_01751_),
    .A2(_07199_),
    .Y(_07224_),
    .B1(_07221_));
 sg13g2_nor2_1 _15925_ (.A(net2460),
    .B(_03670_),
    .Y(_07225_));
 sg13g2_nand3_1 _15926_ (.B(_07218_),
    .C(_07225_),
    .A(\i_uart_rx.rxd_reg[0] ),
    .Y(_07226_));
 sg13g2_nand3_1 _15927_ (.B(_07224_),
    .C(_07226_),
    .A(_07223_),
    .Y(_07227_));
 sg13g2_a22oi_1 _15928_ (.Y(_07228_),
    .B1(_07222_),
    .B2(_07227_),
    .A2(_03670_),
    .A1(net2460));
 sg13g2_and3_1 _15929_ (.X(_07229_),
    .A(net2460),
    .B(_03670_),
    .C(_07195_));
 sg13g2_nor3_1 _15930_ (.A(net2418),
    .B(net5336),
    .C(_07229_),
    .Y(_01371_));
 sg13g2_nand2b_1 _15931_ (.Y(_07230_),
    .B(_07225_),
    .A_N(_07220_));
 sg13g2_nand2_1 _15932_ (.Y(_07231_),
    .A(_07223_),
    .B(_07230_));
 sg13g2_a21oi_1 _15933_ (.A1(net2459),
    .A2(_03668_),
    .Y(_07232_),
    .B1(net2460));
 sg13g2_a21oi_1 _15934_ (.A1(net2459),
    .A2(net2460),
    .Y(_07233_),
    .B1(_07232_));
 sg13g2_o21ai_1 _15935_ (.B1(_07222_),
    .Y(_07234_),
    .A1(_07231_),
    .A2(_07233_));
 sg13g2_nand3_1 _15936_ (.B(_03668_),
    .C(_07200_),
    .A(net2459),
    .Y(_07235_));
 sg13g2_a21oi_1 _15937_ (.A1(_07234_),
    .A2(_07235_),
    .Y(_01372_),
    .B1(net2418));
 sg13g2_nand3_1 _15938_ (.B(net2460),
    .C(_07222_),
    .A(net2459),
    .Y(_07236_));
 sg13g2_nand3_1 _15939_ (.B(\i_uart_rx.fsm_state[1] ),
    .C(net2460),
    .A(net4787),
    .Y(_07237_));
 sg13g2_nand4_1 _15940_ (.B(net2459),
    .C(net2460),
    .A(net4787),
    .Y(_07238_),
    .D(_07195_));
 sg13g2_nand3_1 _15941_ (.B(_07221_),
    .C(_07238_),
    .A(net2641),
    .Y(_07239_));
 sg13g2_a21oi_1 _15942_ (.A1(_01750_),
    .A2(_07236_),
    .Y(_01373_),
    .B1(_07239_));
 sg13g2_xor2_1 _15943_ (.B(_07237_),
    .A(net5236),
    .X(_07240_));
 sg13g2_nand2_1 _15944_ (.Y(_01660_),
    .A(_07195_),
    .B(_07240_));
 sg13g2_a21oi_1 _15945_ (.A1(_07221_),
    .A2(_01660_),
    .Y(_01661_),
    .B1(_07231_));
 sg13g2_nor3_1 _15946_ (.A(net5236),
    .B(_07195_),
    .C(_07199_),
    .Y(_01662_));
 sg13g2_nor3_1 _15947_ (.A(net2418),
    .B(_01661_),
    .C(net5237),
    .Y(_01374_));
 sg13g2_nor4_1 _15948_ (.A(_04730_),
    .B(_04776_),
    .C(_04778_),
    .D(net1795),
    .Y(_01375_));
 sg13g2_nor2_1 _15949_ (.A(net2443),
    .B(net1801),
    .Y(_01663_));
 sg13g2_a22oi_1 _15950_ (.Y(_01376_),
    .B1(_01663_),
    .B2(_02004_),
    .A2(net1801),
    .A1(_02035_));
 sg13g2_a22oi_1 _15951_ (.Y(_01377_),
    .B1(_01663_),
    .B2(_02009_),
    .A2(net1801),
    .A1(_02036_));
 sg13g2_nand2_1 _15952_ (.Y(_01664_),
    .A(net2626),
    .B(_06758_));
 sg13g2_nand2_1 _15953_ (.Y(_01665_),
    .A(net3542),
    .B(_01664_));
 sg13g2_o21ai_1 _15954_ (.B1(_01665_),
    .Y(_01378_),
    .A1(_01797_),
    .A2(_01664_));
 sg13g2_nand2_2 _15955_ (.Y(_01666_),
    .A(net2629),
    .B(_06756_));
 sg13g2_a21o_1 _15956_ (.A2(net4740),
    .A1(net2454),
    .B1(_01666_),
    .X(_01667_));
 sg13g2_a21oi_1 _15957_ (.A1(_01747_),
    .A2(_01749_),
    .Y(_01379_),
    .B1(_01667_));
 sg13g2_and3_2 _15958_ (.X(_01668_),
    .A(net2454),
    .B(net3619),
    .C(net4740));
 sg13g2_a21oi_1 _15959_ (.A1(net2454),
    .A2(\i_spi.clock_count[0] ),
    .Y(_01669_),
    .B1(net3619));
 sg13g2_nor3_1 _15960_ (.A(_01666_),
    .B(_01668_),
    .C(net3620),
    .Y(_01380_));
 sg13g2_nand2_1 _15961_ (.Y(_01670_),
    .A(\i_spi.clock_count[2] ),
    .B(_01668_));
 sg13g2_xnor2_1 _15962_ (.Y(_01671_),
    .A(net4771),
    .B(_01668_));
 sg13g2_nor2_1 _15963_ (.A(_01666_),
    .B(_01671_),
    .Y(_01381_));
 sg13g2_xor2_1 _15964_ (.B(_01670_),
    .A(net4744),
    .X(_01672_));
 sg13g2_nor2_1 _15965_ (.A(_01666_),
    .B(net4745),
    .Y(_01382_));
 sg13g2_nor2_2 _15966_ (.A(net5007),
    .B(_06756_),
    .Y(_01673_));
 sg13g2_o21ai_1 _15967_ (.B1(_01673_),
    .Y(_01674_),
    .A1(net4199),
    .A2(_01979_));
 sg13g2_nand3_1 _15968_ (.B(_06760_),
    .C(_01674_),
    .A(net2629),
    .Y(_01675_));
 sg13g2_nand2_1 _15969_ (.Y(_01676_),
    .A(net2454),
    .B(net4));
 sg13g2_o21ai_1 _15970_ (.B1(_01676_),
    .Y(_01677_),
    .A1(net2454),
    .A2(_01779_));
 sg13g2_mux2_1 _15971_ (.A0(_01677_),
    .A1(net4784),
    .S(_01675_),
    .X(_01383_));
 sg13g2_nand2_1 _15972_ (.Y(_01678_),
    .A(net2626),
    .B(_06759_));
 sg13g2_nor4_2 _15973_ (.A(net4199),
    .B(net4603),
    .C(net4916),
    .Y(_01679_),
    .D(net4229));
 sg13g2_a21oi_1 _15974_ (.A1(net2458),
    .A2(_01679_),
    .Y(_01680_),
    .B1(_06761_));
 sg13g2_nand2_1 _15975_ (.Y(_01681_),
    .A(net4229),
    .B(_06761_));
 sg13g2_nand2b_2 _15976_ (.Y(_01682_),
    .B(_01680_),
    .A_N(net4229));
 sg13g2_a21oi_1 _15977_ (.A1(net4230),
    .A2(_01682_),
    .Y(_01384_),
    .B1(_01678_));
 sg13g2_xor2_1 _15978_ (.B(_01682_),
    .A(net4916),
    .X(_01683_));
 sg13g2_nor2_1 _15979_ (.A(_01678_),
    .B(_01683_),
    .Y(_01385_));
 sg13g2_o21ai_1 _15980_ (.B1(net4603),
    .Y(_01684_),
    .A1(\i_spi.bits_remaining[1] ),
    .A2(_01682_));
 sg13g2_or3_1 _15981_ (.A(net4603),
    .B(\i_spi.bits_remaining[1] ),
    .C(_01682_),
    .X(_01685_));
 sg13g2_a21oi_1 _15982_ (.A1(net4604),
    .A2(_01685_),
    .Y(_01386_),
    .B1(_01678_));
 sg13g2_nand3_1 _15983_ (.B(net2626),
    .C(_01685_),
    .A(net4199),
    .Y(_01686_));
 sg13g2_nand2_1 _15984_ (.Y(_01387_),
    .A(_01664_),
    .B(net4200));
 sg13g2_nand2_1 _15985_ (.Y(_01687_),
    .A(_01673_),
    .B(_01679_));
 sg13g2_a221oi_1 _15986_ (.B2(_01679_),
    .C1(net2413),
    .B1(_01673_),
    .A1(_01747_),
    .Y(_01388_),
    .A2(_06757_));
 sg13g2_nand3_1 _15987_ (.B(_06759_),
    .C(_01687_),
    .A(net4250),
    .Y(_01688_));
 sg13g2_nand4_1 _15988_ (.B(net3542),
    .C(_01673_),
    .A(net2454),
    .Y(_01689_),
    .D(_01679_));
 sg13g2_nand3_1 _15989_ (.B(net4251),
    .C(_01689_),
    .A(net2629),
    .Y(_01389_));
 sg13g2_a21oi_1 _15990_ (.A1(_02075_),
    .A2(_06392_),
    .Y(_01390_),
    .B1(_06408_));
 sg13g2_nand2_1 _15991_ (.Y(_01690_),
    .A(_06760_),
    .B(_01679_));
 sg13g2_o21ai_1 _15992_ (.B1(_01690_),
    .Y(_01691_),
    .A1(net5007),
    .A2(_06760_));
 sg13g2_nor3_1 _15993_ (.A(net2413),
    .B(_06762_),
    .C(_01691_),
    .Y(_01391_));
 sg13g2_o21ai_1 _15994_ (.B1(_06786_),
    .Y(_01692_),
    .A1(net2465),
    .A2(_02755_));
 sg13g2_o21ai_1 _15995_ (.B1(_01692_),
    .Y(_01640_),
    .A1(_02111_),
    .A2(_06787_));
 sg13g2_nand2_1 _15996_ (.Y(_01693_),
    .A(net2619),
    .B(net2332));
 sg13g2_o21ai_1 _15997_ (.B1(net4329),
    .Y(_01694_),
    .A1(_05370_),
    .A2(_05400_));
 sg13g2_nor2_1 _15998_ (.A(_01693_),
    .B(net4330),
    .Y(_01641_));
 sg13g2_a21oi_1 _15999_ (.A1(net2465),
    .A2(_06785_),
    .Y(_01695_),
    .B1(net5024));
 sg13g2_nor2_1 _16000_ (.A(_06789_),
    .B(net5025),
    .Y(_01642_));
 sg13g2_nand3_1 _16001_ (.B(_05394_),
    .C(_06821_),
    .A(_05356_),
    .Y(_01696_));
 sg13g2_o21ai_1 _16002_ (.B1(_05369_),
    .Y(_01697_),
    .A1(net2544),
    .A2(_05366_));
 sg13g2_nand3_1 _16003_ (.B(_01696_),
    .C(_01697_),
    .A(_05881_),
    .Y(_01698_));
 sg13g2_a221oi_1 _16004_ (.B2(\i_i2c_peri.i_i2c.data_reg[6] ),
    .C1(net1922),
    .B1(net2223),
    .A1(\i_i2c_peri.i_i2c.s_axis_data_tdata[7] ),
    .Y(_01699_),
    .A2(_05372_));
 sg13g2_a21oi_1 _16005_ (.A1(_02088_),
    .A2(net1922),
    .Y(_01643_),
    .B1(_01699_));
 sg13g2_a221oi_1 _16006_ (.B2(\i_i2c_peri.i_i2c.data_reg[5] ),
    .C1(net1922),
    .B1(net2222),
    .A1(\i_i2c_peri.i_i2c.s_axis_data_tdata[6] ),
    .Y(_01700_),
    .A2(net2283));
 sg13g2_a21oi_1 _16007_ (.A1(_02033_),
    .A2(net1922),
    .Y(_01644_),
    .B1(_01700_));
 sg13g2_a221oi_1 _16008_ (.B2(net4367),
    .C1(net1921),
    .B1(net2222),
    .A1(\i_i2c_peri.i_i2c.s_axis_data_tdata[5] ),
    .Y(_01701_),
    .A2(net2283));
 sg13g2_a21oi_1 _16009_ (.A1(_02032_),
    .A2(net1922),
    .Y(_01645_),
    .B1(_01701_));
 sg13g2_a221oi_1 _16010_ (.B2(\i_i2c_peri.i_i2c.data_reg[3] ),
    .C1(net1921),
    .B1(net2222),
    .A1(\i_i2c_peri.i_i2c.s_axis_data_tdata[4] ),
    .Y(_01702_),
    .A2(net2283));
 sg13g2_a21oi_1 _16011_ (.A1(_02031_),
    .A2(_01698_),
    .Y(_01646_),
    .B1(_01702_));
 sg13g2_a221oi_1 _16012_ (.B2(\i_i2c_peri.i_i2c.data_reg[2] ),
    .C1(net1921),
    .B1(net2222),
    .A1(\i_i2c_peri.i_i2c.s_axis_data_tdata[3] ),
    .Y(_01703_),
    .A2(net2283));
 sg13g2_a21oi_1 _16013_ (.A1(_02030_),
    .A2(net1922),
    .Y(_01647_),
    .B1(_01703_));
 sg13g2_a221oi_1 _16014_ (.B2(\i_i2c_peri.i_i2c.data_reg[1] ),
    .C1(net1921),
    .B1(net2223),
    .A1(\i_i2c_peri.i_i2c.s_axis_data_tdata[2] ),
    .Y(_01704_),
    .A2(net2283));
 sg13g2_a21oi_1 _16015_ (.A1(_02029_),
    .A2(net1921),
    .Y(_01648_),
    .B1(_01704_));
 sg13g2_a221oi_1 _16016_ (.B2(net4339),
    .C1(net1921),
    .B1(net2223),
    .A1(\i_i2c_peri.i_i2c.s_axis_data_tdata[1] ),
    .Y(_01705_),
    .A2(_05372_));
 sg13g2_a21oi_1 _16017_ (.A1(_02028_),
    .A2(net1921),
    .Y(_01649_),
    .B1(_01705_));
 sg13g2_a221oi_1 _16018_ (.B2(net4329),
    .C1(net1922),
    .B1(net2223),
    .A1(net4470),
    .Y(_01706_),
    .A2(_05372_));
 sg13g2_a21oi_1 _16019_ (.A1(_02027_),
    .A2(net1921),
    .Y(_01650_),
    .B1(net4471));
 sg13g2_a21oi_1 _16020_ (.A1(net4271),
    .A2(_05361_),
    .Y(_01707_),
    .B1(_06800_));
 sg13g2_and3_1 _16021_ (.X(_01651_),
    .A(net2621),
    .B(_05359_),
    .C(_01707_));
 sg13g2_a21oi_1 _16022_ (.A1(_05373_),
    .A2(_05428_),
    .Y(_01652_),
    .B1(_01693_));
 sg13g2_nand3_1 _16023_ (.B(_02534_),
    .C(_02536_),
    .A(net2528),
    .Y(_01708_));
 sg13g2_nor2_1 _16024_ (.A(_03139_),
    .B(_03393_),
    .Y(_01709_));
 sg13g2_o21ai_1 _16025_ (.B1(net2530),
    .Y(_01710_),
    .A1(net2528),
    .A2(_02810_));
 sg13g2_nand2_1 _16026_ (.Y(_01711_),
    .A(_02537_),
    .B(_05904_));
 sg13g2_nand2_1 _16027_ (.Y(_01712_),
    .A(net2530),
    .B(_01711_));
 sg13g2_nand3_1 _16028_ (.B(_01708_),
    .C(_01709_),
    .A(_02708_),
    .Y(_01713_));
 sg13g2_o21ai_1 _16029_ (.B1(_05899_),
    .Y(_01714_),
    .A1(_01712_),
    .A2(_01713_));
 sg13g2_a21oi_1 _16030_ (.A1(_01742_),
    .A2(_01713_),
    .Y(_01653_),
    .B1(_01714_));
 sg13g2_nor3_2 _16031_ (.A(_02549_),
    .B(_03139_),
    .C(_03393_),
    .Y(_01715_));
 sg13g2_and4_1 _16032_ (.A(net2530),
    .B(_01708_),
    .C(_01711_),
    .D(_01715_),
    .X(_01716_));
 sg13g2_a21oi_1 _16033_ (.A1(_01708_),
    .A2(_01715_),
    .Y(_01717_),
    .B1(net3556));
 sg13g2_nor3_1 _16034_ (.A(_05900_),
    .B(_01716_),
    .C(_01717_),
    .Y(_01654_));
 sg13g2_o21ai_1 _16035_ (.B1(_01715_),
    .Y(_01718_),
    .A1(_02626_),
    .A2(_05904_));
 sg13g2_nand2_1 _16036_ (.Y(_01719_),
    .A(net4177),
    .B(_01718_));
 sg13g2_nand3_1 _16037_ (.B(_01710_),
    .C(_01715_),
    .A(_02626_),
    .Y(_01720_));
 sg13g2_a21oi_1 _16038_ (.A1(_01719_),
    .A2(_01720_),
    .Y(_01655_),
    .B1(_05900_));
 sg13g2_or2_1 _16039_ (.X(_01721_),
    .B(_05904_),
    .A(_02667_));
 sg13g2_nand2_1 _16040_ (.Y(_01722_),
    .A(_01715_),
    .B(_01721_));
 sg13g2_nand2_1 _16041_ (.Y(_01723_),
    .A(net4122),
    .B(_01722_));
 sg13g2_nand3_1 _16042_ (.B(_02667_),
    .C(_05926_),
    .A(net2324),
    .Y(_01724_));
 sg13g2_nand4_1 _16043_ (.B(_02667_),
    .C(_05926_),
    .A(net2324),
    .Y(_01725_),
    .D(_01709_));
 sg13g2_a21oi_1 _16044_ (.A1(_01723_),
    .A2(_01725_),
    .Y(_01656_),
    .B1(_05900_));
 sg13g2_or2_1 _16045_ (.X(_01726_),
    .B(_05904_),
    .A(_02703_));
 sg13g2_nand2_1 _16046_ (.Y(_01727_),
    .A(_01715_),
    .B(_01726_));
 sg13g2_and3_1 _16047_ (.X(_01728_),
    .A(net2324),
    .B(_02703_),
    .C(_01710_));
 sg13g2_a22oi_1 _16048_ (.Y(_01729_),
    .B1(_01728_),
    .B2(_01709_),
    .A2(_01727_),
    .A1(net4828));
 sg13g2_nor2_1 _16049_ (.A(_05900_),
    .B(_01729_),
    .Y(_01657_));
 sg13g2_or2_1 _16050_ (.X(_01730_),
    .B(_03139_),
    .A(_02547_));
 sg13g2_o21ai_1 _16051_ (.B1(_02551_),
    .Y(_01731_),
    .A1(_03380_),
    .A2(_01730_));
 sg13g2_o21ai_1 _16052_ (.B1(_01731_),
    .Y(_01732_),
    .A1(_02549_),
    .A2(_01721_));
 sg13g2_nor2b_1 _16053_ (.A(net4205),
    .B_N(net4436),
    .Y(_01733_));
 sg13g2_o21ai_1 _16054_ (.B1(_02549_),
    .Y(_01734_),
    .A1(net4637),
    .A2(_01733_));
 sg13g2_nor2b_1 _16055_ (.A(_01732_),
    .B_N(_01724_),
    .Y(_01735_));
 sg13g2_a221oi_1 _16056_ (.B2(_01735_),
    .C1(_05900_),
    .B1(_01734_),
    .A1(_01741_),
    .Y(_01658_),
    .A2(_01732_));
 sg13g2_o21ai_1 _16057_ (.B1(_01731_),
    .Y(_01736_),
    .A1(_02549_),
    .A2(_01726_));
 sg13g2_a21oi_1 _16058_ (.A1(\dio1_sync[1] ),
    .A2(_02087_),
    .Y(_01737_),
    .B1(net4357));
 sg13g2_nor2_1 _16059_ (.A(net2324),
    .B(_01737_),
    .Y(_01738_));
 sg13g2_nor3_1 _16060_ (.A(_01728_),
    .B(_01736_),
    .C(_01738_),
    .Y(_01739_));
 sg13g2_nor2b_1 _16061_ (.A(net4357),
    .B_N(_01736_),
    .Y(_01740_));
 sg13g2_nor3_1 _16062_ (.A(_05900_),
    .B(_01739_),
    .C(_01740_),
    .Y(_01659_));
 sg13g2_inv_1 _16064__3 (.Y(net2723),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _16065__4 (.Y(net2724),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _16066__5 (.Y(net2725),
    .A(clknet_leaf_0_clk));
 sg13g2_inv_1 _16067__6 (.Y(net2726),
    .A(clknet_leaf_65_clk));
 sg13g2_inv_1 _16068__7 (.Y(net2727),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _16069__8 (.Y(net2728),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _16070__9 (.Y(net2729),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _16071__10 (.Y(net2730),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _16072__11 (.Y(net2731),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _16073__12 (.Y(net2732),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _16074__13 (.Y(net2733),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _16075__14 (.Y(net2734),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _16076__15 (.Y(net2735),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _16077__16 (.Y(net2736),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 _16078__17 (.Y(net2737),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _16079__18 (.Y(net2738),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _16080__19 (.Y(net2739),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _16081__20 (.Y(net2740),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _16082__21 (.Y(net2741),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _16083__22 (.Y(net2742),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 _16084__23 (.Y(net2743),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _16085__24 (.Y(net2744),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _16086__25 (.Y(net2745),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _16087__26 (.Y(net2746),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _16088__27 (.Y(net2747),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _16089__28 (.Y(net2748),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _16090__29 (.Y(net2749),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _16091__30 (.Y(net2750),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _16092__31 (.Y(net2751),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _16093__32 (.Y(net2752),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _16094__33 (.Y(net2753),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _16095__34 (.Y(net2754),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _16096__35 (.Y(net2755),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _16097__36 (.Y(net2756),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _16098__37 (.Y(net2757),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _16099__38 (.Y(net2758),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _16100__39 (.Y(net2759),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _16101__40 (.Y(net2760),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _16102__41 (.Y(net2761),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _16103__42 (.Y(net2762),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _16104__43 (.Y(net2763),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _16105__44 (.Y(net2764),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _16106__45 (.Y(net2765),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _16107__46 (.Y(net2766),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _16108__47 (.Y(net2767),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _16109__48 (.Y(net2768),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _16110__49 (.Y(net2769),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _16111__50 (.Y(net2770),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _16112__51 (.Y(net2771),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _16113__52 (.Y(net2772),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _16114__53 (.Y(net2773),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _16115__54 (.Y(net2774),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _16116__55 (.Y(net2775),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _16117__56 (.Y(net2776),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _16118__57 (.Y(net2777),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _16119__58 (.Y(net2778),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _16120__59 (.Y(net2779),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _16121__60 (.Y(net2780),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _16122__61 (.Y(net2781),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _16123__62 (.Y(net2782),
    .A(clknet_leaf_32_clk));
 sg13g2_inv_1 _16124__63 (.Y(net2783),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _16125__64 (.Y(net2784),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _16126__65 (.Y(net2785),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _16127__66 (.Y(net2786),
    .A(clknet_leaf_28_clk));
 sg13g2_inv_1 _16128__67 (.Y(net2787),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _16129__68 (.Y(net2788),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _16130__69 (.Y(net2789),
    .A(clknet_leaf_29_clk));
 sg13g2_inv_1 _16131__70 (.Y(net2790),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _16132__71 (.Y(net2791),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _16133__72 (.Y(net2792),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _16134__73 (.Y(net2793),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _16135__74 (.Y(net2794),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _16136__75 (.Y(net2795),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _16137__76 (.Y(net2796),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _16138__77 (.Y(net2797),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _16139__78 (.Y(net2798),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _16140__79 (.Y(net2799),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _16141__80 (.Y(net2800),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 _16142__81 (.Y(net2801),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _16143__82 (.Y(net2802),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _16144__83 (.Y(net2803),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _16145__84 (.Y(net2804),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _16146__85 (.Y(net2805),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _16147__86 (.Y(net2806),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _16148__87 (.Y(net2807),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 _16149__88 (.Y(net2808),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _16150__89 (.Y(net2809),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _16151__90 (.Y(net2810),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _16152__91 (.Y(net2811),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _16153__92 (.Y(net2812),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 _16154__93 (.Y(net2813),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _16155__94 (.Y(net2814),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _16156__95 (.Y(net2815),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _16157__96 (.Y(net2816),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _16158__97 (.Y(net2817),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _16159__98 (.Y(net2818),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _16160__99 (.Y(net2819),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _16161__100 (.Y(net2820),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _16162__101 (.Y(net2821),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _16163__102 (.Y(net2822),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _16164__103 (.Y(net2823),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _16165__104 (.Y(net2824),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _16166__105 (.Y(net2825),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _16167__106 (.Y(net2826),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _16168__107 (.Y(net2827),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _16169__108 (.Y(net2828),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _16170__109 (.Y(net2829),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _16171__110 (.Y(net2830),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _16172__111 (.Y(net2831),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _16173__112 (.Y(net2832),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _16174__113 (.Y(net2833),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _16175__114 (.Y(net2834),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _16176__115 (.Y(net2835),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _16177__116 (.Y(net2836),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _16178__117 (.Y(net2837),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _16179__118 (.Y(net2838),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _16180__119 (.Y(net2839),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _16181__120 (.Y(net2840),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _16182__121 (.Y(net2841),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _16183__122 (.Y(net2842),
    .A(clknet_leaf_18_clk));
 sg13g2_inv_1 _16184__123 (.Y(net2843),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _16185__124 (.Y(net2844),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _16186__125 (.Y(net2845),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _16187__126 (.Y(net2846),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _16188__127 (.Y(net2847),
    .A(clknet_leaf_4_clk));
 sg13g2_inv_1 _16189__128 (.Y(net2848),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 _16190__129 (.Y(net2849),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 _16191__130 (.Y(net2850),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _16192__131 (.Y(net2851),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 _16193__132 (.Y(net2852),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 _16194__133 (.Y(net2853),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _16195__134 (.Y(net2854),
    .A(clknet_leaf_19_clk));
 sg13g2_inv_1 _16196__135 (.Y(net2855),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 _16197__136 (.Y(net2856),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _16198__137 (.Y(net2857),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _16199__138 (.Y(net2858),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _16200__139 (.Y(net2859),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _16201__140 (.Y(net2860),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _16202__141 (.Y(net2861),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _16203__142 (.Y(net2862),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _16204__143 (.Y(net2863),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _16205__144 (.Y(net2864),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _16206__145 (.Y(net2865),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _16207__146 (.Y(net2866),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 _16208__147 (.Y(net2867),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _16209__148 (.Y(net2868),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _16210__149 (.Y(net2869),
    .A(clknet_leaf_45_clk));
 sg13g2_inv_1 _16211__150 (.Y(net2870),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 _16212__151 (.Y(net2871),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _16213__152 (.Y(net2872),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _16214__153 (.Y(net2873),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _16215__154 (.Y(net2874),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _16216__155 (.Y(net2875),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _16217__156 (.Y(net2876),
    .A(clknet_leaf_54_clk));
 sg13g2_inv_1 _16218__157 (.Y(net2877),
    .A(clknet_leaf_57_clk));
 sg13g2_inv_1 _16219__158 (.Y(net2878),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 _16220__159 (.Y(net2879),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _16221__160 (.Y(net2880),
    .A(clknet_leaf_58_clk));
 sg13g2_inv_1 _16222__161 (.Y(net2881),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _16223__162 (.Y(net2882),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _16224__163 (.Y(net2883),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _16225__164 (.Y(net2884),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _16226__165 (.Y(net2885),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _16227__166 (.Y(net2886),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _16228__167 (.Y(net2887),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 _16229__168 (.Y(net2888),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _16230__169 (.Y(net2889),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _16231__170 (.Y(net2890),
    .A(clknet_leaf_12_clk));
 sg13g2_inv_1 _16232__171 (.Y(net2891),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _16233__172 (.Y(net2892),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _16234__173 (.Y(net2893),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _16235__174 (.Y(net2894),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _16236__175 (.Y(net2895),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _16237__176 (.Y(net2896),
    .A(clknet_leaf_35_clk));
 sg13g2_inv_1 _16238__177 (.Y(net2897),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _16239__178 (.Y(net2898),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _16240__179 (.Y(net2899),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _16241__180 (.Y(net2900),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _16242__181 (.Y(net2901),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 _16243__182 (.Y(net2902),
    .A(clknet_leaf_31_clk));
 sg13g2_inv_1 _16244__183 (.Y(net2903),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _16245__184 (.Y(net2904),
    .A(clknet_leaf_26_clk));
 sg13g2_inv_1 _16246__185 (.Y(net2905),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _16247__186 (.Y(net2906),
    .A(clknet_leaf_20_clk));
 sg13g2_inv_1 _16248__187 (.Y(net2907),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _16249__188 (.Y(net2908),
    .A(clknet_leaf_25_clk));
 sg13g2_inv_1 _16250__189 (.Y(net2909),
    .A(clknet_leaf_24_clk));
 sg13g2_inv_1 _16251__190 (.Y(net2910),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _16252__191 (.Y(net2911),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _16253__192 (.Y(net2912),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 _16254__193 (.Y(net2913),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _16255__194 (.Y(net2914),
    .A(clknet_leaf_27_clk));
 sg13g2_inv_1 _16256__195 (.Y(net2915),
    .A(clknet_leaf_33_clk));
 sg13g2_inv_1 _16257__196 (.Y(net2916),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 _16258__197 (.Y(net2917),
    .A(clknet_leaf_34_clk));
 sg13g2_inv_1 _16259__198 (.Y(net2918),
    .A(clknet_leaf_30_clk));
 sg13g2_inv_1 _16260__199 (.Y(net2919),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 _16261__200 (.Y(net2920),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _16262__201 (.Y(net2921),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 _16263__202 (.Y(net2922),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _16264__203 (.Y(net2923),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _16265__204 (.Y(net2924),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _16266__205 (.Y(net2925),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 _16267__206 (.Y(net2926),
    .A(clknet_leaf_44_clk));
 sg13g2_inv_1 _16268__207 (.Y(net2927),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _16269__208 (.Y(net2928),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _16270__209 (.Y(net2929),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _16271__210 (.Y(net2930),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _16272__211 (.Y(net2931),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _16273__212 (.Y(net2932),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _16274__213 (.Y(net2933),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _16275__214 (.Y(net2934),
    .A(clknet_leaf_21_clk));
 sg13g2_inv_1 _16276__215 (.Y(net2935),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _16277__216 (.Y(net2936),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _16278__217 (.Y(net2937),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _16279__218 (.Y(net2938),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _16280__219 (.Y(net2939),
    .A(clknet_leaf_64_clk));
 sg13g2_inv_1 _16281__220 (.Y(net2940),
    .A(clknet_leaf_60_clk));
 sg13g2_inv_1 _16282__221 (.Y(net2941),
    .A(clknet_leaf_63_clk));
 sg13g2_inv_1 _16283__222 (.Y(net2942),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 _16284__223 (.Y(net2943),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _16285__224 (.Y(net2944),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _16286__225 (.Y(net2945),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _16287__226 (.Y(net2946),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _16288__227 (.Y(net2947),
    .A(clknet_leaf_22_clk));
 sg13g2_inv_1 _16289__228 (.Y(net2948),
    .A(clknet_leaf_59_clk));
 sg13g2_inv_1 _16290__229 (.Y(net2949),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 _16291__230 (.Y(net2950),
    .A(clknet_leaf_23_clk));
 sg13g2_inv_1 _16292__231 (.Y(net2951),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _16293__232 (.Y(net2952),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _16294__233 (.Y(net2953),
    .A(clknet_leaf_8_clk));
 sg13g2_inv_1 _16295__234 (.Y(net2954),
    .A(clknet_leaf_9_clk));
 sg13g2_inv_1 _16296__235 (.Y(net2955),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _16297__236 (.Y(net2956),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _16298__237 (.Y(net2957),
    .A(clknet_leaf_2_clk));
 sg13g2_inv_1 _16299__238 (.Y(net2958),
    .A(clknet_leaf_1_clk));
 sg13g2_inv_1 _16300__239 (.Y(net2959),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _16301__240 (.Y(net2960),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _16302__241 (.Y(net2961),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _16303__242 (.Y(net2962),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _16304__243 (.Y(net2963),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 _16305__244 (.Y(net2964),
    .A(clknet_leaf_55_clk));
 sg13g2_inv_1 _16306__245 (.Y(net2965),
    .A(clknet_leaf_48_clk));
 sg13g2_inv_1 _16307__246 (.Y(net2966),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 _16308__247 (.Y(net2967),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _16309__248 (.Y(net2968),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _16310__249 (.Y(net2969),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _16311__250 (.Y(net2970),
    .A(clknet_leaf_36_clk));
 sg13g2_inv_1 _16312__251 (.Y(net2971),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _16313__252 (.Y(net2972),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 _16314__253 (.Y(net2973),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 _16315__254 (.Y(net2974),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 _16316__255 (.Y(net2975),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _16317__256 (.Y(net2976),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _16318__257 (.Y(net2977),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 _16319__258 (.Y(net2978),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _16320__259 (.Y(net2979),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 _16321__260 (.Y(net2980),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 _16322__261 (.Y(net2981),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 _16323__262 (.Y(net2982),
    .A(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbpq_1 _16324_ (.RESET_B(net90),
    .D(_00361_),
    .Q(\i_tinyqv.cpu.i_core.load_top_bit ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16325_ (.RESET_B(net258),
    .D(_00362_),
    .Q(\gpio_out_sel[0] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _16326_ (.RESET_B(net256),
    .D(_00363_),
    .Q(\gpio_out_sel[1] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _16327_ (.RESET_B(net254),
    .D(net4974),
    .Q(\gpio_out_sel[2] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _16328_ (.RESET_B(net252),
    .D(_00365_),
    .Q(\gpio_out_sel[3] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _16329_ (.RESET_B(net250),
    .D(_00366_),
    .Q(\gpio_out_sel[4] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16330_ (.RESET_B(net248),
    .D(_00367_),
    .Q(\gpio_out_sel[5] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _16331_ (.RESET_B(net246),
    .D(_00368_),
    .Q(\gpio_out_sel[6] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _16332_ (.RESET_B(net244),
    .D(net4827),
    .Q(\gpio_out_sel[7] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _16333_ (.RESET_B(net242),
    .D(net4609),
    .Q(\gpio_out[0] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _16334_ (.RESET_B(net240),
    .D(net3905),
    .Q(\gpio_out[1] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16335_ (.RESET_B(net238),
    .D(net4451),
    .Q(\gpio_out[2] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16336_ (.RESET_B(net236),
    .D(_00373_),
    .Q(\gpio_out[3] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16337_ (.RESET_B(net234),
    .D(net4722),
    .Q(\gpio_out[4] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16338_ (.RESET_B(net232),
    .D(net4457),
    .Q(\gpio_out[5] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _16339_ (.RESET_B(net230),
    .D(net4514),
    .Q(\gpio_out[6] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _16340_ (.RESET_B(net228),
    .D(net4611),
    .Q(\gpio_out[7] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16341_ (.RESET_B(net226),
    .D(net5217),
    .Q(\i_wdt.wdt_reset ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _16342_ (.RESET_B(net225),
    .D(_00379_),
    .Q(\session_ms_div[0] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _16343_ (.RESET_B(net223),
    .D(net3748),
    .Q(\session_ms_div[1] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16344_ (.RESET_B(net221),
    .D(net3417),
    .Q(\session_ms_div[2] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16345_ (.RESET_B(net219),
    .D(net4830),
    .Q(\session_ms_div[3] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16346_ (.RESET_B(net217),
    .D(net3712),
    .Q(\session_ms_div[4] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16347_ (.RESET_B(net215),
    .D(_00384_),
    .Q(\session_ms_div[5] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16348_ (.RESET_B(net213),
    .D(_00385_),
    .Q(\session_ms_div[6] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_2 _16349_ (.RESET_B(net211),
    .D(net3515),
    .Q(\session_ms_div[7] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16350_ (.RESET_B(net209),
    .D(_00387_),
    .Q(\session_ms_div[8] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16351_ (.RESET_B(net207),
    .D(net3415),
    .Q(\session_ms_div[9] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_2 _16352_ (.RESET_B(net205),
    .D(_00389_),
    .Q(\i_seal.session_ctr_in[0] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16353_ (.RESET_B(net203),
    .D(_00390_),
    .Q(\i_seal.session_ctr_in[1] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16354_ (.RESET_B(net201),
    .D(_00391_),
    .Q(\i_seal.session_ctr_in[2] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_2 _16355_ (.RESET_B(net199),
    .D(_00392_),
    .Q(\i_seal.session_ctr_in[3] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16356_ (.RESET_B(net197),
    .D(net3781),
    .Q(\i_seal.session_ctr_in[4] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16357_ (.RESET_B(net195),
    .D(_00394_),
    .Q(\i_seal.session_ctr_in[5] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16358_ (.RESET_B(net193),
    .D(_00395_),
    .Q(\i_seal.session_ctr_in[6] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16359_ (.RESET_B(net191),
    .D(net3991),
    .Q(\i_seal.session_ctr_in[7] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_2 _16360_ (.RESET_B(net189),
    .D(net4694),
    .Q(\pps_count[0] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16361_ (.RESET_B(net187),
    .D(net4043),
    .Q(\pps_count[1] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_2 _16362_ (.RESET_B(net185),
    .D(_00399_),
    .Q(\pps_count[2] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_2 _16363_ (.RESET_B(net183),
    .D(net4855),
    .Q(\pps_count[3] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_2 _16364_ (.RESET_B(net181),
    .D(_00401_),
    .Q(\pps_count[4] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_2 _16365_ (.RESET_B(net179),
    .D(_00402_),
    .Q(\pps_count[5] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16366_ (.RESET_B(net177),
    .D(net4011),
    .Q(\pps_count[6] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16367_ (.RESET_B(net175),
    .D(_00404_),
    .Q(\pps_count[7] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16368_ (.RESET_B(net173),
    .D(net4890),
    .Q(\pps_count[8] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_2 _16369_ (.RESET_B(net171),
    .D(_00406_),
    .Q(\pps_count[9] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16370_ (.RESET_B(net169),
    .D(net4025),
    .Q(\pps_count[10] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16371_ (.RESET_B(net167),
    .D(_00408_),
    .Q(\pps_count[11] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_2 _16372_ (.RESET_B(net165),
    .D(net3571),
    .Q(\pps_count[12] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16373_ (.RESET_B(net163),
    .D(_00410_),
    .Q(\pps_count[13] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16374_ (.RESET_B(net161),
    .D(_00411_),
    .Q(\pps_count[14] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16375_ (.RESET_B(net159),
    .D(net3936),
    .Q(\pps_count[15] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_2 _16376_ (.RESET_B(net157),
    .D(_00413_),
    .Q(\dio1_sync[0] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _16377_ (.RESET_B(net156),
    .D(_00414_),
    .Q(\dio1_sync[1] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16378_ (.RESET_B(net155),
    .D(_00415_),
    .Q(\pps_sync[0] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _16379_ (.RESET_B(net154),
    .D(_00416_),
    .Q(\pps_sync[1] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_2 _16380_ (.RESET_B(net153),
    .D(_00417_),
    .Q(\timer_count[0] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _16381_ (.RESET_B(net151),
    .D(_00418_),
    .Q(\timer_count[1] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _16382_ (.RESET_B(net149),
    .D(_00419_),
    .Q(\timer_count[2] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _16383_ (.RESET_B(net147),
    .D(_00420_),
    .Q(\timer_count[3] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _16384_ (.RESET_B(net145),
    .D(_00421_),
    .Q(\timer_count[4] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _16385_ (.RESET_B(net143),
    .D(_00422_),
    .Q(\timer_count[5] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _16386_ (.RESET_B(net141),
    .D(_00423_),
    .Q(\timer_count[6] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _16387_ (.RESET_B(net139),
    .D(_00424_),
    .Q(\timer_count[7] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _16388_ (.RESET_B(net137),
    .D(_00425_),
    .Q(\timer_count[8] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _16389_ (.RESET_B(net135),
    .D(_00426_),
    .Q(\timer_count[9] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _16390_ (.RESET_B(net133),
    .D(_00427_),
    .Q(\timer_count[10] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _16391_ (.RESET_B(net131),
    .D(net4335),
    .Q(\timer_count[11] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _16392_ (.RESET_B(net129),
    .D(net5155),
    .Q(\timer_count[12] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _16393_ (.RESET_B(net127),
    .D(net5038),
    .Q(\timer_count[13] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _16394_ (.RESET_B(net125),
    .D(_00431_),
    .Q(\timer_count[14] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _16395_ (.RESET_B(net123),
    .D(net4387),
    .Q(\timer_count[15] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _16396_ (.RESET_B(net120),
    .D(_00433_),
    .Q(\timer_count[16] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16397_ (.RESET_B(net118),
    .D(net4915),
    .Q(\timer_count[17] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16398_ (.RESET_B(net116),
    .D(net4757),
    .Q(\timer_count[18] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16399_ (.RESET_B(net114),
    .D(net4913),
    .Q(\timer_count[19] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16400_ (.RESET_B(net112),
    .D(net4801),
    .Q(\timer_count[20] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _16401_ (.RESET_B(net110),
    .D(_00438_),
    .Q(\timer_count[21] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16402_ (.RESET_B(net108),
    .D(net4463),
    .Q(\timer_count[22] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _16403_ (.RESET_B(net106),
    .D(_00440_),
    .Q(\timer_count[23] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _16404_ (.RESET_B(net104),
    .D(_00441_),
    .Q(\timer_count[24] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16405_ (.RESET_B(net102),
    .D(_00442_),
    .Q(\timer_count[25] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16406_ (.RESET_B(net100),
    .D(net4972),
    .Q(\timer_count[26] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_2 _16407_ (.RESET_B(net98),
    .D(_00444_),
    .Q(\timer_count[27] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16408_ (.RESET_B(net96),
    .D(_00445_),
    .Q(\timer_count[28] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16409_ (.RESET_B(net94),
    .D(_00446_),
    .Q(\timer_count[29] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16410_ (.RESET_B(net92),
    .D(_00447_),
    .Q(\timer_count[30] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16411_ (.RESET_B(net89),
    .D(_00448_),
    .Q(\timer_count[31] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16412_ (.RESET_B(net87),
    .D(_00449_),
    .Q(timer_irq),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _16413_ (.RESET_B(net121),
    .D(_00450_),
    .Q(pps_prev),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _16414_ (.RESET_B(net85),
    .D(net3406),
    .Q(\i_crc16.rst_n ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16415_ (.RESET_B(net84),
    .D(net3431),
    .Q(\reset_hold_counter[0] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16416_ (.RESET_B(net82),
    .D(_00452_),
    .Q(\reset_hold_counter[1] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16417_ (.RESET_B(net80),
    .D(_00453_),
    .Q(\reset_hold_counter[2] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16418_ (.RESET_B(net78),
    .D(_00454_),
    .Q(\reset_hold_counter[3] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16419_ (.RESET_B(net76),
    .D(_00455_),
    .Q(\reset_hold_counter[4] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16420_ (.RESET_B(net74),
    .D(_00456_),
    .Q(\i_tinyqv.cpu.i_core.mcause[0] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _16421_ (.RESET_B(net72),
    .D(net4671),
    .Q(\i_tinyqv.cpu.i_core.mcause[1] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _16422_ (.RESET_B(net70),
    .D(net3775),
    .Q(\i_tinyqv.cpu.i_core.mcause[3] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _16423_ (.RESET_B(net68),
    .D(_00459_),
    .Q(\i_tinyqv.cpu.i_core.mcause[4] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _16424_ (.RESET_B(net66),
    .D(net4133),
    .Q(\reset_hold_counter[5] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _16425_ (.RESET_B(net64),
    .D(net4563),
    .Q(\i_tinyqv.cpu.instr_data[1][2] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _16426_ (.RESET_B(net63),
    .D(net4270),
    .Q(\i_tinyqv.cpu.instr_data[1][3] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _16427_ (.RESET_B(net62),
    .D(net4435),
    .Q(\i_tinyqv.cpu.instr_data[1][4] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16428_ (.RESET_B(net61),
    .D(net4465),
    .Q(\i_tinyqv.cpu.instr_data[1][5] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _16429_ (.RESET_B(net60),
    .D(net4615),
    .Q(\i_tinyqv.cpu.instr_data[1][6] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _16430_ (.RESET_B(net59),
    .D(net4419),
    .Q(\i_tinyqv.cpu.instr_data[1][7] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _16431_ (.RESET_B(net58),
    .D(net4164),
    .Q(\i_tinyqv.cpu.instr_data[1][8] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _16432_ (.RESET_B(net57),
    .D(net4595),
    .Q(\i_tinyqv.cpu.instr_data[1][9] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _16433_ (.RESET_B(net56),
    .D(net4485),
    .Q(\i_tinyqv.cpu.instr_data[1][10] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _16434_ (.RESET_B(net55),
    .D(net4593),
    .Q(\i_tinyqv.cpu.instr_data[1][11] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _16435_ (.RESET_B(net54),
    .D(net4522),
    .Q(\i_tinyqv.cpu.instr_data[1][12] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _16436_ (.RESET_B(net53),
    .D(net4476),
    .Q(\i_tinyqv.cpu.instr_data[1][13] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _16437_ (.RESET_B(net52),
    .D(net4517),
    .Q(\i_tinyqv.cpu.instr_data[1][14] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _16438_ (.RESET_B(net51),
    .D(net4483),
    .Q(\i_tinyqv.cpu.instr_data[1][15] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _16439_ (.RESET_B(net50),
    .D(_00475_),
    .Q(\us_divider[0] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_2 _16440_ (.RESET_B(net49),
    .D(_00476_),
    .Q(\us_divider[1] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16441_ (.RESET_B(net48),
    .D(_00477_),
    .Q(\us_divider[2] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16442_ (.RESET_B(net47),
    .D(_00478_),
    .Q(\us_divider[3] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16443_ (.RESET_B(net46),
    .D(_00479_),
    .Q(\us_divider[4] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16444_ (.RESET_B(net297),
    .D(net3653),
    .Q(\i_tinyqv.mem.data_stall ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _16445_ (.RESET_B(net45),
    .D(_00098_),
    .Q(\i_tinyqv.mem.qspi_write_done ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _16446_ (.RESET_B(net43),
    .D(_00481_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _16447_ (.RESET_B(net42),
    .D(_00482_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .CLK(clknet_leaf_195_clk_regs));
 sg13g2_dfrbpq_1 _16448_ (.RESET_B(net41),
    .D(_00483_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _16449_ (.RESET_B(net40),
    .D(_00484_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .CLK(clknet_leaf_195_clk_regs));
 sg13g2_dfrbpq_1 _16450_ (.RESET_B(net39),
    .D(_00485_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _16451_ (.RESET_B(net37),
    .D(_00486_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _16452_ (.RESET_B(net35),
    .D(net4879),
    .Q(\i_tinyqv.cpu.instr_data_in[0] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _16453_ (.RESET_B(net34),
    .D(net4565),
    .Q(\i_tinyqv.cpu.instr_data_in[1] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _16454_ (.RESET_B(net33),
    .D(net5075),
    .Q(\i_tinyqv.cpu.instr_data_in[2] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _16455_ (.RESET_B(net32),
    .D(net4650),
    .Q(\i_tinyqv.cpu.instr_data_in[3] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _16456_ (.RESET_B(net31),
    .D(net5009),
    .Q(\i_tinyqv.cpu.instr_data_in[4] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _16457_ (.RESET_B(net30),
    .D(net5098),
    .Q(\i_tinyqv.cpu.instr_data_in[5] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _16458_ (.RESET_B(net29),
    .D(net5017),
    .Q(\i_tinyqv.cpu.instr_data_in[6] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _16459_ (.RESET_B(net28),
    .D(net5255),
    .Q(\i_tinyqv.cpu.instr_data_in[7] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _16460_ (.RESET_B(net27),
    .D(net3725),
    .Q(\i_tinyqv.mem.qspi_data_buf[8] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16461_ (.RESET_B(net26),
    .D(net4104),
    .Q(\i_tinyqv.mem.qspi_data_buf[9] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _16462_ (.RESET_B(net25),
    .D(net3741),
    .Q(\i_tinyqv.mem.qspi_data_buf[10] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _16463_ (.RESET_B(net24),
    .D(net3824),
    .Q(\i_tinyqv.mem.qspi_data_buf[11] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16464_ (.RESET_B(net23),
    .D(net3849),
    .Q(\i_tinyqv.mem.qspi_data_buf[12] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16465_ (.RESET_B(net22),
    .D(net3879),
    .Q(\i_tinyqv.mem.qspi_data_buf[13] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16466_ (.RESET_B(net21),
    .D(net3981),
    .Q(\i_tinyqv.mem.qspi_data_buf[14] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _16467_ (.RESET_B(net20),
    .D(net3881),
    .Q(\i_tinyqv.mem.qspi_data_buf[15] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _16468_ (.RESET_B(net19),
    .D(net3795),
    .Q(\i_tinyqv.mem.data_from_read[16] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _16469_ (.RESET_B(net18),
    .D(net4176),
    .Q(\i_tinyqv.mem.data_from_read[17] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _16470_ (.RESET_B(net17),
    .D(net4264),
    .Q(\i_tinyqv.mem.data_from_read[18] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _16471_ (.RESET_B(net16),
    .D(net4240),
    .Q(\i_tinyqv.mem.data_from_read[19] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _16472_ (.RESET_B(net15),
    .D(net4097),
    .Q(\i_tinyqv.mem.data_from_read[20] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _16473_ (.RESET_B(net14),
    .D(net4168),
    .Q(\i_tinyqv.mem.data_from_read[21] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _16474_ (.RESET_B(net2720),
    .D(net4196),
    .Q(\i_tinyqv.mem.data_from_read[22] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _16475_ (.RESET_B(net2719),
    .D(net4373),
    .Q(\i_tinyqv.mem.data_from_read[23] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _16476_ (.RESET_B(net2718),
    .D(net3487),
    .Q(\i_tinyqv.mem.qspi_data_buf[24] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16477_ (.RESET_B(net2717),
    .D(net4159),
    .Q(\i_tinyqv.mem.qspi_data_buf[25] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16478_ (.RESET_B(net2716),
    .D(net4146),
    .Q(\i_tinyqv.mem.qspi_data_buf[26] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16479_ (.RESET_B(net2715),
    .D(net4101),
    .Q(\i_tinyqv.mem.qspi_data_buf[27] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _16480_ (.RESET_B(net2714),
    .D(net4089),
    .Q(\i_tinyqv.mem.qspi_data_buf[28] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16481_ (.RESET_B(net2713),
    .D(net4154),
    .Q(\i_tinyqv.mem.qspi_data_buf[29] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _16482_ (.RESET_B(net2712),
    .D(net4131),
    .Q(\i_tinyqv.mem.qspi_data_buf[30] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _16483_ (.RESET_B(net2711),
    .D(net3635),
    .Q(\i_tinyqv.mem.qspi_data_buf[31] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _16484_ (.RESET_B(net2710),
    .D(_00519_),
    .Q(\i_tinyqv.cpu.instr_fetch_started ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _16485_ (.RESET_B(net2709),
    .D(_00520_),
    .Q(\i_tinyqv.mem.instr_active ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _16486_ (.RESET_B(net2707),
    .D(_00521_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16487_ (.RESET_B(net2706),
    .D(_00522_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _16488_ (.RESET_B(net2705),
    .D(_00523_),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _16489_ (.RESET_B(net2704),
    .D(net4911),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _16490_ (.RESET_B(net2703),
    .D(_00525_),
    .Q(\i_tinyqv.mem.q_ctrl.data_req ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _16491_ (.RESET_B(net2702),
    .D(net5034),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _16492_ (.RESET_B(net2700),
    .D(_00527_),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _16493_ (.RESET_B(net2698),
    .D(net4381),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _16494_ (.RESET_B(net2696),
    .D(net4282),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16495_ (.RESET_B(net2694),
    .D(_00530_),
    .Q(\i_tinyqv.mem.q_ctrl.is_writing ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _16496_ (.RESET_B(net2692),
    .D(_00531_),
    .Q(\i_tinyqv.mem.q_ctrl.data_ready ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16497_ (.RESET_B(net2691),
    .D(_00532_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _16498_ (.RESET_B(net2689),
    .D(_00533_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16499_ (.RESET_B(net1773),
    .D(_00534_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16500_ (.RESET_B(net1771),
    .D(_00535_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16501_ (.RESET_B(net1769),
    .D(_00536_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _16502_ (.RESET_B(net1767),
    .D(_00537_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16503_ (.RESET_B(net1765),
    .D(_00538_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _16504_ (.RESET_B(net1763),
    .D(_00539_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_2 _16505_ (.RESET_B(net1761),
    .D(_00540_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _16506_ (.RESET_B(net1759),
    .D(net3721),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16507_ (.RESET_B(net1758),
    .D(net4180),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16508_ (.RESET_B(net1757),
    .D(net4091),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16509_ (.RESET_B(net1756),
    .D(net4126),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _16510_ (.RESET_B(net1755),
    .D(_00545_),
    .Q(\i_tinyqv.cpu.instr_data_in[8] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _16511_ (.RESET_B(net1754),
    .D(_00546_),
    .Q(\i_tinyqv.cpu.instr_data_in[9] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _16512_ (.RESET_B(net1753),
    .D(_00547_),
    .Q(\i_tinyqv.cpu.instr_data_in[10] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _16513_ (.RESET_B(net1752),
    .D(net5273),
    .Q(\i_tinyqv.cpu.instr_data_in[11] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _16514_ (.RESET_B(net1751),
    .D(net5268),
    .Q(\i_tinyqv.cpu.instr_data_in[12] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16515_ (.RESET_B(net1750),
    .D(net5367),
    .Q(\i_tinyqv.cpu.instr_data_in[13] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16516_ (.RESET_B(net1749),
    .D(net5364),
    .Q(\i_tinyqv.cpu.instr_data_in[14] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _16517_ (.RESET_B(net1748),
    .D(net5344),
    .Q(\i_tinyqv.cpu.instr_data_in[15] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _16518_ (.RESET_B(net1747),
    .D(net3562),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _16519_ (.RESET_B(net1746),
    .D(net3745),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _16520_ (.RESET_B(net1745),
    .D(_00555_),
    .Q(\i_tinyqv.cpu.instr_fetch_stopped ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _16521_ (.RESET_B(net1744),
    .D(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_neg ),
    .CLK(net2721));
 sg13g2_dfrbpq_1 _16522_ (.RESET_B(net1743),
    .D(net3680),
    .Q(\i_tinyqv.cpu.instr_data[1][0] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _16523_ (.RESET_B(net1741),
    .D(net3743),
    .Q(\i_tinyqv.cpu.instr_data[1][1] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _16524_ (.RESET_B(net1739),
    .D(_00558_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16525_ (.RESET_B(net1738),
    .D(_00559_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_1 _16526_ (.RESET_B(net1737),
    .D(net4690),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_2 _16527_ (.RESET_B(net1736),
    .D(net4998),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_2 _16528_ (.RESET_B(net1735),
    .D(net4996),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_1 _16529_ (.RESET_B(net1734),
    .D(net4792),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_2 _16530_ (.RESET_B(net1733),
    .D(_00564_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_2 _16531_ (.RESET_B(net1732),
    .D(_00565_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_2 _16532_ (.RESET_B(net1731),
    .D(_00566_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_2 _16533_ (.RESET_B(net1730),
    .D(net5341),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_1 _16534_ (.RESET_B(net1729),
    .D(_00568_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_2 _16535_ (.RESET_B(net1728),
    .D(net5315),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_2 _16536_ (.RESET_B(net1727),
    .D(_00570_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_1 _16537_ (.RESET_B(net1726),
    .D(net4809),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_1 _16538_ (.RESET_B(net1725),
    .D(net4737),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_1 _16539_ (.RESET_B(net1724),
    .D(net4852),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_1 _16540_ (.RESET_B(net1723),
    .D(net4759),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_2 _16541_ (.RESET_B(net1722),
    .D(net4796),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_2 _16542_ (.RESET_B(net1721),
    .D(net4948),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_2 _16543_ (.RESET_B(net1720),
    .D(_00577_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_2 _16544_ (.RESET_B(net1719),
    .D(net4930),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_2 _16545_ (.RESET_B(net1718),
    .D(_00579_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_2 _16546_ (.RESET_B(net1717),
    .D(_00580_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_2 _16547_ (.RESET_B(net1716),
    .D(_00581_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_2 _16548_ (.RESET_B(net1715),
    .D(_00582_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_2 _16549_ (.RESET_B(net1714),
    .D(_00583_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_2 _16550_ (.RESET_B(net1713),
    .D(_00584_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_2 _16551_ (.RESET_B(net1712),
    .D(_00585_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .CLK(clknet_leaf_192_clk_regs));
 sg13g2_dfrbpq_2 _16552_ (.RESET_B(net1711),
    .D(_00586_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_2 _16553_ (.RESET_B(net1710),
    .D(_00587_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_2 _16554_ (.RESET_B(net1709),
    .D(_00588_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_2 _16555_ (.RESET_B(net1708),
    .D(_00589_),
    .Q(\i_tinyqv.cpu.pc[1] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _16556_ (.RESET_B(net1706),
    .D(_00590_),
    .Q(\i_tinyqv.cpu.pc[2] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _16557_ (.RESET_B(net1704),
    .D(_00591_),
    .Q(\i_spi.read_latency ),
    .CLK(net2722));
 sg13g2_dfrbpq_1 _16558_ (.RESET_B(net1702),
    .D(_00592_),
    .Q(\i_spi.clock_divider[0] ),
    .CLK(net2723));
 sg13g2_dfrbpq_1 _16559_ (.RESET_B(net1700),
    .D(_00593_),
    .Q(\i_spi.clock_divider[1] ),
    .CLK(net2724));
 sg13g2_dfrbpq_1 _16560_ (.RESET_B(net1698),
    .D(_00594_),
    .Q(\i_spi.clock_divider[2] ),
    .CLK(net2725));
 sg13g2_dfrbpq_1 _16561_ (.RESET_B(net1696),
    .D(_00595_),
    .Q(\i_spi.clock_divider[3] ),
    .CLK(net2726));
 sg13g2_dfrbpq_1 _16562_ (.RESET_B(net1694),
    .D(_00596_),
    .Q(\i_tinyqv.cpu.instr_data_start[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _16563_ (.RESET_B(net1692),
    .D(_00597_),
    .Q(\i_tinyqv.cpu.instr_data_start[4] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _16564_ (.RESET_B(net1690),
    .D(_00598_),
    .Q(\i_tinyqv.cpu.instr_data_start[5] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _16565_ (.RESET_B(net1688),
    .D(_00599_),
    .Q(\i_tinyqv.cpu.instr_data_start[6] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _16566_ (.RESET_B(net1686),
    .D(_00600_),
    .Q(\i_tinyqv.cpu.instr_data_start[7] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _16567_ (.RESET_B(net1684),
    .D(_00601_),
    .Q(\i_tinyqv.cpu.instr_data_start[8] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _16568_ (.RESET_B(net1682),
    .D(_00602_),
    .Q(\i_tinyqv.cpu.instr_data_start[9] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _16569_ (.RESET_B(net1680),
    .D(_00603_),
    .Q(\i_tinyqv.cpu.instr_data_start[10] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _16570_ (.RESET_B(net1678),
    .D(_00604_),
    .Q(\i_tinyqv.cpu.instr_data_start[11] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _16571_ (.RESET_B(net1676),
    .D(_00605_),
    .Q(\i_tinyqv.cpu.instr_data_start[12] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _16572_ (.RESET_B(net1674),
    .D(_00606_),
    .Q(\i_tinyqv.cpu.instr_data_start[13] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _16573_ (.RESET_B(net1672),
    .D(_00607_),
    .Q(\i_tinyqv.cpu.instr_data_start[14] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _16574_ (.RESET_B(net1670),
    .D(_00608_),
    .Q(\i_tinyqv.cpu.instr_data_start[15] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16575_ (.RESET_B(net1668),
    .D(_00609_),
    .Q(\i_tinyqv.cpu.instr_data_start[16] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _16576_ (.RESET_B(net1666),
    .D(_00610_),
    .Q(\i_tinyqv.cpu.instr_data_start[17] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _16577_ (.RESET_B(net1664),
    .D(_00611_),
    .Q(\i_tinyqv.cpu.instr_data_start[18] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16578_ (.RESET_B(net1662),
    .D(_00612_),
    .Q(\i_tinyqv.cpu.instr_data_start[19] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16579_ (.RESET_B(net1660),
    .D(_00613_),
    .Q(\i_tinyqv.cpu.instr_data_start[20] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16580_ (.RESET_B(net1658),
    .D(_00614_),
    .Q(\i_tinyqv.cpu.instr_data_start[21] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16581_ (.RESET_B(net1656),
    .D(_00615_),
    .Q(\i_tinyqv.cpu.instr_data_start[22] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16582_ (.RESET_B(net1654),
    .D(_00616_),
    .Q(\i_tinyqv.cpu.instr_data_start[23] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16583_ (.RESET_B(net1652),
    .D(_00617_),
    .Q(\i_tinyqv.cpu.instr_fetch_running ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _16584_ (.RESET_B(net1650),
    .D(_00618_),
    .Q(\i_tinyqv.cpu.was_early_branch ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_2 _16585_ (.RESET_B(net1648),
    .D(_00619_),
    .Q(\crc_peri_data[0] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _16586_ (.RESET_B(net1646),
    .D(_00620_),
    .Q(\crc_peri_data[1] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _16587_ (.RESET_B(net1644),
    .D(_00621_),
    .Q(\crc_peri_data[2] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_2 _16588_ (.RESET_B(net1642),
    .D(_00622_),
    .Q(\crc_peri_data[3] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _16589_ (.RESET_B(net1640),
    .D(_00623_),
    .Q(\crc_peri_data[4] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _16590_ (.RESET_B(net1638),
    .D(_00624_),
    .Q(\crc_peri_data[5] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_2 _16591_ (.RESET_B(net1636),
    .D(_00625_),
    .Q(\crc_peri_data[6] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16592_ (.RESET_B(net1634),
    .D(_00626_),
    .Q(\crc_peri_data[7] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _16593_ (.RESET_B(net1632),
    .D(_00627_),
    .Q(\data_to_write[8] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_2 _16594_ (.RESET_B(net1630),
    .D(_00628_),
    .Q(\data_to_write[9] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16595_ (.RESET_B(net1628),
    .D(_00629_),
    .Q(\data_to_write[10] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16596_ (.RESET_B(net1626),
    .D(_00630_),
    .Q(\data_to_write[11] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16597_ (.RESET_B(net1624),
    .D(_00631_),
    .Q(\data_to_write[12] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _16598_ (.RESET_B(net1622),
    .D(_00632_),
    .Q(\data_to_write[13] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _16599_ (.RESET_B(net1620),
    .D(_00633_),
    .Q(\data_to_write[14] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _16600_ (.RESET_B(net1618),
    .D(_00634_),
    .Q(\data_to_write[15] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _16601_ (.RESET_B(net1616),
    .D(_00635_),
    .Q(\data_to_write[16] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _16602_ (.RESET_B(net1614),
    .D(_00636_),
    .Q(\data_to_write[17] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _16603_ (.RESET_B(net1612),
    .D(_00637_),
    .Q(\data_to_write[18] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16604_ (.RESET_B(net1610),
    .D(_00638_),
    .Q(\data_to_write[19] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16605_ (.RESET_B(net1608),
    .D(_00639_),
    .Q(\data_to_write[20] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16606_ (.RESET_B(net1606),
    .D(_00640_),
    .Q(\data_to_write[21] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16607_ (.RESET_B(net1604),
    .D(_00641_),
    .Q(\data_to_write[22] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16608_ (.RESET_B(net1602),
    .D(_00642_),
    .Q(\data_to_write[23] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16609_ (.RESET_B(net1600),
    .D(_00643_),
    .Q(\data_to_write[24] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16610_ (.RESET_B(net1598),
    .D(_00644_),
    .Q(\data_to_write[25] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16611_ (.RESET_B(net1596),
    .D(_00645_),
    .Q(\data_to_write[26] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _16612_ (.RESET_B(net1594),
    .D(_00646_),
    .Q(\data_to_write[27] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16613_ (.RESET_B(net1592),
    .D(_00647_),
    .Q(\data_to_write[28] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _16614_ (.RESET_B(net1590),
    .D(_00648_),
    .Q(\data_to_write[29] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _16615_ (.RESET_B(net1588),
    .D(_00649_),
    .Q(\data_to_write[30] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _16616_ (.RESET_B(net1586),
    .D(_00650_),
    .Q(\data_to_write[31] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _16617_ (.RESET_B(net1584),
    .D(_00651_),
    .Q(\i_tinyqv.cpu.data_write_n[0] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _16618_ (.RESET_B(net1582),
    .D(_00652_),
    .Q(\i_tinyqv.cpu.data_write_n[1] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _16619_ (.RESET_B(net1580),
    .D(net4922),
    .Q(\i_tinyqv.cpu.data_read_n[0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _16620_ (.RESET_B(net375),
    .D(net4950),
    .Q(\i_tinyqv.cpu.data_read_n[1] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _16621_ (.RESET_B(net1578),
    .D(_00044_),
    .Q(debug_data_continue),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _16622_ (.RESET_B(net1576),
    .D(_00655_),
    .Q(\i_tinyqv.cpu.no_write_in_progress ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _16623_ (.RESET_B(net1574),
    .D(net3861),
    .Q(\i_tinyqv.cpu.load_started ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _16624_ (.RESET_B(net1572),
    .D(_00657_),
    .Q(\i_i2c_peri.i_i2c.state_reg[0] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _16625_ (.RESET_B(net1570),
    .D(net4978),
    .Q(\i_i2c_peri.i_i2c.state_reg[1] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _16626_ (.RESET_B(net1568),
    .D(_00659_),
    .Q(\i_i2c_peri.i_i2c.state_reg[2] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _16627_ (.RESET_B(net1566),
    .D(_00660_),
    .Q(\i_i2c_peri.i_i2c.state_reg[3] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _16628_ (.RESET_B(net1564),
    .D(_00661_),
    .Q(\i_tinyqv.cpu.counter[2] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _16629_ (.RESET_B(net1563),
    .D(_00662_),
    .Q(\i_tinyqv.cpu.counter[3] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_2 _16630_ (.RESET_B(net1562),
    .D(_00663_),
    .Q(\i_tinyqv.cpu.counter[4] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _16631_ (.RESET_B(net1561),
    .D(net4310),
    .Q(\i_tinyqv.cpu.data_ready_sync ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _16632_ (.RESET_B(net1559),
    .D(_00665_),
    .Q(\i_tinyqv.cpu.data_ready_latch ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _16633_ (.RESET_B(net1558),
    .D(_00666_),
    .Q(\i_tinyqv.cpu.is_load ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _16634_ (.RESET_B(net1556),
    .D(_00667_),
    .Q(\i_tinyqv.cpu.is_alu_imm ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _16635_ (.RESET_B(net1554),
    .D(_00668_),
    .Q(\i_tinyqv.cpu.is_auipc ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16636_ (.RESET_B(net1552),
    .D(_00669_),
    .Q(\i_tinyqv.cpu.is_store ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _16637_ (.RESET_B(net1550),
    .D(_00670_),
    .Q(\i_tinyqv.cpu.is_alu_reg ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _16638_ (.RESET_B(net1548),
    .D(_00671_),
    .Q(\i_tinyqv.cpu.is_lui ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _16639_ (.RESET_B(net1546),
    .D(_00672_),
    .Q(\i_tinyqv.cpu.is_branch ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _16640_ (.RESET_B(net1544),
    .D(_00673_),
    .Q(\i_tinyqv.cpu.is_jalr ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _16641_ (.RESET_B(net1542),
    .D(net4743),
    .Q(\i_tinyqv.cpu.is_jal ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_2 _16642_ (.RESET_B(net1540),
    .D(_00675_),
    .Q(\i_tinyqv.cpu.is_system ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _16643_ (.RESET_B(net1538),
    .D(_00676_),
    .Q(\i_tinyqv.cpu.instr_len[1] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _16644_ (.RESET_B(net1536),
    .D(_00677_),
    .Q(\i_tinyqv.cpu.instr_len[2] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _16645_ (.RESET_B(net1534),
    .D(_00678_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16646_ (.RESET_B(net1533),
    .D(_00679_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16647_ (.RESET_B(net1532),
    .D(_00680_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16648_ (.RESET_B(net1531),
    .D(_00681_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _16649_ (.RESET_B(net1530),
    .D(_00682_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16650_ (.RESET_B(net1529),
    .D(_00683_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16651_ (.RESET_B(net1528),
    .D(_00684_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _16652_ (.RESET_B(net1527),
    .D(_00685_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16653_ (.RESET_B(net1526),
    .D(_00686_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16654_ (.RESET_B(net1525),
    .D(_00687_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16655_ (.RESET_B(net1524),
    .D(_00688_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _16656_ (.RESET_B(net1523),
    .D(_00689_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16657_ (.RESET_B(net1522),
    .D(_00690_),
    .Q(\i_tinyqv.cpu.imm[12] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16658_ (.RESET_B(net1521),
    .D(_00691_),
    .Q(\i_tinyqv.cpu.imm[13] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16659_ (.RESET_B(net1520),
    .D(_00692_),
    .Q(\i_tinyqv.cpu.imm[14] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16660_ (.RESET_B(net1519),
    .D(_00693_),
    .Q(\i_tinyqv.cpu.imm[15] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16661_ (.RESET_B(net1518),
    .D(_00694_),
    .Q(\i_tinyqv.cpu.imm[16] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16662_ (.RESET_B(net1517),
    .D(_00695_),
    .Q(\i_tinyqv.cpu.imm[17] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16663_ (.RESET_B(net1516),
    .D(_00696_),
    .Q(\i_tinyqv.cpu.imm[18] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16664_ (.RESET_B(net1515),
    .D(_00697_),
    .Q(\i_tinyqv.cpu.imm[19] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16665_ (.RESET_B(net1514),
    .D(_00698_),
    .Q(\i_tinyqv.cpu.imm[20] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16666_ (.RESET_B(net1513),
    .D(_00699_),
    .Q(\i_tinyqv.cpu.imm[21] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16667_ (.RESET_B(net1512),
    .D(_00700_),
    .Q(\i_tinyqv.cpu.imm[22] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16668_ (.RESET_B(net1511),
    .D(_00701_),
    .Q(\i_tinyqv.cpu.imm[23] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16669_ (.RESET_B(net1510),
    .D(_00702_),
    .Q(\i_tinyqv.cpu.imm[24] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16670_ (.RESET_B(net1509),
    .D(_00703_),
    .Q(\i_tinyqv.cpu.imm[25] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16671_ (.RESET_B(net1508),
    .D(_00704_),
    .Q(\i_tinyqv.cpu.imm[26] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16672_ (.RESET_B(net1507),
    .D(_00705_),
    .Q(\i_tinyqv.cpu.imm[27] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _16673_ (.RESET_B(net1506),
    .D(_00706_),
    .Q(\i_tinyqv.cpu.imm[28] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16674_ (.RESET_B(net1505),
    .D(_00707_),
    .Q(\i_tinyqv.cpu.imm[29] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _16675_ (.RESET_B(net1504),
    .D(_00708_),
    .Q(\i_tinyqv.cpu.imm[30] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _16676_ (.RESET_B(net1503),
    .D(_00709_),
    .Q(\i_tinyqv.cpu.imm[31] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16677_ (.RESET_B(net1502),
    .D(_00710_),
    .Q(\i_tinyqv.cpu.alu_op[0] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _16678_ (.RESET_B(net1501),
    .D(_00711_),
    .Q(\i_tinyqv.cpu.alu_op[1] ),
    .CLK(clknet_leaf_195_clk_regs));
 sg13g2_dfrbpq_1 _16679_ (.RESET_B(net1500),
    .D(_00712_),
    .Q(\i_tinyqv.cpu.alu_op[2] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16680_ (.RESET_B(net1499),
    .D(_00713_),
    .Q(\i_tinyqv.cpu.alu_op[3] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16681_ (.RESET_B(net1498),
    .D(_00714_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_2 _16682_ (.RESET_B(net1497),
    .D(_00715_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _16683_ (.RESET_B(net1496),
    .D(_00716_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_2 _16684_ (.RESET_B(net1495),
    .D(_00717_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16685_ (.RESET_B(net1494),
    .D(_00718_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_2 _16686_ (.RESET_B(net1493),
    .D(_00719_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_2 _16687_ (.RESET_B(net1492),
    .D(_00720_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _16688_ (.RESET_B(net1491),
    .D(net3945),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_2 _16689_ (.RESET_B(net1490),
    .D(_00722_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_2 _16690_ (.RESET_B(net1489),
    .D(_00723_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_2 _16691_ (.RESET_B(net1488),
    .D(_00724_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_2 _16692_ (.RESET_B(net1487),
    .D(_00725_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16693_ (.RESET_B(net1485),
    .D(net5051),
    .Q(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _16694_ (.RESET_B(net1483),
    .D(_00727_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16695_ (.RESET_B(net1481),
    .D(_00728_),
    .Q(\i_tinyqv.cpu.mem_op_increment_reg ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_2 _16696_ (.RESET_B(net1479),
    .D(_00729_),
    .Q(\i_tinyqv.cpu.i_core.is_interrupt ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _16697_ (.RESET_B(net1477),
    .D(_00730_),
    .Q(debug_instr_valid),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_2 _16698_ (.RESET_B(net376),
    .D(_00731_),
    .Q(\i_tinyqv.cpu.instr_write_offset[3] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _16699_ (.RESET_B(net377),
    .D(net3288),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_2 _16700_ (.RESET_B(net378),
    .D(net3269),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _16701_ (.RESET_B(net379),
    .D(net3148),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_2 _16702_ (.RESET_B(net380),
    .D(net3347),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _16703_ (.RESET_B(net381),
    .D(net3236),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _16704_ (.RESET_B(net382),
    .D(net3255),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _16705_ (.RESET_B(net383),
    .D(net3281),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _16706_ (.RESET_B(net384),
    .D(net3270),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16707_ (.RESET_B(net385),
    .D(net3283),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _16708_ (.RESET_B(net386),
    .D(net3293),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _16709_ (.RESET_B(net387),
    .D(net3077),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _16710_ (.RESET_B(net388),
    .D(net3116),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16711_ (.RESET_B(net389),
    .D(net2997),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _16712_ (.RESET_B(net390),
    .D(net3096),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _16713_ (.RESET_B(net391),
    .D(net3103),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _16714_ (.RESET_B(net392),
    .D(net3284),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _16715_ (.RESET_B(net393),
    .D(net3314),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _16716_ (.RESET_B(net394),
    .D(net3278),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _16717_ (.RESET_B(net395),
    .D(net3127),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _16718_ (.RESET_B(net396),
    .D(net3100),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _16719_ (.RESET_B(net397),
    .D(net3246),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _16720_ (.RESET_B(net398),
    .D(net3235),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _16721_ (.RESET_B(net399),
    .D(net3368),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _16722_ (.RESET_B(net400),
    .D(net3271),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _16723_ (.RESET_B(net401),
    .D(net3147),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _16724_ (.RESET_B(net402),
    .D(net3136),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .CLK(clknet_leaf_185_clk_regs));
 sg13g2_dfrbpq_1 _16725_ (.RESET_B(net408),
    .D(net3168),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_1 _16726_ (.RESET_B(net1475),
    .D(net3233),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _16727_ (.RESET_B(net1474),
    .D(net5070),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _16728_ (.RESET_B(net1473),
    .D(_00733_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _16729_ (.RESET_B(net1472),
    .D(_00734_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16730_ (.RESET_B(net1471),
    .D(net4399),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16731_ (.RESET_B(net409),
    .D(net4624),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.cy ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_2 _16732_ (.RESET_B(net410),
    .D(net3394),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _16733_ (.RESET_B(net411),
    .D(net3383),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_2 _16734_ (.RESET_B(net412),
    .D(net3393),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_2 _16735_ (.RESET_B(net413),
    .D(net3078),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _16736_ (.RESET_B(net414),
    .D(net3349),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16737_ (.RESET_B(net415),
    .D(net3357),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _16738_ (.RESET_B(net416),
    .D(net3252),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _16739_ (.RESET_B(net417),
    .D(net3360),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _16740_ (.RESET_B(net418),
    .D(net3307),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16741_ (.RESET_B(net419),
    .D(net3185),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _16742_ (.RESET_B(net420),
    .D(net3274),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _16743_ (.RESET_B(net421),
    .D(net3298),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _16744_ (.RESET_B(net422),
    .D(net3007),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16745_ (.RESET_B(net423),
    .D(net3154),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16746_ (.RESET_B(net424),
    .D(net3013),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _16747_ (.RESET_B(net425),
    .D(net2995),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _16748_ (.RESET_B(net426),
    .D(net3207),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16749_ (.RESET_B(net427),
    .D(net2994),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16750_ (.RESET_B(net428),
    .D(net3231),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16751_ (.RESET_B(net429),
    .D(net3247),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _16752_ (.RESET_B(net430),
    .D(net3213),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16753_ (.RESET_B(net431),
    .D(net3050),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _16754_ (.RESET_B(net432),
    .D(net3258),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16755_ (.RESET_B(net433),
    .D(net3114),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _16756_ (.RESET_B(net434),
    .D(net3351),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16757_ (.RESET_B(net435),
    .D(net3220),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_1 _16758_ (.RESET_B(net442),
    .D(net3040),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16759_ (.RESET_B(net1470),
    .D(net3155),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _16760_ (.RESET_B(net1469),
    .D(net4673),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _16761_ (.RESET_B(net1468),
    .D(_00738_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _16762_ (.RESET_B(net1467),
    .D(net5092),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _16763_ (.RESET_B(net1466),
    .D(net5067),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .CLK(clknet_leaf_184_clk_regs));
 sg13g2_dfrbpq_1 _16764_ (.RESET_B(net1465),
    .D(_00741_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_1 _16765_ (.RESET_B(net443),
    .D(_00742_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .CLK(clknet_leaf_182_clk_regs));
 sg13g2_dfrbpq_2 _16766_ (.RESET_B(net444),
    .D(net3183),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_2 _16767_ (.RESET_B(net445),
    .D(net3031),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_2 _16768_ (.RESET_B(net446),
    .D(net3250),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_2 _16769_ (.RESET_B(net447),
    .D(net3107),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16770_ (.RESET_B(net448),
    .D(net3180),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16771_ (.RESET_B(net449),
    .D(net3212),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16772_ (.RESET_B(net450),
    .D(net3311),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16773_ (.RESET_B(net451),
    .D(net3290),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16774_ (.RESET_B(net452),
    .D(net3104),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16775_ (.RESET_B(net453),
    .D(net3170),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16776_ (.RESET_B(net454),
    .D(net3263),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16777_ (.RESET_B(net455),
    .D(net3072),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16778_ (.RESET_B(net456),
    .D(net3365),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16779_ (.RESET_B(net457),
    .D(net3176),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16780_ (.RESET_B(net458),
    .D(net3065),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16781_ (.RESET_B(net459),
    .D(net3184),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16782_ (.RESET_B(net460),
    .D(net3162),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16783_ (.RESET_B(net461),
    .D(net3018),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16784_ (.RESET_B(net462),
    .D(net3097),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16785_ (.RESET_B(net463),
    .D(net3141),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16786_ (.RESET_B(net464),
    .D(net3260),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16787_ (.RESET_B(net465),
    .D(net3122),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16788_ (.RESET_B(net466),
    .D(net3005),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16789_ (.RESET_B(net467),
    .D(net3265),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16790_ (.RESET_B(net468),
    .D(net3068),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16791_ (.RESET_B(net469),
    .D(net3140),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16792_ (.RESET_B(net470),
    .D(net3309),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16793_ (.RESET_B(net471),
    .D(net3029),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16794_ (.RESET_B(net472),
    .D(_00066_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16795_ (.RESET_B(net473),
    .D(_00067_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16796_ (.RESET_B(net474),
    .D(_00068_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16797_ (.RESET_B(net475),
    .D(_00069_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_2 _16798_ (.RESET_B(net476),
    .D(net3124),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_2 _16799_ (.RESET_B(net477),
    .D(net3033),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_2 _16800_ (.RESET_B(net478),
    .D(net3194),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_2 _16801_ (.RESET_B(net479),
    .D(net3102),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16802_ (.RESET_B(net480),
    .D(net3086),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16803_ (.RESET_B(net481),
    .D(net3316),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16804_ (.RESET_B(net482),
    .D(net3313),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16805_ (.RESET_B(net483),
    .D(net3080),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16806_ (.RESET_B(net484),
    .D(net3280),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16807_ (.RESET_B(net485),
    .D(net3081),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16808_ (.RESET_B(net486),
    .D(net3094),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16809_ (.RESET_B(net487),
    .D(net3125),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16810_ (.RESET_B(net488),
    .D(net2987),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16811_ (.RESET_B(net489),
    .D(net3276),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16812_ (.RESET_B(net490),
    .D(net3014),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16813_ (.RESET_B(net491),
    .D(net3156),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16814_ (.RESET_B(net492),
    .D(net3244),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _16815_ (.RESET_B(net493),
    .D(net3164),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16816_ (.RESET_B(net494),
    .D(net3203),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16817_ (.RESET_B(net495),
    .D(net3253),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16818_ (.RESET_B(net496),
    .D(net3024),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _16819_ (.RESET_B(net497),
    .D(net3110),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16820_ (.RESET_B(net498),
    .D(net3279),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16821_ (.RESET_B(net499),
    .D(net3099),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16822_ (.RESET_B(net500),
    .D(net3208),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _16823_ (.RESET_B(net501),
    .D(net3058),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16824_ (.RESET_B(net502),
    .D(net3041),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16825_ (.RESET_B(net503),
    .D(net3083),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16826_ (.RESET_B(net504),
    .D(_00062_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16827_ (.RESET_B(net505),
    .D(_00063_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16828_ (.RESET_B(net506),
    .D(_00064_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16829_ (.RESET_B(net507),
    .D(_00065_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_2 _16830_ (.RESET_B(net508),
    .D(net3322),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_2 _16831_ (.RESET_B(net509),
    .D(net3223),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_2 _16832_ (.RESET_B(net510),
    .D(net3025),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_2 _16833_ (.RESET_B(net511),
    .D(net3046),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16834_ (.RESET_B(net512),
    .D(net3079),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16835_ (.RESET_B(net513),
    .D(net3205),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16836_ (.RESET_B(net514),
    .D(net3228),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _16837_ (.RESET_B(net515),
    .D(net3308),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16838_ (.RESET_B(net516),
    .D(net3002),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16839_ (.RESET_B(net517),
    .D(net3323),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16840_ (.RESET_B(net518),
    .D(net3137),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _16841_ (.RESET_B(net519),
    .D(net3112),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16842_ (.RESET_B(net520),
    .D(net3135),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16843_ (.RESET_B(net521),
    .D(net3062),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16844_ (.RESET_B(net522),
    .D(net3142),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _16845_ (.RESET_B(net523),
    .D(net3305),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _16846_ (.RESET_B(net524),
    .D(net3085),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16847_ (.RESET_B(net525),
    .D(net3109),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16848_ (.RESET_B(net526),
    .D(net3098),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _16849_ (.RESET_B(net527),
    .D(net3042),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _16850_ (.RESET_B(net528),
    .D(net3174),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16851_ (.RESET_B(net529),
    .D(net3003),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16852_ (.RESET_B(net530),
    .D(net3259),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _16853_ (.RESET_B(net531),
    .D(net3264),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _16854_ (.RESET_B(net532),
    .D(net3158),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16855_ (.RESET_B(net533),
    .D(net3172),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16856_ (.RESET_B(net534),
    .D(net3076),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _16857_ (.RESET_B(net535),
    .D(net3015),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _16858_ (.RESET_B(net536),
    .D(_00058_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _16859_ (.RESET_B(net537),
    .D(_00059_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _16860_ (.RESET_B(net538),
    .D(_00060_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _16861_ (.RESET_B(net539),
    .D(_00061_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _16862_ (.RESET_B(net540),
    .D(net3192),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16863_ (.RESET_B(net541),
    .D(net3128),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _16864_ (.RESET_B(net542),
    .D(net3056),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_2 _16865_ (.RESET_B(net543),
    .D(net3240),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16866_ (.RESET_B(net544),
    .D(net3036),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _16867_ (.RESET_B(net545),
    .D(net3242),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _16868_ (.RESET_B(net546),
    .D(net3222),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16869_ (.RESET_B(net547),
    .D(net3209),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16870_ (.RESET_B(net548),
    .D(net3226),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _16871_ (.RESET_B(net549),
    .D(net3173),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _16872_ (.RESET_B(net550),
    .D(net3130),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _16873_ (.RESET_B(net551),
    .D(net3275),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16874_ (.RESET_B(net552),
    .D(net3249),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16875_ (.RESET_B(net553),
    .D(net3219),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16876_ (.RESET_B(net554),
    .D(net3134),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16877_ (.RESET_B(net555),
    .D(net3118),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16878_ (.RESET_B(net556),
    .D(net3334),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16879_ (.RESET_B(net557),
    .D(net3328),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16880_ (.RESET_B(net558),
    .D(net3088),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16881_ (.RESET_B(net559),
    .D(net3167),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _16882_ (.RESET_B(net560),
    .D(net3282),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16883_ (.RESET_B(net561),
    .D(net3367),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16884_ (.RESET_B(net562),
    .D(net3251),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16885_ (.RESET_B(net563),
    .D(net3286),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _16886_ (.RESET_B(net564),
    .D(net3115),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16887_ (.RESET_B(net565),
    .D(net3069),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _16888_ (.RESET_B(net566),
    .D(net3238),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16889_ (.RESET_B(net567),
    .D(net3333),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _16890_ (.RESET_B(net568),
    .D(_00054_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16891_ (.RESET_B(net569),
    .D(_00055_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16892_ (.RESET_B(net570),
    .D(_00056_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _16893_ (.RESET_B(net571),
    .D(_00057_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _16894_ (.RESET_B(net572),
    .D(net3189),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_2 _16895_ (.RESET_B(net573),
    .D(net2984),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_2 _16896_ (.RESET_B(net574),
    .D(net3089),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_2 _16897_ (.RESET_B(net575),
    .D(net3337),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16898_ (.RESET_B(net576),
    .D(net3364),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16899_ (.RESET_B(net577),
    .D(net3294),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _16900_ (.RESET_B(net578),
    .D(net2990),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16901_ (.RESET_B(net579),
    .D(net3296),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16902_ (.RESET_B(net580),
    .D(net3161),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16903_ (.RESET_B(net581),
    .D(net3206),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16904_ (.RESET_B(net582),
    .D(net3303),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _16905_ (.RESET_B(net583),
    .D(net3129),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16906_ (.RESET_B(net584),
    .D(net3295),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16907_ (.RESET_B(net585),
    .D(net3262),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16908_ (.RESET_B(net586),
    .D(net3053),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16909_ (.RESET_B(net587),
    .D(net3171),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16910_ (.RESET_B(net588),
    .D(net3350),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16911_ (.RESET_B(net589),
    .D(net3061),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16912_ (.RESET_B(net590),
    .D(net3256),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16913_ (.RESET_B(net591),
    .D(net3151),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16914_ (.RESET_B(net592),
    .D(net3175),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _16915_ (.RESET_B(net593),
    .D(net3359),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16916_ (.RESET_B(net594),
    .D(net3245),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16917_ (.RESET_B(net595),
    .D(net3266),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16918_ (.RESET_B(net596),
    .D(net3084),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _16919_ (.RESET_B(net597),
    .D(net3106),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16920_ (.RESET_B(net598),
    .D(net3375),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16921_ (.RESET_B(net599),
    .D(net3361),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16922_ (.RESET_B(net600),
    .D(_00050_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _16923_ (.RESET_B(net601),
    .D(_00051_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16924_ (.RESET_B(net602),
    .D(_00052_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _16925_ (.RESET_B(net603),
    .D(_00053_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_2 _16926_ (.RESET_B(net604),
    .D(net3318),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16927_ (.RESET_B(net605),
    .D(net3201),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_2 _16928_ (.RESET_B(net606),
    .D(net3225),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_2 _16929_ (.RESET_B(net607),
    .D(net3178),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16930_ (.RESET_B(net608),
    .D(net3145),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _16931_ (.RESET_B(net609),
    .D(net3071),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16932_ (.RESET_B(net610),
    .D(net3059),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16933_ (.RESET_B(net611),
    .D(net3248),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16934_ (.RESET_B(net612),
    .D(net3067),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16935_ (.RESET_B(net613),
    .D(net3234),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16936_ (.RESET_B(net614),
    .D(net3196),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16937_ (.RESET_B(net615),
    .D(net3119),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16938_ (.RESET_B(net616),
    .D(net3016),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16939_ (.RESET_B(net617),
    .D(net3277),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16940_ (.RESET_B(net618),
    .D(net3306),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16941_ (.RESET_B(net619),
    .D(net3291),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16942_ (.RESET_B(net620),
    .D(net3074),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16943_ (.RESET_B(net621),
    .D(net3064),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16944_ (.RESET_B(net622),
    .D(net3021),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16945_ (.RESET_B(net623),
    .D(net3300),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16946_ (.RESET_B(net624),
    .D(net2996),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16947_ (.RESET_B(net625),
    .D(net3181),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16948_ (.RESET_B(net626),
    .D(net3329),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16949_ (.RESET_B(net627),
    .D(net2992),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16950_ (.RESET_B(net628),
    .D(net3150),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16951_ (.RESET_B(net629),
    .D(net3120),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16952_ (.RESET_B(net630),
    .D(net2998),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16953_ (.RESET_B(net631),
    .D(net3057),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16954_ (.RESET_B(net632),
    .D(_00046_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16955_ (.RESET_B(net633),
    .D(_00047_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16956_ (.RESET_B(net634),
    .D(_00048_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16957_ (.RESET_B(net635),
    .D(_00049_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_2 _16958_ (.RESET_B(net636),
    .D(net3163),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16959_ (.RESET_B(net637),
    .D(net3144),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16960_ (.RESET_B(net638),
    .D(net2991),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16961_ (.RESET_B(net639),
    .D(net3320),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16962_ (.RESET_B(net640),
    .D(net3028),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _16963_ (.RESET_B(net641),
    .D(net3193),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _16964_ (.RESET_B(net642),
    .D(net3343),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _16965_ (.RESET_B(net643),
    .D(net3371),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16966_ (.RESET_B(net644),
    .D(net3202),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _16967_ (.RESET_B(net645),
    .D(net3195),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16968_ (.RESET_B(net646),
    .D(net2989),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16969_ (.RESET_B(net647),
    .D(net3332),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16970_ (.RESET_B(net648),
    .D(net3045),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16971_ (.RESET_B(net649),
    .D(net3082),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16972_ (.RESET_B(net650),
    .D(net3139),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16973_ (.RESET_B(net651),
    .D(net3022),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16974_ (.RESET_B(net652),
    .D(net2986),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16975_ (.RESET_B(net653),
    .D(net3075),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16976_ (.RESET_B(net654),
    .D(net3070),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16977_ (.RESET_B(net655),
    .D(net3063),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16978_ (.RESET_B(net656),
    .D(net3335),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16979_ (.RESET_B(net657),
    .D(net3191),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16980_ (.RESET_B(net658),
    .D(net3060),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16981_ (.RESET_B(net659),
    .D(net3241),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16982_ (.RESET_B(net660),
    .D(net2988),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16983_ (.RESET_B(net661),
    .D(net3004),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16984_ (.RESET_B(net662),
    .D(net3008),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16985_ (.RESET_B(net663),
    .D(net3304),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16986_ (.RESET_B(net664),
    .D(_00094_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16987_ (.RESET_B(net665),
    .D(_00095_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16988_ (.RESET_B(net666),
    .D(_00096_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16989_ (.RESET_B(net667),
    .D(_00097_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_2 _16990_ (.RESET_B(net668),
    .D(net3325),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_2 _16991_ (.RESET_B(net669),
    .D(net3330),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_2 _16992_ (.RESET_B(net670),
    .D(net3159),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_2 _16993_ (.RESET_B(net671),
    .D(net3363),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16994_ (.RESET_B(net672),
    .D(net3273),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16995_ (.RESET_B(net673),
    .D(net3043),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16996_ (.RESET_B(net674),
    .D(net3312),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16997_ (.RESET_B(net675),
    .D(net3232),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16998_ (.RESET_B(net676),
    .D(net3237),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16999_ (.RESET_B(net677),
    .D(net3011),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _17000_ (.RESET_B(net678),
    .D(net3034),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _17001_ (.RESET_B(net679),
    .D(net3048),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _17002_ (.RESET_B(net680),
    .D(net3038),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _17003_ (.RESET_B(net681),
    .D(net3030),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _17004_ (.RESET_B(net682),
    .D(net3010),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _17005_ (.RESET_B(net683),
    .D(net3166),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _17006_ (.RESET_B(net684),
    .D(net3138),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _17007_ (.RESET_B(net685),
    .D(net3091),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _17008_ (.RESET_B(net686),
    .D(net3037),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _17009_ (.RESET_B(net687),
    .D(net3324),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _17010_ (.RESET_B(net688),
    .D(net3101),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _17011_ (.RESET_B(net689),
    .D(net3093),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _17012_ (.RESET_B(net690),
    .D(net3210),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _17013_ (.RESET_B(net691),
    .D(net3352),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _17014_ (.RESET_B(net692),
    .D(net3105),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _17015_ (.RESET_B(net693),
    .D(net3123),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _17016_ (.RESET_B(net694),
    .D(net3204),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _17017_ (.RESET_B(net695),
    .D(net3297),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _17018_ (.RESET_B(net696),
    .D(_00090_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _17019_ (.RESET_B(net697),
    .D(_00091_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _17020_ (.RESET_B(net698),
    .D(_00092_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _17021_ (.RESET_B(net699),
    .D(net4679),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_2 _17022_ (.RESET_B(net700),
    .D(net3177),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_2 _17023_ (.RESET_B(net701),
    .D(net3224),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_2 _17024_ (.RESET_B(net702),
    .D(net3218),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_2 _17025_ (.RESET_B(net703),
    .D(net3302),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _17026_ (.RESET_B(net704),
    .D(net3310),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _17027_ (.RESET_B(net705),
    .D(net3182),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _17028_ (.RESET_B(net706),
    .D(net3111),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17029_ (.RESET_B(net707),
    .D(net3019),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17030_ (.RESET_B(net708),
    .D(net3285),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17031_ (.RESET_B(net709),
    .D(net3292),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _17032_ (.RESET_B(net710),
    .D(net3289),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _17033_ (.RESET_B(net711),
    .D(net3319),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _17034_ (.RESET_B(net712),
    .D(net3261),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17035_ (.RESET_B(net713),
    .D(net3032),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _17036_ (.RESET_B(net714),
    .D(net3047),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _17037_ (.RESET_B(net715),
    .D(net3301),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17038_ (.RESET_B(net716),
    .D(net3327),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17039_ (.RESET_B(net717),
    .D(net3321),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _17040_ (.RESET_B(net718),
    .D(net3268),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _17041_ (.RESET_B(net719),
    .D(net2993),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17042_ (.RESET_B(net720),
    .D(net3152),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _17043_ (.RESET_B(net721),
    .D(net3169),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17044_ (.RESET_B(net722),
    .D(net3254),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17045_ (.RESET_B(net723),
    .D(net3230),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _17046_ (.RESET_B(net724),
    .D(net3346),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17047_ (.RESET_B(net725),
    .D(net3340),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17048_ (.RESET_B(net726),
    .D(net3336),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17049_ (.RESET_B(net727),
    .D(net3179),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _17050_ (.RESET_B(net728),
    .D(_00086_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _17051_ (.RESET_B(net729),
    .D(_00087_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _17052_ (.RESET_B(net730),
    .D(_00088_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17053_ (.RESET_B(net731),
    .D(_00089_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_2 _17054_ (.RESET_B(net732),
    .D(net3160),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_2 _17055_ (.RESET_B(net733),
    .D(net3117),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_2 _17056_ (.RESET_B(net734),
    .D(net2999),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_2 _17057_ (.RESET_B(net735),
    .D(net3143),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _17058_ (.RESET_B(net736),
    .D(net3132),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _17059_ (.RESET_B(net737),
    .D(net3229),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _17060_ (.RESET_B(net738),
    .D(net3366),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _17061_ (.RESET_B(net739),
    .D(net3214),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _17062_ (.RESET_B(net740),
    .D(net3197),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _17063_ (.RESET_B(net741),
    .D(net3362),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _17064_ (.RESET_B(net742),
    .D(net3017),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _17065_ (.RESET_B(net743),
    .D(net3354),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _17066_ (.RESET_B(net744),
    .D(net3341),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _17067_ (.RESET_B(net745),
    .D(net3188),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _17068_ (.RESET_B(net746),
    .D(net3035),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _17069_ (.RESET_B(net747),
    .D(net3039),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17070_ (.RESET_B(net748),
    .D(net3315),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17071_ (.RESET_B(net749),
    .D(net3227),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _17072_ (.RESET_B(net750),
    .D(net3131),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _17073_ (.RESET_B(net751),
    .D(net3066),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17074_ (.RESET_B(net752),
    .D(net3095),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _17075_ (.RESET_B(net753),
    .D(net3113),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17076_ (.RESET_B(net754),
    .D(net3149),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _17077_ (.RESET_B(net755),
    .D(net3073),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17078_ (.RESET_B(net756),
    .D(net3267),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _17079_ (.RESET_B(net757),
    .D(net3023),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17080_ (.RESET_B(net758),
    .D(net3054),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _17081_ (.RESET_B(net759),
    .D(net3026),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17082_ (.RESET_B(net760),
    .D(net4284),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _17083_ (.RESET_B(net761),
    .D(_00083_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _17084_ (.RESET_B(net762),
    .D(_00084_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _17085_ (.RESET_B(net763),
    .D(_00085_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _17086_ (.RESET_B(net764),
    .D(net3353),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_2 _17087_ (.RESET_B(net765),
    .D(net3348),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_2 _17088_ (.RESET_B(net766),
    .D(net3001),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_2 _17089_ (.RESET_B(net767),
    .D(net3108),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _17090_ (.RESET_B(net768),
    .D(net3027),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _17091_ (.RESET_B(net769),
    .D(net3272),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _17092_ (.RESET_B(net770),
    .D(net3338),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _17093_ (.RESET_B(net771),
    .D(net3221),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _17094_ (.RESET_B(net772),
    .D(net3052),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _17095_ (.RESET_B(net773),
    .D(net3121),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _17096_ (.RESET_B(net774),
    .D(net3000),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _17097_ (.RESET_B(net775),
    .D(net3287),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _17098_ (.RESET_B(net776),
    .D(net3090),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _17099_ (.RESET_B(net777),
    .D(net3153),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _17100_ (.RESET_B(net778),
    .D(net3215),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _17101_ (.RESET_B(net779),
    .D(net3009),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _17102_ (.RESET_B(net780),
    .D(net3356),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _17103_ (.RESET_B(net781),
    .D(net3199),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _17104_ (.RESET_B(net782),
    .D(net3257),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _17105_ (.RESET_B(net783),
    .D(net3200),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _17106_ (.RESET_B(net784),
    .D(net3216),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _17107_ (.RESET_B(net785),
    .D(net3339),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _17108_ (.RESET_B(net786),
    .D(net3055),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _17109_ (.RESET_B(net787),
    .D(net3217),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _17110_ (.RESET_B(net788),
    .D(net3345),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _17111_ (.RESET_B(net789),
    .D(net3372),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _17112_ (.RESET_B(net790),
    .D(net3376),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _17113_ (.RESET_B(net791),
    .D(net3157),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _17114_ (.RESET_B(net792),
    .D(_00078_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _17115_ (.RESET_B(net793),
    .D(_00079_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _17116_ (.RESET_B(net794),
    .D(_00080_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _17117_ (.RESET_B(net795),
    .D(_00081_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_2 _17118_ (.RESET_B(net796),
    .D(net2983),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_2 _17119_ (.RESET_B(net797),
    .D(net3190),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_2 _17120_ (.RESET_B(net798),
    .D(net3373),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_2 _17121_ (.RESET_B(net799),
    .D(net3049),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _17122_ (.RESET_B(net800),
    .D(net3146),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _17123_ (.RESET_B(net801),
    .D(net3165),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _17124_ (.RESET_B(net802),
    .D(net2985),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _17125_ (.RESET_B(net803),
    .D(net3370),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _17126_ (.RESET_B(net804),
    .D(net3299),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _17127_ (.RESET_B(net805),
    .D(net3126),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _17128_ (.RESET_B(net806),
    .D(net3369),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _17129_ (.RESET_B(net807),
    .D(net3243),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _17130_ (.RESET_B(net808),
    .D(net3187),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _17131_ (.RESET_B(net809),
    .D(net3087),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _17132_ (.RESET_B(net810),
    .D(net3006),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _17133_ (.RESET_B(net811),
    .D(net3051),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _17134_ (.RESET_B(net812),
    .D(net3012),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _17135_ (.RESET_B(net813),
    .D(net3344),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _17136_ (.RESET_B(net814),
    .D(net3198),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _17137_ (.RESET_B(net815),
    .D(net3020),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _17138_ (.RESET_B(net816),
    .D(net3133),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _17139_ (.RESET_B(net817),
    .D(net3342),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _17140_ (.RESET_B(net818),
    .D(net3044),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _17141_ (.RESET_B(net819),
    .D(net3239),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17142_ (.RESET_B(net820),
    .D(net3378),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _17143_ (.RESET_B(net821),
    .D(net3355),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _17144_ (.RESET_B(net822),
    .D(net3186),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _17145_ (.RESET_B(net823),
    .D(net3092),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _17146_ (.RESET_B(net824),
    .D(_00074_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _17147_ (.RESET_B(net825),
    .D(_00075_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _17148_ (.RESET_B(net826),
    .D(_00076_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _17149_ (.RESET_B(net827),
    .D(_00077_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _17150_ (.RESET_B(net828),
    .D(net3396),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _17151_ (.RESET_B(net829),
    .D(net3398),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_2 _17152_ (.RESET_B(net830),
    .D(net3403),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_2 _17153_ (.RESET_B(net831),
    .D(net3399),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_2 _17154_ (.RESET_B(net832),
    .D(net3387),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_2 _17155_ (.RESET_B(net833),
    .D(net3391),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_2 _17156_ (.RESET_B(net834),
    .D(net3392),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _17157_ (.RESET_B(net835),
    .D(net3382),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _17158_ (.RESET_B(net836),
    .D(net3388),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17159_ (.RESET_B(net837),
    .D(net3395),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17160_ (.RESET_B(net838),
    .D(net3389),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17161_ (.RESET_B(net839),
    .D(net3390),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _17162_ (.RESET_B(net840),
    .D(net3377),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _17163_ (.RESET_B(net841),
    .D(net3386),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _17164_ (.RESET_B(net842),
    .D(net3385),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17165_ (.RESET_B(net843),
    .D(net3381),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _17166_ (.RESET_B(net844),
    .D(net3384),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _17167_ (.RESET_B(net845),
    .D(net3374),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _17168_ (.RESET_B(net846),
    .D(net3380),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _17169_ (.RESET_B(net847),
    .D(net3379),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_1 _17170_ (.RESET_B(net848),
    .D(net3401),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_1 _17171_ (.RESET_B(net849),
    .D(net3404),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _17172_ (.RESET_B(net850),
    .D(net3400),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _17173_ (.RESET_B(net851),
    .D(net3402),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_2 _17174_ (.RESET_B(net852),
    .D(net3331),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_2 _17175_ (.RESET_B(net853),
    .D(net3211),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_2 _17176_ (.RESET_B(net854),
    .D(net3358),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_2 _17177_ (.RESET_B(net855),
    .D(net3326),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _17178_ (.RESET_B(net875),
    .D(\i_tinyqv.cpu.i_core.cy_out ),
    .Q(\i_tinyqv.cpu.i_core.cy ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _17179_ (.RESET_B(net1464),
    .D(\i_tinyqv.cpu.i_core.cmp_out ),
    .Q(\i_tinyqv.cpu.i_core.cmp ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_2 _17180_ (.RESET_B(net1463),
    .D(net4944),
    .Q(\crc16_read[8] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _17181_ (.RESET_B(net1461),
    .D(_00744_),
    .Q(\crc16_read[9] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _17182_ (.RESET_B(net1459),
    .D(_00745_),
    .Q(\crc16_read[10] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17183_ (.RESET_B(net1457),
    .D(net4939),
    .Q(\crc16_read[11] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17184_ (.RESET_B(net1455),
    .D(net4753),
    .Q(\crc16_read[12] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _17185_ (.RESET_B(net1453),
    .D(_00748_),
    .Q(\crc16_read[13] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17186_ (.RESET_B(net1451),
    .D(net4786),
    .Q(\crc16_read[14] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17187_ (.RESET_B(net1449),
    .D(_00750_),
    .Q(\crc16_read[15] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_1 _17188_ (.RESET_B(net1447),
    .D(net3867),
    .Q(\i_tinyqv.cpu.i_core.load_done ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_2 _17189_ (.RESET_B(net1446),
    .D(_00752_),
    .Q(\i_tinyqv.cpu.i_core.cycle[0] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _17190_ (.RESET_B(net1444),
    .D(_00753_),
    .Q(\i_tinyqv.cpu.i_core.cycle[1] ),
    .CLK(clknet_leaf_178_clk_regs));
 sg13g2_dfrbpq_1 _17191_ (.RESET_B(net1442),
    .D(_00754_),
    .Q(\i_i2c_peri.i_i2c.bit_count_reg[0] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _17192_ (.RESET_B(net1440),
    .D(_00755_),
    .Q(\i_i2c_peri.i_i2c.bit_count_reg[1] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _17193_ (.RESET_B(net1438),
    .D(_00756_),
    .Q(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _17194_ (.RESET_B(net1436),
    .D(net4866),
    .Q(\i_i2c_peri.i_i2c.bit_count_reg[3] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _17195_ (.RESET_B(net1434),
    .D(net3615),
    .Q(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_1 _17196_ (.RESET_B(net1433),
    .D(_00759_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _17197_ (.RESET_B(net1431),
    .D(_00760_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _17198_ (.RESET_B(net914),
    .D(net3961),
    .Q(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _17199_ (.RESET_B(net1429),
    .D(_00045_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.add ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _17200_ (.RESET_B(net1427),
    .D(net4152),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _17201_ (.RESET_B(net1426),
    .D(net4206),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_2 _17202_ (.RESET_B(net1425),
    .D(net4062),
    .Q(\i_tinyqv.cpu.i_core.mepc[20] ),
    .CLK(clknet_leaf_180_clk_regs));
 sg13g2_dfrbpq_1 _17203_ (.RESET_B(net1423),
    .D(_00765_),
    .Q(\i_tinyqv.cpu.i_core.mepc[21] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_1 _17204_ (.RESET_B(net1421),
    .D(net4276),
    .Q(\i_tinyqv.cpu.i_core.mepc[22] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _17205_ (.RESET_B(net1419),
    .D(net4351),
    .Q(\i_tinyqv.cpu.i_core.mepc[23] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _17206_ (.RESET_B(net1417),
    .D(_00768_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_2 _17207_ (.RESET_B(net1415),
    .D(_00769_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _17208_ (.RESET_B(net1413),
    .D(net3965),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_2 _17209_ (.RESET_B(net1411),
    .D(_00771_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_2 _17210_ (.RESET_B(net1410),
    .D(net4106),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_2 _17211_ (.RESET_B(net1409),
    .D(_00773_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _17212_ (.RESET_B(net1408),
    .D(_00774_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _17213_ (.RESET_B(net1407),
    .D(_00775_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _17214_ (.RESET_B(net1406),
    .D(net4212),
    .Q(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _17215_ (.RESET_B(net1405),
    .D(net3839),
    .Q(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17216_ (.RESET_B(net1404),
    .D(_00778_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17217_ (.RESET_B(net1403),
    .D(net3829),
    .Q(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17218_ (.RESET_B(net1402),
    .D(net4773),
    .Q(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17219_ (.RESET_B(net1401),
    .D(net3604),
    .Q(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17220_ (.RESET_B(net1400),
    .D(_00782_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17221_ (.RESET_B(net1399),
    .D(net3628),
    .Q(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _17222_ (.RESET_B(net1398),
    .D(net3750),
    .Q(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17223_ (.RESET_B(net1397),
    .D(_00785_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17224_ (.RESET_B(net1396),
    .D(net3626),
    .Q(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17225_ (.RESET_B(net1395),
    .D(net4286),
    .Q(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _17226_ (.RESET_B(net1394),
    .D(_00788_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17227_ (.RESET_B(net1393),
    .D(_00789_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17228_ (.RESET_B(net1392),
    .D(net3888),
    .Q(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17229_ (.RESET_B(net1391),
    .D(_00791_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _17230_ (.RESET_B(net1390),
    .D(net3815),
    .Q(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _17231_ (.RESET_B(net1389),
    .D(_00793_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17232_ (.RESET_B(net1388),
    .D(net4390),
    .Q(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17233_ (.RESET_B(net1387),
    .D(net3943),
    .Q(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17234_ (.RESET_B(net1385),
    .D(_00796_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17235_ (.RESET_B(net1383),
    .D(net3567),
    .Q(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _17236_ (.RESET_B(net1381),
    .D(net3977),
    .Q(\i_tinyqv.cpu.instr_data[2][0] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _17237_ (.RESET_B(net915),
    .D(net3911),
    .Q(\i_tinyqv.cpu.instr_data[2][1] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17238_ (.RESET_B(net916),
    .D(_00070_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _17239_ (.RESET_B(net917),
    .D(_00071_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _17240_ (.RESET_B(net918),
    .D(_00072_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _17241_ (.RESET_B(net1228),
    .D(_00073_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _17242_ (.RESET_B(net1379),
    .D(net2620),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _17243_ (.RESET_B(net1377),
    .D(net3482),
    .Q(\i_crc16.bit_cnt[0] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _17244_ (.RESET_B(net1375),
    .D(_00801_),
    .Q(\i_crc16.bit_cnt[1] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _17245_ (.RESET_B(net1372),
    .D(net4172),
    .Q(\i_crc16.bit_cnt[2] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _17246_ (.RESET_B(net1370),
    .D(_00803_),
    .Q(\i_wdt.enabled ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17247_ (.RESET_B(net1368),
    .D(_00804_),
    .Q(\i_wdt.counter[0] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17248_ (.RESET_B(net1366),
    .D(net5144),
    .Q(\i_wdt.counter[1] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17249_ (.RESET_B(net1364),
    .D(_00806_),
    .Q(\i_wdt.counter[2] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17250_ (.RESET_B(net1362),
    .D(net4629),
    .Q(\i_wdt.counter[3] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17251_ (.RESET_B(net1360),
    .D(_00808_),
    .Q(\i_wdt.counter[4] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17252_ (.RESET_B(net1358),
    .D(net4718),
    .Q(\i_wdt.counter[5] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17253_ (.RESET_B(net1356),
    .D(_00810_),
    .Q(\i_wdt.counter[6] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17254_ (.RESET_B(net1354),
    .D(net4396),
    .Q(\i_wdt.counter[7] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17255_ (.RESET_B(net1352),
    .D(_00812_),
    .Q(\i_wdt.counter[8] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17256_ (.RESET_B(net1350),
    .D(_00813_),
    .Q(\i_wdt.counter[9] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17257_ (.RESET_B(net1348),
    .D(_00814_),
    .Q(\i_wdt.counter[10] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17258_ (.RESET_B(net1346),
    .D(_00815_),
    .Q(\i_wdt.counter[11] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _17259_ (.RESET_B(net1344),
    .D(_00816_),
    .Q(\i_wdt.counter[12] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _17260_ (.RESET_B(net1342),
    .D(_00817_),
    .Q(\i_wdt.counter[13] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _17261_ (.RESET_B(net1340),
    .D(net5212),
    .Q(\i_wdt.counter[14] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _17262_ (.RESET_B(net1338),
    .D(_00819_),
    .Q(\i_wdt.counter[15] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _17263_ (.RESET_B(net1335),
    .D(_00820_),
    .Q(\i_wdt.counter[16] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _17264_ (.RESET_B(net1333),
    .D(net4819),
    .Q(\i_wdt.counter[17] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _17265_ (.RESET_B(net1331),
    .D(net5028),
    .Q(\i_wdt.counter[18] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _17266_ (.RESET_B(net1329),
    .D(net4703),
    .Q(\i_wdt.counter[19] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _17267_ (.RESET_B(net1327),
    .D(_00824_),
    .Q(\i_wdt.counter[20] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _17268_ (.RESET_B(net1325),
    .D(net4665),
    .Q(\i_wdt.counter[21] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _17269_ (.RESET_B(net1323),
    .D(_00826_),
    .Q(\i_wdt.counter[22] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _17270_ (.RESET_B(net1321),
    .D(_00827_),
    .Q(\i_wdt.counter[23] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _17271_ (.RESET_B(net1319),
    .D(net4238),
    .Q(\i_wdt.counter[24] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17272_ (.RESET_B(net1317),
    .D(net4266),
    .Q(\i_wdt.counter[25] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_2 _17273_ (.RESET_B(net1315),
    .D(net4433),
    .Q(\i_wdt.counter[26] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17274_ (.RESET_B(net1313),
    .D(_00831_),
    .Q(\i_wdt.counter[27] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17275_ (.RESET_B(net1311),
    .D(net4894),
    .Q(\i_wdt.counter[28] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _17276_ (.RESET_B(net1309),
    .D(_00833_),
    .Q(\i_wdt.counter[29] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _17277_ (.RESET_B(net1307),
    .D(net4348),
    .Q(\i_wdt.counter[30] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _17278_ (.RESET_B(net1305),
    .D(net4392),
    .Q(\i_wdt.counter[31] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _17279_ (.RESET_B(net1303),
    .D(net4941),
    .Q(\i_uart_tx.txd_reg ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _17280_ (.RESET_B(net1302),
    .D(_00837_),
    .Q(\i_rtc.us_count[0] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _17281_ (.RESET_B(net1300),
    .D(net3769),
    .Q(\i_rtc.us_count[1] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_2 _17282_ (.RESET_B(net1298),
    .D(net3522),
    .Q(\i_rtc.us_count[2] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _17283_ (.RESET_B(net1296),
    .D(_00840_),
    .Q(\i_rtc.us_count[3] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_2 _17284_ (.RESET_B(net1294),
    .D(_00841_),
    .Q(\i_rtc.us_count[4] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_2 _17285_ (.RESET_B(net1292),
    .D(_00842_),
    .Q(\i_rtc.us_count[5] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_2 _17286_ (.RESET_B(net1290),
    .D(_00843_),
    .Q(\i_rtc.us_count[6] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_2 _17287_ (.RESET_B(net1288),
    .D(_00844_),
    .Q(\i_rtc.us_count[7] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _17288_ (.RESET_B(net1286),
    .D(net4014),
    .Q(\i_rtc.us_count[8] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _17289_ (.RESET_B(net1284),
    .D(net4502),
    .Q(\i_rtc.us_count[9] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _17290_ (.RESET_B(net1282),
    .D(_00847_),
    .Q(\i_rtc.us_count[10] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_2 _17291_ (.RESET_B(net1280),
    .D(_00848_),
    .Q(\i_rtc.us_count[11] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_2 _17292_ (.RESET_B(net1278),
    .D(net4218),
    .Q(\i_rtc.us_count[12] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_2 _17293_ (.RESET_B(net1276),
    .D(_00850_),
    .Q(\i_rtc.us_count[13] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _17294_ (.RESET_B(net1274),
    .D(_00851_),
    .Q(\i_rtc.us_count[14] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _17295_ (.RESET_B(net1272),
    .D(net4307),
    .Q(\i_rtc.us_count[15] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _17296_ (.RESET_B(net1270),
    .D(_00853_),
    .Q(\i_rtc.us_count[16] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_2 _17297_ (.RESET_B(net1268),
    .D(net3608),
    .Q(\i_rtc.us_count[17] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _17298_ (.RESET_B(net1266),
    .D(_00855_),
    .Q(\i_rtc.us_count[18] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _17299_ (.RESET_B(net1264),
    .D(_00856_),
    .Q(\i_rtc.us_count[19] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_2 _17300_ (.RESET_B(net1262),
    .D(_00857_),
    .Q(\i_rtc.seconds_out[0] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17301_ (.RESET_B(net1260),
    .D(_00858_),
    .Q(\i_rtc.seconds_out[1] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17302_ (.RESET_B(net1258),
    .D(_00859_),
    .Q(\i_rtc.seconds_out[2] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _17303_ (.RESET_B(net1256),
    .D(_00860_),
    .Q(\i_rtc.seconds_out[3] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17304_ (.RESET_B(net1254),
    .D(_00861_),
    .Q(\i_rtc.seconds_out[4] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17305_ (.RESET_B(net1252),
    .D(_00862_),
    .Q(\i_rtc.seconds_out[5] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17306_ (.RESET_B(net1250),
    .D(_00863_),
    .Q(\i_rtc.seconds_out[6] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _17307_ (.RESET_B(net1248),
    .D(_00864_),
    .Q(\i_rtc.seconds_out[7] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17308_ (.RESET_B(net1246),
    .D(_00865_),
    .Q(\i_rtc.seconds_out[8] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _17309_ (.RESET_B(net1244),
    .D(_00866_),
    .Q(\i_rtc.seconds_out[9] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _17310_ (.RESET_B(net1242),
    .D(net5233),
    .Q(\i_rtc.seconds_out[10] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _17311_ (.RESET_B(net1240),
    .D(net5183),
    .Q(\i_rtc.seconds_out[11] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _17312_ (.RESET_B(net1226),
    .D(net5294),
    .Q(\i_rtc.seconds_out[12] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _17313_ (.RESET_B(net1224),
    .D(_00870_),
    .Q(\i_rtc.seconds_out[13] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _17314_ (.RESET_B(net1222),
    .D(_00871_),
    .Q(\i_rtc.seconds_out[14] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _17315_ (.RESET_B(net1220),
    .D(_00872_),
    .Q(\i_rtc.seconds_out[15] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_2 _17316_ (.RESET_B(net1218),
    .D(_00873_),
    .Q(\i_rtc.seconds_out[16] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _17317_ (.RESET_B(net1216),
    .D(_00874_),
    .Q(\i_rtc.seconds_out[17] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_2 _17318_ (.RESET_B(net1214),
    .D(_00875_),
    .Q(\i_rtc.seconds_out[18] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _17319_ (.RESET_B(net1212),
    .D(_00876_),
    .Q(\i_rtc.seconds_out[19] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_2 _17320_ (.RESET_B(net1210),
    .D(_00877_),
    .Q(\i_rtc.seconds_out[20] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _17321_ (.RESET_B(net1208),
    .D(_00878_),
    .Q(\i_rtc.seconds_out[21] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _17322_ (.RESET_B(net1206),
    .D(_00879_),
    .Q(\i_rtc.seconds_out[22] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _17323_ (.RESET_B(net1204),
    .D(_00880_),
    .Q(\i_rtc.seconds_out[23] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _17324_ (.RESET_B(net1202),
    .D(net4735),
    .Q(\i_rtc.seconds_out[24] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _17325_ (.RESET_B(net1200),
    .D(_00882_),
    .Q(\i_rtc.seconds_out[25] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _17326_ (.RESET_B(net1198),
    .D(net5089),
    .Q(\i_rtc.seconds_out[26] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _17327_ (.RESET_B(net1196),
    .D(net5080),
    .Q(\i_rtc.seconds_out[27] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _17328_ (.RESET_B(net1194),
    .D(_00885_),
    .Q(\i_rtc.seconds_out[28] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _17329_ (.RESET_B(net1192),
    .D(_00886_),
    .Q(\i_rtc.seconds_out[29] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _17330_ (.RESET_B(net1190),
    .D(_00887_),
    .Q(\i_rtc.seconds_out[30] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _17331_ (.RESET_B(net1188),
    .D(net5021),
    .Q(\i_rtc.seconds_out[31] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_2 _17332_ (.RESET_B(net1186),
    .D(_00889_),
    .Q(\i_seal.crc_feed ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _17333_ (.RESET_B(net1185),
    .D(_00890_),
    .Q(\i_seal.byte_sent ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _17334_ (.RESET_B(net1183),
    .D(_00891_),
    .Q(\i_seal.byte_idx[0] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _17335_ (.RESET_B(net1181),
    .D(_00892_),
    .Q(\i_seal.byte_idx[1] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _17336_ (.RESET_B(net1179),
    .D(_00893_),
    .Q(\i_seal.byte_idx[2] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _17337_ (.RESET_B(net1177),
    .D(net5121),
    .Q(\i_seal.byte_idx[3] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _17338_ (.RESET_B(net1175),
    .D(net4683),
    .Q(\i_seal.sealed_crc[0] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _17339_ (.RESET_B(net1173),
    .D(net4688),
    .Q(\i_seal.sealed_crc[1] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _17340_ (.RESET_B(net1171),
    .D(net4748),
    .Q(\i_seal.sealed_crc[2] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _17341_ (.RESET_B(net1169),
    .D(net4844),
    .Q(\i_seal.sealed_crc[3] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _17342_ (.RESET_B(net1167),
    .D(net4720),
    .Q(\i_seal.sealed_crc[4] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _17343_ (.RESET_B(net1165),
    .D(net4528),
    .Q(\i_seal.sealed_crc[5] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _17344_ (.RESET_B(net1163),
    .D(net4587),
    .Q(\i_seal.sealed_crc[6] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _17345_ (.RESET_B(net1161),
    .D(net4530),
    .Q(\i_seal.sealed_crc[7] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _17346_ (.RESET_B(net1159),
    .D(net3555),
    .Q(\i_seal.sealed_crc[8] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _17347_ (.RESET_B(net1157),
    .D(net3678),
    .Q(\i_seal.sealed_crc[9] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _17348_ (.RESET_B(net1155),
    .D(net3565),
    .Q(\i_seal.sealed_crc[10] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17349_ (.RESET_B(net1153),
    .D(net3545),
    .Q(\i_seal.sealed_crc[11] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _17350_ (.RESET_B(net1151),
    .D(net3669),
    .Q(\i_seal.sealed_crc[12] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _17351_ (.RESET_B(net1149),
    .D(net4654),
    .Q(\i_seal.sealed_crc[13] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _17352_ (.RESET_B(net1147),
    .D(net3589),
    .Q(\i_seal.sealed_crc[14] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _17353_ (.RESET_B(net1145),
    .D(net3569),
    .Q(\i_seal.sealed_crc[15] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _17354_ (.RESET_B(net1143),
    .D(net4188),
    .Q(\i_seal.sealed_mono[0] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _17355_ (.RESET_B(net1141),
    .D(net4111),
    .Q(\i_seal.sealed_mono[1] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _17356_ (.RESET_B(net1139),
    .D(net4080),
    .Q(\i_seal.sealed_mono[2] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _17357_ (.RESET_B(net1137),
    .D(net4627),
    .Q(\i_seal.sealed_mono[3] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _17358_ (.RESET_B(net1135),
    .D(net4115),
    .Q(\i_seal.sealed_mono[4] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _17359_ (.RESET_B(net1133),
    .D(_00916_),
    .Q(\i_seal.sealed_mono[5] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _17360_ (.RESET_B(net1131),
    .D(net4577),
    .Q(\i_seal.sealed_mono[6] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17361_ (.RESET_B(net1129),
    .D(net4254),
    .Q(\i_seal.sealed_mono[7] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17362_ (.RESET_B(net1127),
    .D(_00919_),
    .Q(\i_seal.sealed_mono[8] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17363_ (.RESET_B(net1125),
    .D(net4639),
    .Q(\i_seal.sealed_mono[9] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _17364_ (.RESET_B(net1123),
    .D(net4556),
    .Q(\i_seal.sealed_mono[10] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _17365_ (.RESET_B(net1121),
    .D(net3923),
    .Q(\i_seal.sealed_mono[11] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _17366_ (.RESET_B(net1119),
    .D(net3766),
    .Q(\i_seal.sealed_mono[12] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _17367_ (.RESET_B(net1117),
    .D(_00924_),
    .Q(\i_seal.sealed_mono[13] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _17368_ (.RESET_B(net1115),
    .D(net4778),
    .Q(\i_seal.sealed_mono[14] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _17369_ (.RESET_B(net1113),
    .D(net3947),
    .Q(\i_seal.sealed_mono[15] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _17370_ (.RESET_B(net1111),
    .D(net4656),
    .Q(\i_seal.sealed_mono[16] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17371_ (.RESET_B(net1109),
    .D(net4148),
    .Q(\i_seal.sealed_mono[17] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _17372_ (.RESET_B(net1107),
    .D(_00929_),
    .Q(\i_seal.sealed_mono[18] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17373_ (.RESET_B(net1105),
    .D(_00930_),
    .Q(\i_seal.sealed_mono[19] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17374_ (.RESET_B(net1103),
    .D(net4544),
    .Q(\i_seal.sealed_mono[20] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17375_ (.RESET_B(net1101),
    .D(net4337),
    .Q(\i_seal.sealed_mono[21] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _17376_ (.RESET_B(net1099),
    .D(net4560),
    .Q(\i_seal.sealed_mono[22] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _17377_ (.RESET_B(net1097),
    .D(net4366),
    .Q(\i_seal.sealed_mono[23] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _17378_ (.RESET_B(net1095),
    .D(net4174),
    .Q(\i_seal.sealed_mono[24] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _17379_ (.RESET_B(net1093),
    .D(net3826),
    .Q(\i_seal.sealed_mono[25] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _17380_ (.RESET_B(net1091),
    .D(net3983),
    .Q(\i_seal.sealed_mono[26] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _17381_ (.RESET_B(net1089),
    .D(net4143),
    .Q(\i_seal.sealed_mono[27] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17382_ (.RESET_B(net1087),
    .D(net3845),
    .Q(\i_seal.sealed_mono[28] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _17383_ (.RESET_B(net1085),
    .D(_00940_),
    .Q(\i_seal.sealed_mono[29] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17384_ (.RESET_B(net1083),
    .D(_00941_),
    .Q(\i_seal.sealed_mono[30] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _17385_ (.RESET_B(net1081),
    .D(_00942_),
    .Q(\i_seal.sealed_mono[31] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17386_ (.RESET_B(net1079),
    .D(net4542),
    .Q(\i_seal.sealed_value[0] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _17387_ (.RESET_B(net1077),
    .D(net4573),
    .Q(\i_seal.sealed_value[1] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _17388_ (.RESET_B(net1075),
    .D(net4421),
    .Q(\i_seal.sealed_value[2] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _17389_ (.RESET_B(net1073),
    .D(net4480),
    .Q(\i_seal.sealed_value[3] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _17390_ (.RESET_B(net1071),
    .D(net3957),
    .Q(\i_seal.sealed_value[4] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17391_ (.RESET_B(net1069),
    .D(net4444),
    .Q(\i_seal.sealed_value[5] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17392_ (.RESET_B(net1067),
    .D(net3951),
    .Q(\i_seal.sealed_value[6] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17393_ (.RESET_B(net1065),
    .D(net3927),
    .Q(\i_seal.sealed_value[7] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17394_ (.RESET_B(net1063),
    .D(net3786),
    .Q(\i_seal.sealed_value[8] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _17395_ (.RESET_B(net1061),
    .D(net4198),
    .Q(\i_seal.sealed_value[9] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _17396_ (.RESET_B(net1059),
    .D(net4268),
    .Q(\i_seal.sealed_value[10] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17397_ (.RESET_B(net1057),
    .D(net4431),
    .Q(\i_seal.sealed_value[11] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _17398_ (.RESET_B(net1055),
    .D(net4597),
    .Q(\i_seal.sealed_value[12] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _17399_ (.RESET_B(net1053),
    .D(net4222),
    .Q(\i_seal.sealed_value[13] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _17400_ (.RESET_B(net1051),
    .D(net4030),
    .Q(\i_seal.sealed_value[14] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _17401_ (.RESET_B(net1049),
    .D(net4119),
    .Q(\i_seal.sealed_value[15] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _17402_ (.RESET_B(net1047),
    .D(net4006),
    .Q(\i_seal.sealed_value[16] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _17403_ (.RESET_B(net1045),
    .D(net3963),
    .Q(\i_seal.sealed_value[17] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17404_ (.RESET_B(net1043),
    .D(net4017),
    .Q(\i_seal.sealed_value[18] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17405_ (.RESET_B(net1041),
    .D(net4318),
    .Q(\i_seal.sealed_value[19] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _17406_ (.RESET_B(net1039),
    .D(net4008),
    .Q(\i_seal.sealed_value[20] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17407_ (.RESET_B(net1037),
    .D(net4156),
    .Q(\i_seal.sealed_value[21] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _17408_ (.RESET_B(net1035),
    .D(net4099),
    .Q(\i_seal.sealed_value[22] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17409_ (.RESET_B(net1033),
    .D(net4135),
    .Q(\i_seal.sealed_value[23] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _17410_ (.RESET_B(net1031),
    .D(net4190),
    .Q(\i_seal.sealed_value[24] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _17411_ (.RESET_B(net1029),
    .D(net4394),
    .Q(\i_seal.sealed_value[25] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _17412_ (.RESET_B(net1027),
    .D(net4325),
    .Q(\i_seal.sealed_value[26] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _17413_ (.RESET_B(net1025),
    .D(net4328),
    .Q(\i_seal.sealed_value[27] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _17414_ (.RESET_B(net1023),
    .D(net4072),
    .Q(\i_seal.sealed_value[28] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _17415_ (.RESET_B(net1021),
    .D(net4383),
    .Q(\i_seal.sealed_value[29] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _17416_ (.RESET_B(net1019),
    .D(net4078),
    .Q(\i_seal.sealed_value[30] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17417_ (.RESET_B(net1017),
    .D(net4228),
    .Q(\i_seal.sealed_value[31] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17418_ (.RESET_B(net1015),
    .D(_00975_),
    .Q(\i_seal.session_locked ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17419_ (.RESET_B(net1013),
    .D(net4086),
    .Q(\i_seal.sealed_sid[0] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _17420_ (.RESET_B(net1011),
    .D(net3790),
    .Q(\i_seal.sealed_sid[1] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _17421_ (.RESET_B(net1009),
    .D(net4312),
    .Q(\i_seal.sealed_sid[2] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _17422_ (.RESET_B(net1007),
    .D(net4139),
    .Q(\i_seal.sealed_sid[3] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _17423_ (.RESET_B(net1005),
    .D(_00980_),
    .Q(\i_seal.sealed_sid[4] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _17424_ (.RESET_B(net1003),
    .D(net3886),
    .Q(\i_seal.sealed_sid[5] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _17425_ (.RESET_B(net1001),
    .D(net3929),
    .Q(\i_seal.sealed_sid[6] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _17426_ (.RESET_B(net999),
    .D(net3994),
    .Q(\i_seal.sealed_sid[7] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _17427_ (.RESET_B(net997),
    .D(_00984_),
    .Q(\i_seal.mono_count[0] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _17428_ (.RESET_B(net995),
    .D(_00985_),
    .Q(\i_seal.mono_count[1] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _17429_ (.RESET_B(net993),
    .D(net4053),
    .Q(\i_seal.mono_count[2] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _17430_ (.RESET_B(net991),
    .D(_00987_),
    .Q(\i_seal.mono_count[3] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _17431_ (.RESET_B(net989),
    .D(_00988_),
    .Q(\i_seal.mono_count[4] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _17432_ (.RESET_B(net987),
    .D(_00989_),
    .Q(\i_seal.mono_count[5] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _17433_ (.RESET_B(net985),
    .D(net3891),
    .Q(\i_seal.mono_count[6] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_2 _17434_ (.RESET_B(net983),
    .D(_00991_),
    .Q(\i_seal.mono_count[7] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _17435_ (.RESET_B(net981),
    .D(net3933),
    .Q(\i_seal.mono_count[8] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _17436_ (.RESET_B(net979),
    .D(_00993_),
    .Q(\i_seal.mono_count[9] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _17437_ (.RESET_B(net977),
    .D(_00994_),
    .Q(\i_seal.mono_count[10] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_2 _17438_ (.RESET_B(net975),
    .D(_00995_),
    .Q(\i_seal.mono_count[11] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _17439_ (.RESET_B(net973),
    .D(net3897),
    .Q(\i_seal.mono_count[12] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_2 _17440_ (.RESET_B(net971),
    .D(_00997_),
    .Q(\i_seal.mono_count[13] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _17441_ (.RESET_B(net969),
    .D(_00998_),
    .Q(\i_seal.mono_count[14] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _17442_ (.RESET_B(net967),
    .D(_00999_),
    .Q(\i_seal.mono_count[15] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _17443_ (.RESET_B(net965),
    .D(_01000_),
    .Q(\i_seal.mono_count[16] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _17444_ (.RESET_B(net963),
    .D(_01001_),
    .Q(\i_seal.mono_count[17] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _17445_ (.RESET_B(net961),
    .D(net3973),
    .Q(\i_seal.mono_count[18] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _17446_ (.RESET_B(net959),
    .D(_01003_),
    .Q(\i_seal.mono_count[19] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _17447_ (.RESET_B(net957),
    .D(_01004_),
    .Q(\i_seal.mono_count[20] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _17448_ (.RESET_B(net955),
    .D(_01005_),
    .Q(\i_seal.mono_count[21] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _17449_ (.RESET_B(net953),
    .D(_01006_),
    .Q(\i_seal.mono_count[22] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _17450_ (.RESET_B(net951),
    .D(_01007_),
    .Q(\i_seal.mono_count[23] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _17451_ (.RESET_B(net949),
    .D(_01008_),
    .Q(\i_seal.mono_count[24] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_2 _17452_ (.RESET_B(net947),
    .D(_01009_),
    .Q(\i_seal.mono_count[25] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _17453_ (.RESET_B(net945),
    .D(net3552),
    .Q(\i_seal.mono_count[26] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _17454_ (.RESET_B(net943),
    .D(_01011_),
    .Q(\i_seal.mono_count[27] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _17455_ (.RESET_B(net941),
    .D(_01012_),
    .Q(\i_seal.mono_count[28] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_2 _17456_ (.RESET_B(net939),
    .D(net3540),
    .Q(\i_seal.mono_count[29] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _17457_ (.RESET_B(net937),
    .D(net3687),
    .Q(\i_seal.mono_count[30] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _17458_ (.RESET_B(net935),
    .D(net3938),
    .Q(\i_seal.mono_count[31] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _17459_ (.RESET_B(net933),
    .D(_01016_),
    .Q(\i_seal.cur_mono[0] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_2 _17460_ (.RESET_B(net931),
    .D(_01017_),
    .Q(\i_seal.cur_mono[1] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_2 _17461_ (.RESET_B(net929),
    .D(_01018_),
    .Q(\i_seal.cur_mono[2] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_2 _17462_ (.RESET_B(net927),
    .D(net3955),
    .Q(\i_seal.cur_mono[3] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _17463_ (.RESET_B(net925),
    .D(_01020_),
    .Q(\i_seal.cur_mono[4] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _17464_ (.RESET_B(net923),
    .D(_01021_),
    .Q(\i_seal.cur_mono[5] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_2 _17465_ (.RESET_B(net921),
    .D(net3714),
    .Q(\i_seal.cur_mono[6] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _17466_ (.RESET_B(net919),
    .D(_01023_),
    .Q(\i_seal.cur_mono[7] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _17467_ (.RESET_B(net912),
    .D(_01024_),
    .Q(\i_seal.cur_mono[8] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _17468_ (.RESET_B(net910),
    .D(net3655),
    .Q(\i_seal.cur_mono[9] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_2 _17469_ (.RESET_B(net908),
    .D(net3728),
    .Q(\i_seal.cur_mono[10] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_2 _17470_ (.RESET_B(net906),
    .D(_01027_),
    .Q(\i_seal.cur_mono[11] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_2 _17471_ (.RESET_B(net904),
    .D(_01028_),
    .Q(\i_seal.cur_mono[12] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _17472_ (.RESET_B(net902),
    .D(_01029_),
    .Q(\i_seal.cur_mono[13] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _17473_ (.RESET_B(net900),
    .D(net3865),
    .Q(\i_seal.cur_mono[14] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_2 _17474_ (.RESET_B(net898),
    .D(net3871),
    .Q(\i_seal.cur_mono[15] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _17475_ (.RESET_B(net896),
    .D(net3893),
    .Q(\i_seal.cur_mono[16] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _17476_ (.RESET_B(net894),
    .D(net4040),
    .Q(\i_seal.cur_mono[17] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _17477_ (.RESET_B(net892),
    .D(_01034_),
    .Q(\i_seal.cur_mono[18] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_2 _17478_ (.RESET_B(net890),
    .D(_01035_),
    .Q(\i_seal.cur_mono[19] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_2 _17479_ (.RESET_B(net888),
    .D(net3666),
    .Q(\i_seal.cur_mono[20] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_2 _17480_ (.RESET_B(net886),
    .D(net3836),
    .Q(\i_seal.cur_mono[21] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _17481_ (.RESET_B(net884),
    .D(net4032),
    .Q(\i_seal.cur_mono[22] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_2 _17482_ (.RESET_B(net882),
    .D(net4000),
    .Q(\i_seal.cur_mono[23] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _17483_ (.RESET_B(net880),
    .D(net3674),
    .Q(\i_seal.cur_mono[24] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _17484_ (.RESET_B(net878),
    .D(_01041_),
    .Q(\i_seal.cur_mono[25] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _17485_ (.RESET_B(net876),
    .D(_01042_),
    .Q(\i_seal.cur_mono[26] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_2 _17486_ (.RESET_B(net873),
    .D(net3918),
    .Q(\i_seal.cur_mono[27] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_2 _17487_ (.RESET_B(net871),
    .D(_01044_),
    .Q(\i_seal.cur_mono[28] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_2 _17488_ (.RESET_B(net869),
    .D(_01045_),
    .Q(\i_seal.cur_mono[29] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_2 _17489_ (.RESET_B(net867),
    .D(_01046_),
    .Q(\i_seal.cur_mono[30] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_2 _17490_ (.RESET_B(net865),
    .D(_01047_),
    .Q(\i_seal.cur_mono[31] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _17491_ (.RESET_B(net863),
    .D(net3528),
    .Q(\i_seal.sensor_id_reg[0] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _17492_ (.RESET_B(net861),
    .D(net3676),
    .Q(\i_seal.sensor_id_reg[1] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _17493_ (.RESET_B(net859),
    .D(net3613),
    .Q(\i_seal.sensor_id_reg[2] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_1 _17494_ (.RESET_B(net857),
    .D(net3646),
    .Q(\i_seal.sensor_id_reg[3] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17495_ (.RESET_B(net441),
    .D(net3648),
    .Q(\i_seal.sensor_id_reg[4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17496_ (.RESET_B(net439),
    .D(net3617),
    .Q(\i_seal.sensor_id_reg[5] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17497_ (.RESET_B(net437),
    .D(net3913),
    .Q(\i_seal.sensor_id_reg[6] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _17498_ (.RESET_B(net407),
    .D(net4038),
    .Q(\i_seal.sensor_id_reg[7] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_2 _17499_ (.RESET_B(net405),
    .D(_01056_),
    .Q(\i_seal.value_reg[0] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17500_ (.RESET_B(net403),
    .D(_01057_),
    .Q(\i_seal.value_reg[1] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_2 _17501_ (.RESET_B(net373),
    .D(_01058_),
    .Q(\i_seal.value_reg[2] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_2 _17502_ (.RESET_B(net371),
    .D(_01059_),
    .Q(\i_seal.value_reg[3] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _17503_ (.RESET_B(net369),
    .D(_01060_),
    .Q(\i_seal.value_reg[4] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_2 _17504_ (.RESET_B(net367),
    .D(_01061_),
    .Q(\i_seal.value_reg[5] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _17505_ (.RESET_B(net365),
    .D(_01062_),
    .Q(\i_seal.value_reg[6] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_2 _17506_ (.RESET_B(net363),
    .D(_01063_),
    .Q(\i_seal.value_reg[7] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _17507_ (.RESET_B(net361),
    .D(_01064_),
    .Q(\i_seal.value_reg[8] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _17508_ (.RESET_B(net359),
    .D(_01065_),
    .Q(\i_seal.value_reg[9] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _17509_ (.RESET_B(net357),
    .D(_01066_),
    .Q(\i_seal.value_reg[10] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _17510_ (.RESET_B(net355),
    .D(_01067_),
    .Q(\i_seal.value_reg[11] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _17511_ (.RESET_B(net353),
    .D(net5096),
    .Q(\i_seal.value_reg[12] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _17512_ (.RESET_B(net351),
    .D(_01069_),
    .Q(\i_seal.value_reg[13] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _17513_ (.RESET_B(net349),
    .D(_01070_),
    .Q(\i_seal.value_reg[14] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _17514_ (.RESET_B(net347),
    .D(_01071_),
    .Q(\i_seal.value_reg[15] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _17515_ (.RESET_B(net345),
    .D(_01072_),
    .Q(\i_seal.value_reg[16] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _17516_ (.RESET_B(net343),
    .D(_01073_),
    .Q(\i_seal.value_reg[17] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _17517_ (.RESET_B(net341),
    .D(_01074_),
    .Q(\i_seal.value_reg[18] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_2 _17518_ (.RESET_B(net339),
    .D(_01075_),
    .Q(\i_seal.value_reg[19] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17519_ (.RESET_B(net337),
    .D(_01076_),
    .Q(\i_seal.value_reg[20] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _17520_ (.RESET_B(net335),
    .D(_01077_),
    .Q(\i_seal.value_reg[21] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _17521_ (.RESET_B(net333),
    .D(_01078_),
    .Q(\i_seal.value_reg[22] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_2 _17522_ (.RESET_B(net331),
    .D(_01079_),
    .Q(\i_seal.value_reg[23] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _17523_ (.RESET_B(net329),
    .D(_01080_),
    .Q(\i_seal.value_reg[24] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17524_ (.RESET_B(net327),
    .D(_01081_),
    .Q(\i_seal.value_reg[25] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17525_ (.RESET_B(net325),
    .D(_01082_),
    .Q(\i_seal.value_reg[26] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17526_ (.RESET_B(net323),
    .D(_01083_),
    .Q(\i_seal.value_reg[27] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_2 _17527_ (.RESET_B(net321),
    .D(_01084_),
    .Q(\i_seal.value_reg[28] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_2 _17528_ (.RESET_B(net319),
    .D(_01085_),
    .Q(\i_seal.value_reg[29] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_2 _17529_ (.RESET_B(net317),
    .D(_01086_),
    .Q(\i_seal.value_reg[30] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_2 _17530_ (.RESET_B(net315),
    .D(_01087_),
    .Q(\i_seal.value_reg[31] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_2 _17531_ (.RESET_B(net313),
    .D(_01088_),
    .Q(\i_seal.state[0] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _17532_ (.RESET_B(net311),
    .D(_01089_),
    .Q(\i_seal.state[1] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _17533_ (.RESET_B(net309),
    .D(_01090_),
    .Q(\i_seal.crc_init ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _17534_ (.RESET_B(net308),
    .D(net3959),
    .Q(\i_seal.crc_byte[0] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _17535_ (.RESET_B(net306),
    .D(net4192),
    .Q(\i_seal.crc_byte[1] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_2 _17536_ (.RESET_B(net304),
    .D(net4304),
    .Q(\i_seal.crc_byte[2] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_2 _17537_ (.RESET_B(net302),
    .D(net4141),
    .Q(\i_seal.crc_byte[3] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_2 _17538_ (.RESET_B(net300),
    .D(net4214),
    .Q(\i_seal.crc_byte[4] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _17539_ (.RESET_B(net298),
    .D(net4244),
    .Q(\i_seal.crc_byte[5] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _17540_ (.RESET_B(net295),
    .D(net4909),
    .Q(\i_seal.crc_byte[6] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _17541_ (.RESET_B(net293),
    .D(net3969),
    .Q(\i_seal.crc_byte[7] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _17542_ (.RESET_B(net291),
    .D(_01099_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[0] ),
    .CLK(net2727));
 sg13g2_dfrbpq_1 _17543_ (.RESET_B(net289),
    .D(_01100_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[1] ),
    .CLK(net2728));
 sg13g2_dfrbpq_1 _17544_ (.RESET_B(net287),
    .D(_01101_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[2] ),
    .CLK(net2729));
 sg13g2_dfrbpq_1 _17545_ (.RESET_B(net285),
    .D(_01102_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[3] ),
    .CLK(net2730));
 sg13g2_dfrbpq_1 _17546_ (.RESET_B(net283),
    .D(_01103_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[4] ),
    .CLK(net2731));
 sg13g2_dfrbpq_1 _17547_ (.RESET_B(net281),
    .D(_01104_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[5] ),
    .CLK(net2732));
 sg13g2_dfrbpq_1 _17548_ (.RESET_B(net279),
    .D(_01105_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[6] ),
    .CLK(net2733));
 sg13g2_dfrbpq_1 _17549_ (.RESET_B(net277),
    .D(_01106_),
    .Q(\i_latch_mem.genblk1[9].l_ram.data_out[7] ),
    .CLK(net2734));
 sg13g2_dfrbpq_1 _17550_ (.RESET_B(net275),
    .D(_01107_),
    .Q(\i_seal.read_seq[0] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17551_ (.RESET_B(net1229),
    .D(_01108_),
    .Q(\i_seal.read_seq[1] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17552_ (.RESET_B(net1230),
    .D(_00000_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .CLK(clknet_leaf_183_clk_regs));
 sg13g2_dfrbpq_1 _17553_ (.RESET_B(net1231),
    .D(_00003_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _17554_ (.RESET_B(net1232),
    .D(_00004_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_1 _17555_ (.RESET_B(net1233),
    .D(_00005_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .CLK(clknet_leaf_186_clk_regs));
 sg13g2_dfrbpq_2 _17556_ (.RESET_B(net1234),
    .D(_00006_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .CLK(clknet_leaf_187_clk_regs));
 sg13g2_dfrbpq_2 _17557_ (.RESET_B(net1235),
    .D(_00007_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .CLK(clknet_leaf_193_clk_regs));
 sg13g2_dfrbpq_1 _17558_ (.RESET_B(net1236),
    .D(_00008_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _17559_ (.RESET_B(net1237),
    .D(_00009_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _17560_ (.RESET_B(net1238),
    .D(_00010_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _17561_ (.RESET_B(net1239),
    .D(_00011_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _17562_ (.RESET_B(net1336),
    .D(_00001_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _17563_ (.RESET_B(net273),
    .D(_00002_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .CLK(clknet_leaf_194_clk_regs));
 sg13g2_dfrbpq_1 _17564_ (.RESET_B(net271),
    .D(_01109_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_1 _17565_ (.RESET_B(net270),
    .D(_01110_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_2 _17566_ (.RESET_B(net269),
    .D(net4569),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_1 _17567_ (.RESET_B(net268),
    .D(net4417),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_2 _17568_ (.RESET_B(net267),
    .D(net3683),
    .Q(\i_tinyqv.cpu.i_core.mepc[0] ),
    .CLK(clknet_leaf_179_clk_regs));
 sg13g2_dfrbpq_2 _17569_ (.RESET_B(net266),
    .D(net4439),
    .Q(\i_tinyqv.cpu.i_core.mepc[1] ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_2 _17570_ (.RESET_B(net265),
    .D(_01115_),
    .Q(\i_tinyqv.cpu.i_core.mepc[2] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_2 _17571_ (.RESET_B(net264),
    .D(_01116_),
    .Q(\i_tinyqv.cpu.i_core.mepc[3] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_1 _17572_ (.RESET_B(net263),
    .D(_01117_),
    .Q(\i_tinyqv.cpu.i_core.mepc[4] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_1 _17573_ (.RESET_B(net262),
    .D(_01118_),
    .Q(\i_tinyqv.cpu.i_core.mepc[5] ),
    .CLK(clknet_leaf_188_clk_regs));
 sg13g2_dfrbpq_1 _17574_ (.RESET_B(net261),
    .D(net4511),
    .Q(\i_tinyqv.cpu.i_core.mepc[6] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_1 _17575_ (.RESET_B(net260),
    .D(_01120_),
    .Q(\i_tinyqv.cpu.i_core.mepc[7] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_1 _17576_ (.RESET_B(net259),
    .D(net4411),
    .Q(\i_tinyqv.cpu.i_core.mepc[8] ),
    .CLK(clknet_leaf_189_clk_regs));
 sg13g2_dfrbpq_1 _17577_ (.RESET_B(net257),
    .D(_01122_),
    .Q(\i_tinyqv.cpu.i_core.mepc[9] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_1 _17578_ (.RESET_B(net255),
    .D(net4589),
    .Q(\i_tinyqv.cpu.i_core.mepc[10] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_1 _17579_ (.RESET_B(net253),
    .D(net4405),
    .Q(\i_tinyqv.cpu.i_core.mepc[11] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_1 _17580_ (.RESET_B(net251),
    .D(net4643),
    .Q(\i_tinyqv.cpu.i_core.mepc[12] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_1 _17581_ (.RESET_B(net249),
    .D(_01126_),
    .Q(\i_tinyqv.cpu.i_core.mepc[13] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_1 _17582_ (.RESET_B(net247),
    .D(net4414),
    .Q(\i_tinyqv.cpu.i_core.mepc[14] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _17583_ (.RESET_B(net245),
    .D(_01128_),
    .Q(\i_tinyqv.cpu.i_core.mepc[15] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_1 _17584_ (.RESET_B(net243),
    .D(_01129_),
    .Q(\i_tinyqv.cpu.i_core.mepc[16] ),
    .CLK(clknet_leaf_190_clk_regs));
 sg13g2_dfrbpq_1 _17585_ (.RESET_B(net241),
    .D(net4004),
    .Q(\i_tinyqv.cpu.i_core.mepc[17] ),
    .CLK(clknet_leaf_191_clk_regs));
 sg13g2_dfrbpq_1 _17586_ (.RESET_B(net239),
    .D(net3953),
    .Q(\i_tinyqv.cpu.i_core.mepc[18] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _17587_ (.RESET_B(net237),
    .D(net4297),
    .Q(\i_tinyqv.cpu.i_core.mepc[19] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _17588_ (.RESET_B(net235),
    .D(net4585),
    .Q(\i_tinyqv.cpu.instr_data[0][2] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17589_ (.RESET_B(net233),
    .D(net3985),
    .Q(\i_tinyqv.cpu.instr_data[0][3] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _17590_ (.RESET_B(net231),
    .D(net4558),
    .Q(\i_tinyqv.cpu.instr_data[0][4] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _17591_ (.RESET_B(net229),
    .D(net4504),
    .Q(\i_tinyqv.cpu.instr_data[0][5] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _17592_ (.RESET_B(net227),
    .D(net4658),
    .Q(\i_tinyqv.cpu.instr_data[0][6] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _17593_ (.RESET_B(net224),
    .D(net4499),
    .Q(\i_tinyqv.cpu.instr_data[0][7] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17594_ (.RESET_B(net222),
    .D(net4210),
    .Q(\i_tinyqv.cpu.instr_data[0][8] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17595_ (.RESET_B(net220),
    .D(net4453),
    .Q(\i_tinyqv.cpu.instr_data[0][9] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _17596_ (.RESET_B(net218),
    .D(net4583),
    .Q(\i_tinyqv.cpu.instr_data[0][10] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17597_ (.RESET_B(net216),
    .D(net4497),
    .Q(\i_tinyqv.cpu.instr_data[0][11] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _17598_ (.RESET_B(net214),
    .D(net4455),
    .Q(\i_tinyqv.cpu.instr_data[0][12] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _17599_ (.RESET_B(net212),
    .D(net4506),
    .Q(\i_tinyqv.cpu.instr_data[0][13] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _17600_ (.RESET_B(net210),
    .D(net4571),
    .Q(\i_tinyqv.cpu.instr_data[0][14] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _17601_ (.RESET_B(net208),
    .D(net4493),
    .Q(\i_tinyqv.cpu.instr_data[0][15] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _17602_ (.RESET_B(net206),
    .D(_01147_),
    .Q(\i_tinyqv.cpu.instr_write_offset[1] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17603_ (.RESET_B(net204),
    .D(_01148_),
    .Q(\i_tinyqv.cpu.instr_write_offset[2] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _17604_ (.RESET_B(net202),
    .D(_01149_),
    .Q(\addr[24] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _17605_ (.RESET_B(net198),
    .D(_01150_),
    .Q(\addr[25] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _17606_ (.RESET_B(net194),
    .D(_01151_),
    .Q(\addr[26] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _17607_ (.RESET_B(net190),
    .D(_01152_),
    .Q(\addr[27] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_2 _17608_ (.RESET_B(net186),
    .D(net5248),
    .Q(\addr[0] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _17609_ (.RESET_B(net184),
    .D(_01154_),
    .Q(\addr[1] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _17610_ (.RESET_B(net182),
    .D(_01155_),
    .Q(\addr[2] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _17611_ (.RESET_B(net180),
    .D(_01156_),
    .Q(\addr[3] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17612_ (.RESET_B(net178),
    .D(_01157_),
    .Q(\addr[4] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _17613_ (.RESET_B(net176),
    .D(net5264),
    .Q(\addr[5] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17614_ (.RESET_B(net174),
    .D(_01159_),
    .Q(\addr[6] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _17615_ (.RESET_B(net172),
    .D(net4233),
    .Q(\addr[7] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17616_ (.RESET_B(net170),
    .D(net4235),
    .Q(\addr[8] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17617_ (.RESET_B(net168),
    .D(net4343),
    .Q(\addr[9] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _17618_ (.RESET_B(net166),
    .D(net4117),
    .Q(\addr[10] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _17619_ (.RESET_B(net164),
    .D(net4226),
    .Q(\addr[11] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _17620_ (.RESET_B(net162),
    .D(net4631),
    .Q(\addr[12] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17621_ (.RESET_B(net160),
    .D(net4186),
    .Q(\addr[13] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _17622_ (.RESET_B(net158),
    .D(net4401),
    .Q(\addr[14] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _17623_ (.RESET_B(net152),
    .D(net4532),
    .Q(\addr[15] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17624_ (.RESET_B(net150),
    .D(net4660),
    .Q(\addr[16] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _17625_ (.RESET_B(net148),
    .D(_01170_),
    .Q(\addr[17] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _17626_ (.RESET_B(net146),
    .D(net4302),
    .Q(\addr[18] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _17627_ (.RESET_B(net144),
    .D(net4579),
    .Q(\addr[19] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _17628_ (.RESET_B(net142),
    .D(net4780),
    .Q(\addr[20] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17629_ (.RESET_B(net140),
    .D(_01174_),
    .Q(\addr[21] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17630_ (.RESET_B(net138),
    .D(net4300),
    .Q(\addr[22] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _17631_ (.RESET_B(net136),
    .D(_01176_),
    .Q(\addr[23] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17632_ (.RESET_B(net134),
    .D(net3630),
    .Q(\i_spi.data[1] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _17633_ (.RESET_B(net132),
    .D(_01178_),
    .Q(\i_spi.data[2] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17634_ (.RESET_B(net130),
    .D(net3671),
    .Q(\i_spi.data[3] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17635_ (.RESET_B(net128),
    .D(net3644),
    .Q(\i_spi.data[4] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _17636_ (.RESET_B(net126),
    .D(net3660),
    .Q(\i_spi.data[5] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _17637_ (.RESET_B(net124),
    .D(net3851),
    .Q(\i_spi.data[6] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _17638_ (.RESET_B(net122),
    .D(net3717),
    .Q(\i_spi.data[7] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17639_ (.RESET_B(net119),
    .D(_01184_),
    .Q(\i_latch_mem.cycle[0] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _17640_ (.RESET_B(net117),
    .D(net4279),
    .Q(\i_crc16.bit_cnt[3] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _17641_ (.RESET_B(net113),
    .D(net4546),
    .Q(\i_tinyqv.cpu.instr_data[2][2] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17642_ (.RESET_B(net111),
    .D(net3637),
    .Q(\i_tinyqv.cpu.instr_data[2][3] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17643_ (.RESET_B(net109),
    .D(net4591),
    .Q(\i_tinyqv.cpu.instr_data[2][4] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _17644_ (.RESET_B(net107),
    .D(net4519),
    .Q(\i_tinyqv.cpu.instr_data[2][5] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _17645_ (.RESET_B(net105),
    .D(net4622),
    .Q(\i_tinyqv.cpu.instr_data[2][6] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _17646_ (.RESET_B(net103),
    .D(net4575),
    .Q(\i_tinyqv.cpu.instr_data[2][7] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17647_ (.RESET_B(net101),
    .D(net3694),
    .Q(\i_tinyqv.cpu.instr_data[2][8] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17648_ (.RESET_B(net99),
    .D(net4474),
    .Q(\i_tinyqv.cpu.instr_data[2][9] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17649_ (.RESET_B(net97),
    .D(net4669),
    .Q(\i_tinyqv.cpu.instr_data[2][10] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17650_ (.RESET_B(net95),
    .D(net4524),
    .Q(\i_tinyqv.cpu.instr_data[2][11] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17651_ (.RESET_B(net93),
    .D(net4645),
    .Q(\i_tinyqv.cpu.instr_data[2][12] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _17652_ (.RESET_B(net91),
    .D(net4602),
    .Q(\i_tinyqv.cpu.instr_data[2][13] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _17653_ (.RESET_B(net88),
    .D(net4459),
    .Q(\i_tinyqv.cpu.instr_data[2][14] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _17654_ (.RESET_B(net86),
    .D(net4526),
    .Q(\i_tinyqv.cpu.instr_data[2][15] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _17655_ (.RESET_B(net83),
    .D(net3842),
    .Q(\i_tinyqv.cpu.instr_data[3][0] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _17656_ (.RESET_B(net81),
    .D(net4050),
    .Q(\i_tinyqv.cpu.instr_data[3][1] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _17657_ (.RESET_B(net79),
    .D(_01202_),
    .Q(\i_i2c_peri.i_i2c.busy_reg ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _17658_ (.RESET_B(net77),
    .D(net4824),
    .Q(\i_i2c_peri.i_i2c.sda_o_reg ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _17659_ (.RESET_B(net1374),
    .D(net4446),
    .Q(\i_i2c_peri.i_i2c.scl_o_reg ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _17660_ (.RESET_B(net73),
    .D(net3317),
    .Q(\i_i2c_peri.i_i2c.sda_i_reg ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17661_ (.RESET_B(net69),
    .D(net4162),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[0] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _17662_ (.RESET_B(net67),
    .D(net4340),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[1] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _17663_ (.RESET_B(net65),
    .D(net3949),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[2] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_2 _17664_ (.RESET_B(net44),
    .D(net4262),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[3] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _17665_ (.RESET_B(net38),
    .D(net4208),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[4] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _17666_ (.RESET_B(net36),
    .D(net4109),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[5] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _17667_ (.RESET_B(net2708),
    .D(net4058),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[6] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17668_ (.RESET_B(net2701),
    .D(net3832),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[7] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17669_ (.RESET_B(net2699),
    .D(net3410),
    .Q(\i_i2c_peri.i_i2c.delay_sda_reg ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _17670_ (.RESET_B(net2695),
    .D(_01214_),
    .Q(\i_i2c_peri.i_i2c.phy_rx_data_reg ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _17671_ (.RESET_B(net2693),
    .D(net3633),
    .Q(\i_i2c_peri.i_i2c.bus_active_reg ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_2 _17672_ (.RESET_B(net2688),
    .D(net3989),
    .Q(\i_i2c_peri.i_i2c.mode_stop_reg ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _17673_ (.RESET_B(net1772),
    .D(_01217_),
    .Q(\i_i2c_peri.sda_sync[0] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _17674_ (.RESET_B(net1770),
    .D(_01218_),
    .Q(\i_i2c_peri.i_i2c.sda_i ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17675_ (.RESET_B(net1768),
    .D(net4166),
    .Q(\i_i2c_peri.i_i2c.last_reg ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _17676_ (.RESET_B(net1766),
    .D(_01220_),
    .Q(\i_i2c_peri.i_i2c.m_axis_data_tvalid_reg ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _17677_ (.RESET_B(net1764),
    .D(_01221_),
    .Q(\i_i2c_peri.i_i2c.delay_reg[0] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _17678_ (.RESET_B(net1760),
    .D(net4936),
    .Q(\i_i2c_peri.i_i2c.delay_reg[1] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _17679_ (.RESET_B(net1740),
    .D(net4886),
    .Q(\i_i2c_peri.i_i2c.delay_reg[2] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _17680_ (.RESET_B(net1705),
    .D(net4761),
    .Q(\i_i2c_peri.i_i2c.delay_reg[3] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _17681_ (.RESET_B(net1701),
    .D(net4696),
    .Q(\i_i2c_peri.i_i2c.delay_reg[4] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _17682_ (.RESET_B(net1697),
    .D(net4872),
    .Q(\i_i2c_peri.i_i2c.delay_reg[5] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _17683_ (.RESET_B(net1693),
    .D(_01227_),
    .Q(\i_i2c_peri.i_i2c.delay_reg[6] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _17684_ (.RESET_B(net1689),
    .D(net4247),
    .Q(\i_i2c_peri.i_i2c.delay_reg[7] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _17685_ (.RESET_B(net1685),
    .D(net4701),
    .Q(\i_i2c_peri.i_i2c.delay_reg[8] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _17686_ (.RESET_B(net1681),
    .D(net4620),
    .Q(\i_i2c_peri.i_i2c.delay_reg[9] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _17687_ (.RESET_B(net1677),
    .D(_01231_),
    .Q(\i_i2c_peri.i_i2c.delay_reg[10] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _17688_ (.RESET_B(net1673),
    .D(net4900),
    .Q(\i_i2c_peri.i_i2c.delay_reg[11] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _17689_ (.RESET_B(net1669),
    .D(net4074),
    .Q(\i_i2c_peri.i_i2c.delay_reg[12] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _17690_ (.RESET_B(net1665),
    .D(_01234_),
    .Q(\i_i2c_peri.i_i2c.delay_reg[13] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _17691_ (.RESET_B(net1661),
    .D(_01235_),
    .Q(\i_i2c_peri.i_i2c.delay_reg[14] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _17692_ (.RESET_B(net1657),
    .D(net4925),
    .Q(\i_i2c_peri.i_i2c.delay_reg[15] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _17693_ (.RESET_B(net1653),
    .D(net4184),
    .Q(\i_i2c_peri.i_i2c.delay_reg[16] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _17694_ (.RESET_B(net1649),
    .D(net5161),
    .Q(\i_i2c_peri.i_i2c.phy_state_reg[0] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _17695_ (.RESET_B(net1645),
    .D(_01239_),
    .Q(\i_i2c_peri.i_i2c.phy_state_reg[1] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _17696_ (.RESET_B(net1641),
    .D(_01240_),
    .Q(\i_i2c_peri.i_i2c.phy_state_reg[2] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _17697_ (.RESET_B(net1774),
    .D(net5351),
    .Q(\i_i2c_peri.i_i2c.phy_state_reg[3] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _17698_ (.RESET_B(net1637),
    .D(net3397),
    .Q(\i_i2c_peri.i_i2c.last_sda_i_reg ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17699_ (.RESET_B(net1633),
    .D(net3651),
    .Q(\i_i2c_peri.i_i2c.mode_write_multiple_reg ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _17700_ (.RESET_B(net1631),
    .D(_01243_),
    .Q(\i_i2c_peri.i_i2c.addr_reg[0] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _17701_ (.RESET_B(net1629),
    .D(_01244_),
    .Q(\i_i2c_peri.i_i2c.addr_reg[1] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _17702_ (.RESET_B(net1627),
    .D(net4242),
    .Q(\i_i2c_peri.i_i2c.addr_reg[2] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _17703_ (.RESET_B(net1625),
    .D(net4128),
    .Q(\i_i2c_peri.i_i2c.addr_reg[3] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _17704_ (.RESET_B(net1623),
    .D(net4069),
    .Q(\i_i2c_peri.i_i2c.addr_reg[4] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _17705_ (.RESET_B(net1621),
    .D(net4249),
    .Q(\i_i2c_peri.i_i2c.addr_reg[5] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _17706_ (.RESET_B(net1619),
    .D(_01249_),
    .Q(\i_i2c_peri.i_i2c.addr_reg[6] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _17707_ (.RESET_B(net1617),
    .D(net4567),
    .Q(\i_i2c_peri.i_i2c.mode_read_reg ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _17708_ (.RESET_B(net1615),
    .D(_01251_),
    .Q(\i_i2c_peri.i_i2c.delay_scl_reg ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _17709_ (.RESET_B(net1613),
    .D(net3480),
    .Q(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _17710_ (.RESET_B(net1609),
    .D(net4550),
    .Q(\i_tinyqv.cpu.instr_data[3][2] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17711_ (.RESET_B(net1607),
    .D(net3730),
    .Q(\i_tinyqv.cpu.instr_data[3][3] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17712_ (.RESET_B(net1605),
    .D(net4667),
    .Q(\i_tinyqv.cpu.instr_data[3][4] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _17713_ (.RESET_B(net1603),
    .D(net4449),
    .Q(\i_tinyqv.cpu.instr_data[3][5] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _17714_ (.RESET_B(net1601),
    .D(net4495),
    .Q(\i_tinyqv.cpu.instr_data[3][6] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _17715_ (.RESET_B(net1599),
    .D(net4428),
    .Q(\i_tinyqv.cpu.instr_data[3][7] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17716_ (.RESET_B(net1597),
    .D(net3803),
    .Q(\i_tinyqv.cpu.instr_data[3][8] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17717_ (.RESET_B(net1595),
    .D(net4408),
    .Q(\i_tinyqv.cpu.instr_data[3][9] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _17718_ (.RESET_B(net1593),
    .D(net4662),
    .Q(\i_tinyqv.cpu.instr_data[3][10] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17719_ (.RESET_B(net1591),
    .D(net4425),
    .Q(\i_tinyqv.cpu.instr_data[3][11] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _17720_ (.RESET_B(net1589),
    .D(net4488),
    .Q(\i_tinyqv.cpu.instr_data[3][12] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _17721_ (.RESET_B(net1587),
    .D(net4617),
    .Q(\i_tinyqv.cpu.instr_data[3][13] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _17722_ (.RESET_B(net1585),
    .D(net4548),
    .Q(\i_tinyqv.cpu.instr_data[3][14] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _17723_ (.RESET_B(net1583),
    .D(net4635),
    .Q(\i_tinyqv.cpu.instr_data[3][15] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _17724_ (.RESET_B(net1581),
    .D(net4652),
    .Q(\i2c_config_out[0] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17725_ (.RESET_B(net1577),
    .D(net4370),
    .Q(\i2c_config_out[1] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17726_ (.RESET_B(net1573),
    .D(net4955),
    .Q(\i2c_config_out[2] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _17727_ (.RESET_B(net1569),
    .D(net4806),
    .Q(\i2c_config_out[3] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _17728_ (.RESET_B(net1565),
    .D(_01271_),
    .Q(\i2c_config_out[4] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _17729_ (.RESET_B(net1557),
    .D(_01272_),
    .Q(\i2c_config_out[5] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _17730_ (.RESET_B(net1553),
    .D(_01273_),
    .Q(\i2c_config_out[6] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _17731_ (.RESET_B(net1549),
    .D(_01274_),
    .Q(\i2c_config_out[7] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _17732_ (.RESET_B(net1545),
    .D(_01275_),
    .Q(\i2c_config_out[8] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _17733_ (.RESET_B(net1541),
    .D(_01276_),
    .Q(\i2c_config_out[9] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17734_ (.RESET_B(net1537),
    .D(_01277_),
    .Q(\i2c_config_out[10] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17735_ (.RESET_B(net1486),
    .D(net5003),
    .Q(\i2c_config_out[11] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17736_ (.RESET_B(net1482),
    .D(net5127),
    .Q(\i2c_config_out[12] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17737_ (.RESET_B(net1478),
    .D(_01280_),
    .Q(\i2c_config_out[13] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17738_ (.RESET_B(net1462),
    .D(_01281_),
    .Q(\i2c_config_out[14] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17739_ (.RESET_B(net1458),
    .D(_01282_),
    .Q(\i2c_config_out[15] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _17740_ (.RESET_B(net1454),
    .D(_01283_),
    .Q(\i_i2c_peri.addr_latch[0] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _17741_ (.RESET_B(net1450),
    .D(_01284_),
    .Q(\i_i2c_peri.addr_latch[1] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17742_ (.RESET_B(net1445),
    .D(_01285_),
    .Q(\i_i2c_peri.addr_latch[2] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _17743_ (.RESET_B(net1441),
    .D(_01286_),
    .Q(\i_i2c_peri.addr_latch[3] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _17744_ (.RESET_B(net1437),
    .D(_01287_),
    .Q(\i_i2c_peri.addr_latch[4] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _17745_ (.RESET_B(net1432),
    .D(_01288_),
    .Q(\i_i2c_peri.addr_latch[5] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _17746_ (.RESET_B(net1428),
    .D(_01289_),
    .Q(\i_i2c_peri.addr_latch[6] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _17747_ (.RESET_B(net1422),
    .D(net4056),
    .Q(\i_i2c_peri.cmd_stop_reg ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _17748_ (.RESET_B(net1418),
    .D(_01291_),
    .Q(\i_i2c_peri.cmd_write_m_reg ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _17749_ (.RESET_B(net1414),
    .D(net4724),
    .Q(\i_i2c_peri.cmd_read_reg ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _17750_ (.RESET_B(net1386),
    .D(_01293_),
    .Q(\i_i2c_peri.cmd_start_reg ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _17751_ (.RESET_B(net1382),
    .D(net3752),
    .Q(\i_i2c_peri.cmd_addr_reg[0] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _17752_ (.RESET_B(net1378),
    .D(net4224),
    .Q(\i_i2c_peri.cmd_addr_reg[1] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _17753_ (.RESET_B(net1373),
    .D(net4360),
    .Q(\i_i2c_peri.cmd_addr_reg[2] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _17754_ (.RESET_B(net1369),
    .D(net4332),
    .Q(\i_i2c_peri.cmd_addr_reg[3] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _17755_ (.RESET_B(net1365),
    .D(_01298_),
    .Q(\i_i2c_peri.cmd_addr_reg[4] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _17756_ (.RESET_B(net1361),
    .D(net4259),
    .Q(\i_i2c_peri.cmd_addr_reg[5] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _17757_ (.RESET_B(net1357),
    .D(net3801),
    .Q(\i_i2c_peri.cmd_addr_reg[6] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _17758_ (.RESET_B(net1353),
    .D(_01301_),
    .Q(\i_i2c_peri.cmd_pending ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _17759_ (.RESET_B(net1349),
    .D(net4613),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tlast ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _17760_ (.RESET_B(net1345),
    .D(_01303_),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[0] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _17761_ (.RESET_B(net1341),
    .D(_01304_),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[1] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _17762_ (.RESET_B(net1337),
    .D(net4726),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[2] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _17763_ (.RESET_B(net1332),
    .D(_01306_),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[3] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _17764_ (.RESET_B(net1328),
    .D(net4750),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[4] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _17765_ (.RESET_B(net1324),
    .D(net4813),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[5] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _17766_ (.RESET_B(net1320),
    .D(net4508),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[6] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _17767_ (.RESET_B(net1316),
    .D(net4461),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tdata[7] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _17768_ (.RESET_B(net1312),
    .D(_01311_),
    .Q(\i_i2c_peri.tx_pending ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _17769_ (.RESET_B(net1308),
    .D(net4272),
    .Q(\i_i2c_peri.rx_has_data ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _17770_ (.RESET_B(net1304),
    .D(_01313_),
    .Q(\i2c_data_out[0] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _17771_ (.RESET_B(net1299),
    .D(net4027),
    .Q(\i2c_data_out[1] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _17772_ (.RESET_B(net1295),
    .D(_01315_),
    .Q(\i2c_data_out[2] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_2 _17773_ (.RESET_B(net1291),
    .D(net4065),
    .Q(\i2c_data_out[3] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _17774_ (.RESET_B(net1287),
    .D(net4113),
    .Q(\i2c_data_out[4] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _17775_ (.RESET_B(net1283),
    .D(net3975),
    .Q(\i2c_data_out[5] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _17776_ (.RESET_B(net1279),
    .D(_01319_),
    .Q(\i2c_data_out[6] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _17777_ (.RESET_B(net1275),
    .D(net4204),
    .Q(\i2c_data_out[7] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _17778_ (.RESET_B(net1271),
    .D(_01321_),
    .Q(\i2c_data_out[8] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17779_ (.RESET_B(net1267),
    .D(net4833),
    .Q(\crc16_read[0] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17780_ (.RESET_B(net1263),
    .D(net4875),
    .Q(\crc16_read[1] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _17781_ (.RESET_B(net1259),
    .D(_01324_),
    .Q(\crc16_read[2] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17782_ (.RESET_B(net1255),
    .D(_01325_),
    .Q(\crc16_read[3] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17783_ (.RESET_B(net1251),
    .D(net5014),
    .Q(\crc16_read[4] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _17784_ (.RESET_B(net1247),
    .D(net4993),
    .Q(\crc16_read[5] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _17785_ (.RESET_B(net1243),
    .D(net4991),
    .Q(\crc16_read[6] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _17786_ (.RESET_B(net1227),
    .D(_01329_),
    .Q(\crc16_read[7] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _17787_ (.RESET_B(net1223),
    .D(_01330_),
    .Q(\i_uart_tx.data_to_send[0] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17788_ (.RESET_B(net1219),
    .D(_01331_),
    .Q(\i_uart_tx.data_to_send[1] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17789_ (.RESET_B(net1215),
    .D(_01332_),
    .Q(\i_uart_tx.data_to_send[2] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _17790_ (.RESET_B(net1211),
    .D(net4849),
    .Q(\i_uart_tx.data_to_send[3] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17791_ (.RESET_B(net1207),
    .D(net4794),
    .Q(\i_uart_tx.data_to_send[4] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17792_ (.RESET_B(net1203),
    .D(net4815),
    .Q(\i_uart_tx.data_to_send[5] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17793_ (.RESET_B(net1199),
    .D(net4709),
    .Q(\i_uart_tx.data_to_send[6] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17794_ (.RESET_B(net1195),
    .D(net3592),
    .Q(\i_uart_tx.data_to_send[7] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17795_ (.RESET_B(net1191),
    .D(net4356),
    .Q(\i_uart_tx.cycle_counter[0] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _17796_ (.RESET_B(net1187),
    .D(_01339_),
    .Q(\i_uart_tx.cycle_counter[1] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _17797_ (.RESET_B(net1182),
    .D(net3908),
    .Q(\i_uart_tx.cycle_counter[2] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _17798_ (.RESET_B(net1178),
    .D(net4677),
    .Q(\i_uart_tx.cycle_counter[3] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _17799_ (.RESET_B(net1174),
    .D(net4648),
    .Q(\i_uart_tx.cycle_counter[4] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _17800_ (.RESET_B(net1170),
    .D(_01343_),
    .Q(\i_uart_tx.cycle_counter[5] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _17801_ (.RESET_B(net1166),
    .D(net4468),
    .Q(\i_uart_tx.cycle_counter[6] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _17802_ (.RESET_B(net1162),
    .D(net3997),
    .Q(\i_uart_tx.cycle_counter[7] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _17803_ (.RESET_B(net1158),
    .D(_01346_),
    .Q(\i_uart_tx.cycle_counter[8] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _17804_ (.RESET_B(net1154),
    .D(_01347_),
    .Q(\i_uart_tx.fsm_state[0] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _17805_ (.RESET_B(net1150),
    .D(net4022),
    .Q(\i_uart_tx.fsm_state[1] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _17806_ (.RESET_B(net1146),
    .D(net4763),
    .Q(\i_uart_tx.fsm_state[2] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _17807_ (.RESET_B(net1142),
    .D(net4716),
    .Q(\i_uart_tx.fsm_state[3] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17808_ (.RESET_B(net1138),
    .D(net4194),
    .Q(\i_uart_rx.recieved_data[0] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _17809_ (.RESET_B(net1136),
    .D(net4698),
    .Q(\i_uart_rx.recieved_data[1] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17810_ (.RESET_B(net1134),
    .D(_01353_),
    .Q(\i_uart_rx.recieved_data[2] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17811_ (.RESET_B(net1132),
    .D(_01354_),
    .Q(\i_uart_rx.recieved_data[3] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17812_ (.RESET_B(net1130),
    .D(_01355_),
    .Q(\i_uart_rx.recieved_data[4] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17813_ (.RESET_B(net1128),
    .D(net4732),
    .Q(\i_uart_rx.recieved_data[5] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _17814_ (.RESET_B(net1126),
    .D(_01357_),
    .Q(\i_uart_rx.recieved_data[6] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17815_ (.RESET_B(net1124),
    .D(_01358_),
    .Q(\i_uart_rx.recieved_data[7] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _17816_ (.RESET_B(net1122),
    .D(_01359_),
    .Q(\i_uart_rx.cycle_counter[0] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _17817_ (.RESET_B(net1120),
    .D(_01360_),
    .Q(\i_uart_rx.cycle_counter[1] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_2 _17818_ (.RESET_B(net1118),
    .D(_01361_),
    .Q(\i_uart_rx.cycle_counter[2] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _17819_ (.RESET_B(net1116),
    .D(net3813),
    .Q(\i_uart_rx.cycle_counter[3] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _17820_ (.RESET_B(net1114),
    .D(_01363_),
    .Q(\i_uart_rx.cycle_counter[4] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _17821_ (.RESET_B(net1112),
    .D(_01364_),
    .Q(\i_uart_rx.cycle_counter[5] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _17822_ (.RESET_B(net1110),
    .D(net3820),
    .Q(\i_uart_rx.cycle_counter[6] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_2 _17823_ (.RESET_B(net1108),
    .D(_01366_),
    .Q(\i_uart_rx.cycle_counter[7] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _17824_ (.RESET_B(net1106),
    .D(_01367_),
    .Q(\i_uart_rx.cycle_counter[8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _17825_ (.RESET_B(net1104),
    .D(net4046),
    .Q(\i_uart_rx.bit_sample ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _17826_ (.RESET_B(net1100),
    .D(_01369_),
    .Q(\i_uart_rx.rxd_reg[0] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _17827_ (.RESET_B(net1098),
    .D(_01370_),
    .Q(\i_uart_rx.rxd_reg[1] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _17828_ (.RESET_B(net1096),
    .D(_01371_),
    .Q(\i_uart_rx.fsm_state[0] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _17829_ (.RESET_B(net1092),
    .D(_01372_),
    .Q(\i_uart_rx.fsm_state[1] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_2 _17830_ (.RESET_B(net1088),
    .D(net4788),
    .Q(\i_uart_rx.fsm_state[2] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_2 _17831_ (.RESET_B(net1084),
    .D(net5238),
    .Q(\i_uart_rx.fsm_state[3] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _17832_ (.RESET_B(net1080),
    .D(_01375_),
    .Q(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _17833_ (.RESET_B(net1078),
    .D(net3773),
    .Q(\i_tinyqv.cpu.instr_data[0][0] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _17834_ (.RESET_B(net1074),
    .D(net3808),
    .Q(\i_tinyqv.cpu.instr_data[0][1] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _17835_ (.RESET_B(net1070),
    .D(net3543),
    .Q(\i_spi.end_txn_reg ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _17836_ (.RESET_B(net1068),
    .D(net4741),
    .Q(\i_spi.clock_count[0] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _17837_ (.RESET_B(net1064),
    .D(net3621),
    .Q(\i_spi.clock_count[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _17838_ (.RESET_B(net1060),
    .D(_01381_),
    .Q(\i_spi.clock_count[2] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _17839_ (.RESET_B(net1056),
    .D(_01382_),
    .Q(\i_spi.clock_count[3] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _17840_ (.RESET_B(net1052),
    .D(_01383_),
    .Q(\i_spi.data[0] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _17841_ (.RESET_B(net1050),
    .D(net4231),
    .Q(\i_spi.bits_remaining[0] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _17842_ (.RESET_B(net1046),
    .D(_01385_),
    .Q(\i_spi.bits_remaining[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _17843_ (.RESET_B(net1042),
    .D(net4605),
    .Q(\i_spi.bits_remaining[2] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _17844_ (.RESET_B(net1038),
    .D(net4201),
    .Q(\i_spi.bits_remaining[3] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _17845_ (.RESET_B(net1034),
    .D(_01388_),
    .Q(\i_spi.busy ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _17846_ (.RESET_B(net1032),
    .D(net4252),
    .Q(\i_spi.spi_select ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _17847_ (.RESET_B(net1028),
    .D(_01390_),
    .Q(\i_seal.commit_dropped ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17848_ (.RESET_B(net1026),
    .D(_01391_),
    .Q(\i_spi.spi_clk_out ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _17849_ (.RESET_B(net1022),
    .D(_01392_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[0] ),
    .CLK(net2735));
 sg13g2_dfrbpq_1 _17850_ (.RESET_B(net1018),
    .D(_01393_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[1] ),
    .CLK(net2736));
 sg13g2_dfrbpq_1 _17851_ (.RESET_B(net1014),
    .D(_01394_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[2] ),
    .CLK(net2737));
 sg13g2_dfrbpq_1 _17852_ (.RESET_B(net1010),
    .D(_01395_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[3] ),
    .CLK(net2738));
 sg13g2_dfrbpq_1 _17853_ (.RESET_B(net1006),
    .D(_01396_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[4] ),
    .CLK(net2739));
 sg13g2_dfrbpq_1 _17854_ (.RESET_B(net1002),
    .D(_01397_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[5] ),
    .CLK(net2740));
 sg13g2_dfrbpq_1 _17855_ (.RESET_B(net998),
    .D(_01398_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[6] ),
    .CLK(net2741));
 sg13g2_dfrbpq_1 _17856_ (.RESET_B(net994),
    .D(_01399_),
    .Q(\i_latch_mem.genblk1[30].l_ram.data_out[7] ),
    .CLK(net2742));
 sg13g2_dfrbpq_1 _17857_ (.RESET_B(net990),
    .D(_01400_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[0] ),
    .CLK(net2743));
 sg13g2_dfrbpq_1 _17858_ (.RESET_B(net986),
    .D(_01401_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[1] ),
    .CLK(net2744));
 sg13g2_dfrbpq_1 _17859_ (.RESET_B(net982),
    .D(_01402_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[2] ),
    .CLK(net2745));
 sg13g2_dfrbpq_1 _17860_ (.RESET_B(net978),
    .D(_01403_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[3] ),
    .CLK(net2746));
 sg13g2_dfrbpq_1 _17861_ (.RESET_B(net974),
    .D(_01404_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[4] ),
    .CLK(net2747));
 sg13g2_dfrbpq_1 _17862_ (.RESET_B(net970),
    .D(_01405_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[5] ),
    .CLK(net2748));
 sg13g2_dfrbpq_1 _17863_ (.RESET_B(net966),
    .D(_01406_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[6] ),
    .CLK(net2749));
 sg13g2_dfrbpq_1 _17864_ (.RESET_B(net962),
    .D(_01407_),
    .Q(\i_latch_mem.genblk1[2].l_ram.data_out[7] ),
    .CLK(net2750));
 sg13g2_dfrbpq_1 _17865_ (.RESET_B(net958),
    .D(_01408_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[0] ),
    .CLK(net2751));
 sg13g2_dfrbpq_1 _17866_ (.RESET_B(net954),
    .D(_01409_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[1] ),
    .CLK(net2752));
 sg13g2_dfrbpq_1 _17867_ (.RESET_B(net950),
    .D(_01410_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[2] ),
    .CLK(net2753));
 sg13g2_dfrbpq_1 _17868_ (.RESET_B(net946),
    .D(_01411_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[3] ),
    .CLK(net2754));
 sg13g2_dfrbpq_1 _17869_ (.RESET_B(net942),
    .D(_01412_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[4] ),
    .CLK(net2755));
 sg13g2_dfrbpq_1 _17870_ (.RESET_B(net938),
    .D(_01413_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[5] ),
    .CLK(net2756));
 sg13g2_dfrbpq_1 _17871_ (.RESET_B(net934),
    .D(_01414_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[6] ),
    .CLK(net2757));
 sg13g2_dfrbpq_1 _17872_ (.RESET_B(net930),
    .D(_01415_),
    .Q(\i_latch_mem.genblk1[28].l_ram.data_out[7] ),
    .CLK(net2758));
 sg13g2_dfrbpq_1 _17873_ (.RESET_B(net926),
    .D(_01416_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[0] ),
    .CLK(net2759));
 sg13g2_dfrbpq_1 _17874_ (.RESET_B(net922),
    .D(_01417_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[1] ),
    .CLK(net2760));
 sg13g2_dfrbpq_1 _17875_ (.RESET_B(net913),
    .D(_01418_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[2] ),
    .CLK(net2761));
 sg13g2_dfrbpq_1 _17876_ (.RESET_B(net909),
    .D(_01419_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[3] ),
    .CLK(net2762));
 sg13g2_dfrbpq_1 _17877_ (.RESET_B(net905),
    .D(_01420_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[4] ),
    .CLK(net2763));
 sg13g2_dfrbpq_1 _17878_ (.RESET_B(net901),
    .D(_01421_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[5] ),
    .CLK(net2764));
 sg13g2_dfrbpq_1 _17879_ (.RESET_B(net897),
    .D(_01422_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[6] ),
    .CLK(net2765));
 sg13g2_dfrbpq_1 _17880_ (.RESET_B(net893),
    .D(_01423_),
    .Q(\i_latch_mem.genblk1[27].l_ram.data_out[7] ),
    .CLK(net2766));
 sg13g2_dfrbpq_1 _17881_ (.RESET_B(net889),
    .D(_01424_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[0] ),
    .CLK(net2767));
 sg13g2_dfrbpq_1 _17882_ (.RESET_B(net885),
    .D(_01425_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[1] ),
    .CLK(net2768));
 sg13g2_dfrbpq_1 _17883_ (.RESET_B(net881),
    .D(_01426_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[2] ),
    .CLK(net2769));
 sg13g2_dfrbpq_1 _17884_ (.RESET_B(net877),
    .D(_01427_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[3] ),
    .CLK(net2770));
 sg13g2_dfrbpq_1 _17885_ (.RESET_B(net872),
    .D(_01428_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[4] ),
    .CLK(net2771));
 sg13g2_dfrbpq_1 _17886_ (.RESET_B(net868),
    .D(_01429_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[5] ),
    .CLK(net2772));
 sg13g2_dfrbpq_1 _17887_ (.RESET_B(net864),
    .D(_01430_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[6] ),
    .CLK(net2773));
 sg13g2_dfrbpq_1 _17888_ (.RESET_B(net860),
    .D(_01431_),
    .Q(\i_latch_mem.genblk1[26].l_ram.data_out[7] ),
    .CLK(net2774));
 sg13g2_dfrbpq_1 _17889_ (.RESET_B(net856),
    .D(_01432_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[0] ),
    .CLK(net2775));
 sg13g2_dfrbpq_1 _17890_ (.RESET_B(net438),
    .D(_01433_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[1] ),
    .CLK(net2776));
 sg13g2_dfrbpq_1 _17891_ (.RESET_B(net406),
    .D(_01434_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[2] ),
    .CLK(net2777));
 sg13g2_dfrbpq_1 _17892_ (.RESET_B(net374),
    .D(_01435_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[3] ),
    .CLK(net2778));
 sg13g2_dfrbpq_1 _17893_ (.RESET_B(net370),
    .D(_01436_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[4] ),
    .CLK(net2779));
 sg13g2_dfrbpq_1 _17894_ (.RESET_B(net366),
    .D(_01437_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[5] ),
    .CLK(net2780));
 sg13g2_dfrbpq_1 _17895_ (.RESET_B(net362),
    .D(_01438_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[6] ),
    .CLK(net2781));
 sg13g2_dfrbpq_1 _17896_ (.RESET_B(net358),
    .D(_01439_),
    .Q(\i_latch_mem.genblk1[25].l_ram.data_out[7] ),
    .CLK(net2782));
 sg13g2_dfrbpq_1 _17897_ (.RESET_B(net354),
    .D(_01440_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[0] ),
    .CLK(net2783));
 sg13g2_dfrbpq_1 _17898_ (.RESET_B(net350),
    .D(_01441_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[1] ),
    .CLK(net2784));
 sg13g2_dfrbpq_1 _17899_ (.RESET_B(net346),
    .D(_01442_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[2] ),
    .CLK(net2785));
 sg13g2_dfrbpq_1 _17900_ (.RESET_B(net342),
    .D(_01443_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[3] ),
    .CLK(net2786));
 sg13g2_dfrbpq_1 _17901_ (.RESET_B(net338),
    .D(_01444_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[4] ),
    .CLK(net2787));
 sg13g2_dfrbpq_1 _17902_ (.RESET_B(net334),
    .D(_01445_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[5] ),
    .CLK(net2788));
 sg13g2_dfrbpq_1 _17903_ (.RESET_B(net330),
    .D(_01446_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[6] ),
    .CLK(net2789));
 sg13g2_dfrbpq_1 _17904_ (.RESET_B(net326),
    .D(_01447_),
    .Q(\i_latch_mem.genblk1[24].l_ram.data_out[7] ),
    .CLK(net2790));
 sg13g2_dfrbpq_1 _17905_ (.RESET_B(net322),
    .D(_01448_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[0] ),
    .CLK(net2791));
 sg13g2_dfrbpq_1 _17906_ (.RESET_B(net318),
    .D(_01449_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[1] ),
    .CLK(net2792));
 sg13g2_dfrbpq_1 _17907_ (.RESET_B(net314),
    .D(_01450_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[2] ),
    .CLK(net2793));
 sg13g2_dfrbpq_1 _17908_ (.RESET_B(net310),
    .D(_01451_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[3] ),
    .CLK(net2794));
 sg13g2_dfrbpq_1 _17909_ (.RESET_B(net305),
    .D(_01452_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[4] ),
    .CLK(net2795));
 sg13g2_dfrbpq_1 _17910_ (.RESET_B(net301),
    .D(_01453_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[5] ),
    .CLK(net2796));
 sg13g2_dfrbpq_1 _17911_ (.RESET_B(net296),
    .D(_01454_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[6] ),
    .CLK(net2797));
 sg13g2_dfrbpq_1 _17912_ (.RESET_B(net292),
    .D(_01455_),
    .Q(\i_latch_mem.genblk1[23].l_ram.data_out[7] ),
    .CLK(net2798));
 sg13g2_dfrbpq_1 _17913_ (.RESET_B(net288),
    .D(_01456_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[0] ),
    .CLK(net2799));
 sg13g2_dfrbpq_1 _17914_ (.RESET_B(net284),
    .D(_01457_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[1] ),
    .CLK(net2800));
 sg13g2_dfrbpq_1 _17915_ (.RESET_B(net280),
    .D(_01458_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[2] ),
    .CLK(net2801));
 sg13g2_dfrbpq_1 _17916_ (.RESET_B(net276),
    .D(_01459_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[3] ),
    .CLK(net2802));
 sg13g2_dfrbpq_1 _17917_ (.RESET_B(net272),
    .D(_01460_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[4] ),
    .CLK(net2803));
 sg13g2_dfrbpq_1 _17918_ (.RESET_B(net196),
    .D(_01461_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[5] ),
    .CLK(net2804));
 sg13g2_dfrbpq_1 _17919_ (.RESET_B(net188),
    .D(_01462_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[6] ),
    .CLK(net2805));
 sg13g2_dfrbpq_1 _17920_ (.RESET_B(net75),
    .D(_01463_),
    .Q(\i_latch_mem.genblk1[22].l_ram.data_out[7] ),
    .CLK(net2806));
 sg13g2_dfrbpq_1 _17921_ (.RESET_B(net2697),
    .D(_01464_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[0] ),
    .CLK(net2807));
 sg13g2_dfrbpq_1 _17922_ (.RESET_B(net1762),
    .D(_01465_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[1] ),
    .CLK(net2808));
 sg13g2_dfrbpq_1 _17923_ (.RESET_B(net1707),
    .D(_01466_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[2] ),
    .CLK(net2809));
 sg13g2_dfrbpq_1 _17924_ (.RESET_B(net1699),
    .D(_01467_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[3] ),
    .CLK(net2810));
 sg13g2_dfrbpq_1 _17925_ (.RESET_B(net1691),
    .D(_01468_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[4] ),
    .CLK(net2811));
 sg13g2_dfrbpq_1 _17926_ (.RESET_B(net1683),
    .D(_01469_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[5] ),
    .CLK(net2812));
 sg13g2_dfrbpq_2 _17927_ (.RESET_B(net1675),
    .D(_01470_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[6] ),
    .CLK(net2813));
 sg13g2_dfrbpq_1 _17928_ (.RESET_B(net1667),
    .D(_01471_),
    .Q(\i_latch_mem.genblk1[21].l_ram.data_out[7] ),
    .CLK(net2814));
 sg13g2_dfrbpq_1 _17929_ (.RESET_B(net1659),
    .D(_01472_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[0] ),
    .CLK(net2815));
 sg13g2_dfrbpq_1 _17930_ (.RESET_B(net1651),
    .D(_01473_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[1] ),
    .CLK(net2816));
 sg13g2_dfrbpq_1 _17931_ (.RESET_B(net1643),
    .D(_01474_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[2] ),
    .CLK(net2817));
 sg13g2_dfrbpq_1 _17932_ (.RESET_B(net1635),
    .D(_01475_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[3] ),
    .CLK(net2818));
 sg13g2_dfrbpq_1 _17933_ (.RESET_B(net1579),
    .D(_01476_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[4] ),
    .CLK(net2819));
 sg13g2_dfrbpq_1 _17934_ (.RESET_B(net1571),
    .D(_01477_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[5] ),
    .CLK(net2820));
 sg13g2_dfrbpq_1 _17935_ (.RESET_B(net1560),
    .D(_01478_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[6] ),
    .CLK(net2821));
 sg13g2_dfrbpq_1 _17936_ (.RESET_B(net1551),
    .D(_01479_),
    .Q(\i_latch_mem.genblk1[20].l_ram.data_out[7] ),
    .CLK(net2822));
 sg13g2_dfrbpq_1 _17937_ (.RESET_B(net1543),
    .D(_01480_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[0] ),
    .CLK(net2823));
 sg13g2_dfrbpq_1 _17938_ (.RESET_B(net1535),
    .D(_01481_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[1] ),
    .CLK(net2824));
 sg13g2_dfrbpq_1 _17939_ (.RESET_B(net1480),
    .D(_01482_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[2] ),
    .CLK(net2825));
 sg13g2_dfrbpq_1 _17940_ (.RESET_B(net1460),
    .D(_01483_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[3] ),
    .CLK(net2826));
 sg13g2_dfrbpq_1 _17941_ (.RESET_B(net1452),
    .D(_01484_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[4] ),
    .CLK(net2827));
 sg13g2_dfrbpq_1 _17942_ (.RESET_B(net1443),
    .D(_01485_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[5] ),
    .CLK(net2828));
 sg13g2_dfrbpq_1 _17943_ (.RESET_B(net1435),
    .D(_01486_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[6] ),
    .CLK(net2829));
 sg13g2_dfrbpq_1 _17944_ (.RESET_B(net1424),
    .D(_01487_),
    .Q(\i_latch_mem.genblk1[1].l_ram.data_out[7] ),
    .CLK(net2830));
 sg13g2_dfrbpq_1 _17945_ (.RESET_B(net1416),
    .D(_01488_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[0] ),
    .CLK(net2831));
 sg13g2_dfrbpq_1 _17946_ (.RESET_B(net1384),
    .D(_01489_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[1] ),
    .CLK(net2832));
 sg13g2_dfrbpq_1 _17947_ (.RESET_B(net1376),
    .D(_01490_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[2] ),
    .CLK(net2833));
 sg13g2_dfrbpq_1 _17948_ (.RESET_B(net1367),
    .D(_01491_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[3] ),
    .CLK(net2834));
 sg13g2_dfrbpq_1 _17949_ (.RESET_B(net1359),
    .D(_01492_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[4] ),
    .CLK(net2835));
 sg13g2_dfrbpq_1 _17950_ (.RESET_B(net1351),
    .D(_01493_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[5] ),
    .CLK(net2836));
 sg13g2_dfrbpq_1 _17951_ (.RESET_B(net1343),
    .D(_01494_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[6] ),
    .CLK(net2837));
 sg13g2_dfrbpq_1 _17952_ (.RESET_B(net1334),
    .D(_01495_),
    .Q(\i_latch_mem.genblk1[18].l_ram.data_out[7] ),
    .CLK(net2838));
 sg13g2_dfrbpq_1 _17953_ (.RESET_B(net1326),
    .D(_01496_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[0] ),
    .CLK(net2839));
 sg13g2_dfrbpq_1 _17954_ (.RESET_B(net1318),
    .D(_01497_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[1] ),
    .CLK(net2840));
 sg13g2_dfrbpq_1 _17955_ (.RESET_B(net1310),
    .D(_01498_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[2] ),
    .CLK(net2841));
 sg13g2_dfrbpq_1 _17956_ (.RESET_B(net1301),
    .D(_01499_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[3] ),
    .CLK(net2842));
 sg13g2_dfrbpq_1 _17957_ (.RESET_B(net1293),
    .D(_01500_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[4] ),
    .CLK(net2843));
 sg13g2_dfrbpq_1 _17958_ (.RESET_B(net1285),
    .D(_01501_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[5] ),
    .CLK(net2844));
 sg13g2_dfrbpq_1 _17959_ (.RESET_B(net1277),
    .D(_01502_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[6] ),
    .CLK(net2845));
 sg13g2_dfrbpq_1 _17960_ (.RESET_B(net1269),
    .D(_01503_),
    .Q(\i_latch_mem.genblk1[17].l_ram.data_out[7] ),
    .CLK(net2846));
 sg13g2_dfrbpq_1 _17961_ (.RESET_B(net1261),
    .D(_01504_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[0] ),
    .CLK(net2847));
 sg13g2_dfrbpq_1 _17962_ (.RESET_B(net1253),
    .D(_01505_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[1] ),
    .CLK(net2848));
 sg13g2_dfrbpq_1 _17963_ (.RESET_B(net1245),
    .D(_01506_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[2] ),
    .CLK(net2849));
 sg13g2_dfrbpq_1 _17964_ (.RESET_B(net1225),
    .D(_01507_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[3] ),
    .CLK(net2850));
 sg13g2_dfrbpq_1 _17965_ (.RESET_B(net1217),
    .D(_01508_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[4] ),
    .CLK(net2851));
 sg13g2_dfrbpq_1 _17966_ (.RESET_B(net1209),
    .D(_01509_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[5] ),
    .CLK(net2852));
 sg13g2_dfrbpq_1 _17967_ (.RESET_B(net1201),
    .D(_01510_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[6] ),
    .CLK(net2853));
 sg13g2_dfrbpq_1 _17968_ (.RESET_B(net1193),
    .D(_01511_),
    .Q(\i_latch_mem.genblk1[16].l_ram.data_out[7] ),
    .CLK(net2854));
 sg13g2_dfrbpq_1 _17969_ (.RESET_B(net1184),
    .D(_01512_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[0] ),
    .CLK(net2855));
 sg13g2_dfrbpq_1 _17970_ (.RESET_B(net1176),
    .D(_01513_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[1] ),
    .CLK(net2856));
 sg13g2_dfrbpq_1 _17971_ (.RESET_B(net1168),
    .D(_01514_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[2] ),
    .CLK(net2857));
 sg13g2_dfrbpq_1 _17972_ (.RESET_B(net1160),
    .D(_01515_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[3] ),
    .CLK(net2858));
 sg13g2_dfrbpq_1 _17973_ (.RESET_B(net1152),
    .D(_01516_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[4] ),
    .CLK(net2859));
 sg13g2_dfrbpq_1 _17974_ (.RESET_B(net1144),
    .D(_01517_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[5] ),
    .CLK(net2860));
 sg13g2_dfrbpq_1 _17975_ (.RESET_B(net1102),
    .D(_01518_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[6] ),
    .CLK(net2861));
 sg13g2_dfrbpq_1 _17976_ (.RESET_B(net1090),
    .D(_01519_),
    .Q(\i_latch_mem.genblk1[15].l_ram.data_out[7] ),
    .CLK(net2862));
 sg13g2_dfrbpq_1 _17977_ (.RESET_B(net1082),
    .D(_01520_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[0] ),
    .CLK(net2863));
 sg13g2_dfrbpq_1 _17978_ (.RESET_B(net1072),
    .D(_01521_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[1] ),
    .CLK(net2864));
 sg13g2_dfrbpq_1 _17979_ (.RESET_B(net1062),
    .D(_01522_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[2] ),
    .CLK(net2865));
 sg13g2_dfrbpq_1 _17980_ (.RESET_B(net1054),
    .D(_01523_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[3] ),
    .CLK(net2866));
 sg13g2_dfrbpq_1 _17981_ (.RESET_B(net1044),
    .D(_01524_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[4] ),
    .CLK(net2867));
 sg13g2_dfrbpq_1 _17982_ (.RESET_B(net1036),
    .D(_01525_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[5] ),
    .CLK(net2868));
 sg13g2_dfrbpq_2 _17983_ (.RESET_B(net1024),
    .D(_01526_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[6] ),
    .CLK(net2869));
 sg13g2_dfrbpq_2 _17984_ (.RESET_B(net1016),
    .D(_01527_),
    .Q(\i_latch_mem.genblk1[14].l_ram.data_out[7] ),
    .CLK(net2870));
 sg13g2_dfrbpq_1 _17985_ (.RESET_B(net1008),
    .D(_01528_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[0] ),
    .CLK(net2871));
 sg13g2_dfrbpq_1 _17986_ (.RESET_B(net1000),
    .D(_01529_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[1] ),
    .CLK(net2872));
 sg13g2_dfrbpq_1 _17987_ (.RESET_B(net992),
    .D(_01530_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[2] ),
    .CLK(net2873));
 sg13g2_dfrbpq_1 _17988_ (.RESET_B(net984),
    .D(_01531_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[3] ),
    .CLK(net2874));
 sg13g2_dfrbpq_1 _17989_ (.RESET_B(net976),
    .D(_01532_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[4] ),
    .CLK(net2875));
 sg13g2_dfrbpq_1 _17990_ (.RESET_B(net968),
    .D(_01533_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[5] ),
    .CLK(net2876));
 sg13g2_dfrbpq_1 _17991_ (.RESET_B(net960),
    .D(_01534_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[6] ),
    .CLK(net2877));
 sg13g2_dfrbpq_1 _17992_ (.RESET_B(net952),
    .D(_01535_),
    .Q(\i_latch_mem.genblk1[13].l_ram.data_out[7] ),
    .CLK(net2878));
 sg13g2_dfrbpq_1 _17993_ (.RESET_B(net944),
    .D(_01536_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[0] ),
    .CLK(net2879));
 sg13g2_dfrbpq_1 _17994_ (.RESET_B(net936),
    .D(_01537_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[1] ),
    .CLK(net2880));
 sg13g2_dfrbpq_1 _17995_ (.RESET_B(net928),
    .D(_01538_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[2] ),
    .CLK(net2881));
 sg13g2_dfrbpq_1 _17996_ (.RESET_B(net920),
    .D(_01539_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[3] ),
    .CLK(net2882));
 sg13g2_dfrbpq_1 _17997_ (.RESET_B(net907),
    .D(_01540_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[4] ),
    .CLK(net2883));
 sg13g2_dfrbpq_1 _17998_ (.RESET_B(net899),
    .D(_01541_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[5] ),
    .CLK(net2884));
 sg13g2_dfrbpq_1 _17999_ (.RESET_B(net891),
    .D(_01542_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[6] ),
    .CLK(net2885));
 sg13g2_dfrbpq_1 _18000_ (.RESET_B(net883),
    .D(_01543_),
    .Q(\i_latch_mem.genblk1[12].l_ram.data_out[7] ),
    .CLK(net2886));
 sg13g2_dfrbpq_1 _18001_ (.RESET_B(net874),
    .D(_01544_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[0] ),
    .CLK(net2887));
 sg13g2_dfrbpq_1 _18002_ (.RESET_B(net866),
    .D(_01545_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[1] ),
    .CLK(net2888));
 sg13g2_dfrbpq_1 _18003_ (.RESET_B(net858),
    .D(_01546_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[2] ),
    .CLK(net2889));
 sg13g2_dfrbpq_1 _18004_ (.RESET_B(net436),
    .D(_01547_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[3] ),
    .CLK(net2890));
 sg13g2_dfrbpq_1 _18005_ (.RESET_B(net372),
    .D(_01548_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[4] ),
    .CLK(net2891));
 sg13g2_dfrbpq_1 _18006_ (.RESET_B(net364),
    .D(_01549_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[5] ),
    .CLK(net2892));
 sg13g2_dfrbpq_1 _18007_ (.RESET_B(net356),
    .D(_01550_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[6] ),
    .CLK(net2893));
 sg13g2_dfrbpq_1 _18008_ (.RESET_B(net348),
    .D(_01551_),
    .Q(\i_latch_mem.genblk1[11].l_ram.data_out[7] ),
    .CLK(net2894));
 sg13g2_dfrbpq_1 _18009_ (.RESET_B(net340),
    .D(_01552_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[0] ),
    .CLK(net2895));
 sg13g2_dfrbpq_1 _18010_ (.RESET_B(net332),
    .D(_01553_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[1] ),
    .CLK(net2896));
 sg13g2_dfrbpq_1 _18011_ (.RESET_B(net324),
    .D(_01554_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[2] ),
    .CLK(net2897));
 sg13g2_dfrbpq_2 _18012_ (.RESET_B(net316),
    .D(_01555_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[3] ),
    .CLK(net2898));
 sg13g2_dfrbpq_1 _18013_ (.RESET_B(net307),
    .D(_01556_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[4] ),
    .CLK(net2899));
 sg13g2_dfrbpq_1 _18014_ (.RESET_B(net299),
    .D(_01557_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[5] ),
    .CLK(net2900));
 sg13g2_dfrbpq_1 _18015_ (.RESET_B(net290),
    .D(_01558_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[6] ),
    .CLK(net2901));
 sg13g2_dfrbpq_1 _18016_ (.RESET_B(net282),
    .D(_01559_),
    .Q(\i_latch_mem.genblk1[10].l_ram.data_out[7] ),
    .CLK(net2902));
 sg13g2_dfrbpq_1 _18017_ (.RESET_B(net274),
    .D(_01560_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[0] ),
    .CLK(net2903));
 sg13g2_dfrbpq_1 _18018_ (.RESET_B(net192),
    .D(_01561_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[1] ),
    .CLK(net2904));
 sg13g2_dfrbpq_1 _18019_ (.RESET_B(net71),
    .D(_01562_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[2] ),
    .CLK(net2905));
 sg13g2_dfrbpq_1 _18020_ (.RESET_B(net1742),
    .D(_01563_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[3] ),
    .CLK(net2906));
 sg13g2_dfrbpq_1 _18021_ (.RESET_B(net1695),
    .D(_01564_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[4] ),
    .CLK(net2907));
 sg13g2_dfrbpq_1 _18022_ (.RESET_B(net1679),
    .D(_01565_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[5] ),
    .CLK(net2908));
 sg13g2_dfrbpq_1 _18023_ (.RESET_B(net1663),
    .D(_01566_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[6] ),
    .CLK(net2909));
 sg13g2_dfrbpq_1 _18024_ (.RESET_B(net1647),
    .D(_01567_),
    .Q(\i_latch_mem.genblk1[0].l_ram.data_out[7] ),
    .CLK(net2910));
 sg13g2_dfrbpq_1 _18025_ (.RESET_B(net1611),
    .D(_01568_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[0] ),
    .CLK(net2911));
 sg13g2_dfrbpq_1 _18026_ (.RESET_B(net1567),
    .D(_01569_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[1] ),
    .CLK(net2912));
 sg13g2_dfrbpq_1 _18027_ (.RESET_B(net1547),
    .D(_01570_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[2] ),
    .CLK(net2913));
 sg13g2_dfrbpq_1 _18028_ (.RESET_B(net1484),
    .D(_01571_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[3] ),
    .CLK(net2914));
 sg13g2_dfrbpq_1 _18029_ (.RESET_B(net1456),
    .D(_01572_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[4] ),
    .CLK(net2915));
 sg13g2_dfrbpq_1 _18030_ (.RESET_B(net1439),
    .D(_01573_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[5] ),
    .CLK(net2916));
 sg13g2_dfrbpq_1 _18031_ (.RESET_B(net1420),
    .D(_01574_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[6] ),
    .CLK(net2917));
 sg13g2_dfrbpq_1 _18032_ (.RESET_B(net1380),
    .D(_01575_),
    .Q(\i_latch_mem.genblk1[8].l_ram.data_out[7] ),
    .CLK(net2918));
 sg13g2_dfrbpq_1 _18033_ (.RESET_B(net1363),
    .D(_01576_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[0] ),
    .CLK(net2919));
 sg13g2_dfrbpq_1 _18034_ (.RESET_B(net1347),
    .D(_01577_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[1] ),
    .CLK(net2920));
 sg13g2_dfrbpq_1 _18035_ (.RESET_B(net1330),
    .D(_01578_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[2] ),
    .CLK(net2921));
 sg13g2_dfrbpq_1 _18036_ (.RESET_B(net1314),
    .D(_01579_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[3] ),
    .CLK(net2922));
 sg13g2_dfrbpq_1 _18037_ (.RESET_B(net1297),
    .D(_01580_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[4] ),
    .CLK(net2923));
 sg13g2_dfrbpq_1 _18038_ (.RESET_B(net1281),
    .D(_01581_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[5] ),
    .CLK(net2924));
 sg13g2_dfrbpq_1 _18039_ (.RESET_B(net1265),
    .D(_01582_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[6] ),
    .CLK(net2925));
 sg13g2_dfrbpq_1 _18040_ (.RESET_B(net1249),
    .D(_01583_),
    .Q(\i_latch_mem.genblk1[7].l_ram.data_out[7] ),
    .CLK(net2926));
 sg13g2_dfrbpq_1 _18041_ (.RESET_B(net1221),
    .D(_01584_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[0] ),
    .CLK(net2927));
 sg13g2_dfrbpq_1 _18042_ (.RESET_B(net1205),
    .D(_01585_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[1] ),
    .CLK(net2928));
 sg13g2_dfrbpq_1 _18043_ (.RESET_B(net1189),
    .D(_01586_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[2] ),
    .CLK(net2929));
 sg13g2_dfrbpq_2 _18044_ (.RESET_B(net1172),
    .D(_01587_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[3] ),
    .CLK(net2930));
 sg13g2_dfrbpq_1 _18045_ (.RESET_B(net1156),
    .D(_01588_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[4] ),
    .CLK(net2931));
 sg13g2_dfrbpq_1 _18046_ (.RESET_B(net1140),
    .D(_01589_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[5] ),
    .CLK(net2932));
 sg13g2_dfrbpq_1 _18047_ (.RESET_B(net1086),
    .D(_01590_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[6] ),
    .CLK(net2933));
 sg13g2_dfrbpq_2 _18048_ (.RESET_B(net1066),
    .D(_01591_),
    .Q(\i_latch_mem.genblk1[6].l_ram.data_out[7] ),
    .CLK(net2934));
 sg13g2_dfrbpq_1 _18049_ (.RESET_B(net1048),
    .D(_01592_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[0] ),
    .CLK(net2935));
 sg13g2_dfrbpq_1 _18050_ (.RESET_B(net1030),
    .D(_01593_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[1] ),
    .CLK(net2936));
 sg13g2_dfrbpq_1 _18051_ (.RESET_B(net1012),
    .D(_01594_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[2] ),
    .CLK(net2937));
 sg13g2_dfrbpq_1 _18052_ (.RESET_B(net996),
    .D(_01595_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[3] ),
    .CLK(net2938));
 sg13g2_dfrbpq_1 _18053_ (.RESET_B(net980),
    .D(_01596_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[4] ),
    .CLK(net2939));
 sg13g2_dfrbpq_1 _18054_ (.RESET_B(net964),
    .D(_01597_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[5] ),
    .CLK(net2940));
 sg13g2_dfrbpq_2 _18055_ (.RESET_B(net948),
    .D(_01598_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[6] ),
    .CLK(net2941));
 sg13g2_dfrbpq_2 _18056_ (.RESET_B(net932),
    .D(_01599_),
    .Q(\i_latch_mem.genblk1[5].l_ram.data_out[7] ),
    .CLK(net2942));
 sg13g2_dfrbpq_1 _18057_ (.RESET_B(net911),
    .D(_01600_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[0] ),
    .CLK(net2943));
 sg13g2_dfrbpq_1 _18058_ (.RESET_B(net895),
    .D(_01601_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[1] ),
    .CLK(net2944));
 sg13g2_dfrbpq_1 _18059_ (.RESET_B(net879),
    .D(_01602_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[2] ),
    .CLK(net2945));
 sg13g2_dfrbpq_1 _18060_ (.RESET_B(net862),
    .D(_01603_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[3] ),
    .CLK(net2946));
 sg13g2_dfrbpq_1 _18061_ (.RESET_B(net404),
    .D(_01604_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[4] ),
    .CLK(net2947));
 sg13g2_dfrbpq_1 _18062_ (.RESET_B(net360),
    .D(_01605_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[5] ),
    .CLK(net2948));
 sg13g2_dfrbpq_1 _18063_ (.RESET_B(net344),
    .D(_01606_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[6] ),
    .CLK(net2949));
 sg13g2_dfrbpq_1 _18064_ (.RESET_B(net328),
    .D(_01607_),
    .Q(\i_latch_mem.genblk1[4].l_ram.data_out[7] ),
    .CLK(net2950));
 sg13g2_dfrbpq_1 _18065_ (.RESET_B(net312),
    .D(_01608_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[0] ),
    .CLK(net2951));
 sg13g2_dfrbpq_1 _18066_ (.RESET_B(net294),
    .D(_01609_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[1] ),
    .CLK(net2952));
 sg13g2_dfrbpq_1 _18067_ (.RESET_B(net278),
    .D(_01610_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[2] ),
    .CLK(net2953));
 sg13g2_dfrbpq_1 _18068_ (.RESET_B(net115),
    .D(_01611_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[3] ),
    .CLK(net2954));
 sg13g2_dfrbpq_1 _18069_ (.RESET_B(net1703),
    .D(_01612_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[4] ),
    .CLK(net2955));
 sg13g2_dfrbpq_1 _18070_ (.RESET_B(net1671),
    .D(_01613_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[5] ),
    .CLK(net2956));
 sg13g2_dfrbpq_1 _18071_ (.RESET_B(net1639),
    .D(_01614_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[6] ),
    .CLK(net2957));
 sg13g2_dfrbpq_2 _18072_ (.RESET_B(net1555),
    .D(_01615_),
    .Q(\i_latch_mem.genblk1[3].l_ram.data_out[7] ),
    .CLK(net2958));
 sg13g2_dfrbpq_1 _18073_ (.RESET_B(net1476),
    .D(_01616_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[0] ),
    .CLK(net2959));
 sg13g2_dfrbpq_1 _18074_ (.RESET_B(net1430),
    .D(_01617_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[1] ),
    .CLK(net2960));
 sg13g2_dfrbpq_1 _18075_ (.RESET_B(net1371),
    .D(_01618_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[2] ),
    .CLK(net2961));
 sg13g2_dfrbpq_1 _18076_ (.RESET_B(net1339),
    .D(_01619_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[3] ),
    .CLK(net2962));
 sg13g2_dfrbpq_1 _18077_ (.RESET_B(net1306),
    .D(_01620_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[4] ),
    .CLK(net2963));
 sg13g2_dfrbpq_1 _18078_ (.RESET_B(net1273),
    .D(_01621_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[5] ),
    .CLK(net2964));
 sg13g2_dfrbpq_1 _18079_ (.RESET_B(net1241),
    .D(_01622_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[6] ),
    .CLK(net2965));
 sg13g2_dfrbpq_1 _18080_ (.RESET_B(net1197),
    .D(_01623_),
    .Q(\i_latch_mem.genblk1[31].l_ram.data_out[7] ),
    .CLK(net2966));
 sg13g2_dfrbpq_1 _18081_ (.RESET_B(net1164),
    .D(_01624_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[0] ),
    .CLK(net2967));
 sg13g2_dfrbpq_1 _18082_ (.RESET_B(net1094),
    .D(_01625_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[1] ),
    .CLK(net2968));
 sg13g2_dfrbpq_1 _18083_ (.RESET_B(net1058),
    .D(_01626_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[2] ),
    .CLK(net2969));
 sg13g2_dfrbpq_2 _18084_ (.RESET_B(net1020),
    .D(_01627_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[3] ),
    .CLK(net2970));
 sg13g2_dfrbpq_1 _18085_ (.RESET_B(net988),
    .D(_01628_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[4] ),
    .CLK(net2971));
 sg13g2_dfrbpq_1 _18086_ (.RESET_B(net956),
    .D(_01629_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[5] ),
    .CLK(net2972));
 sg13g2_dfrbpq_2 _18087_ (.RESET_B(net924),
    .D(_01630_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[6] ),
    .CLK(net2973));
 sg13g2_dfrbpq_2 _18088_ (.RESET_B(net887),
    .D(_01631_),
    .Q(\i_latch_mem.genblk1[29].l_ram.data_out[7] ),
    .CLK(net2974));
 sg13g2_dfrbpq_1 _18089_ (.RESET_B(net440),
    .D(_01632_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[0] ),
    .CLK(net2975));
 sg13g2_dfrbpq_1 _18090_ (.RESET_B(net352),
    .D(_01633_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[1] ),
    .CLK(net2976));
 sg13g2_dfrbpq_1 _18091_ (.RESET_B(net320),
    .D(_01634_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[2] ),
    .CLK(net2977));
 sg13g2_dfrbpq_1 _18092_ (.RESET_B(net286),
    .D(_01635_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[3] ),
    .CLK(net2978));
 sg13g2_dfrbpq_1 _18093_ (.RESET_B(net2690),
    .D(_01636_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[4] ),
    .CLK(net2979));
 sg13g2_dfrbpq_1 _18094_ (.RESET_B(net1655),
    .D(_01637_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[5] ),
    .CLK(net2980));
 sg13g2_dfrbpq_1 _18095_ (.RESET_B(net1539),
    .D(_01638_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[6] ),
    .CLK(net2981));
 sg13g2_dfrbpq_1 _18096_ (.RESET_B(net1412),
    .D(_01639_),
    .Q(\i_latch_mem.genblk1[19].l_ram.data_out[7] ),
    .CLK(net2982));
 sg13g2_dfrbpq_1 _18097_ (.RESET_B(net1775),
    .D(_01640_),
    .Q(\i_latch_mem.data_ready ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _18098_ (.RESET_B(net1776),
    .D(_00012_),
    .Q(\i_latch_mem.data_out[0] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _18099_ (.RESET_B(net1777),
    .D(_00023_),
    .Q(\i_latch_mem.data_out[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _18100_ (.RESET_B(net1778),
    .D(_00034_),
    .Q(\i_latch_mem.data_out[2] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _18101_ (.RESET_B(net1779),
    .D(_00037_),
    .Q(\i_latch_mem.data_out[3] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _18102_ (.RESET_B(net1780),
    .D(_00038_),
    .Q(\i_latch_mem.data_out[4] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _18103_ (.RESET_B(net1781),
    .D(_00039_),
    .Q(\i_latch_mem.data_out[5] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18104_ (.RESET_B(net1782),
    .D(_00040_),
    .Q(\i_latch_mem.data_out[6] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _18105_ (.RESET_B(net1783),
    .D(_00041_),
    .Q(\i_latch_mem.data_out[7] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _18106_ (.RESET_B(net1784),
    .D(_00042_),
    .Q(\i_latch_mem.data_out[8] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _18107_ (.RESET_B(net1785),
    .D(_00043_),
    .Q(\i_latch_mem.data_out[9] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _18108_ (.RESET_B(net1786),
    .D(net3854),
    .Q(\i_latch_mem.data_out[10] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _18109_ (.RESET_B(net1787),
    .D(_00014_),
    .Q(\i_latch_mem.data_out[11] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _18110_ (.RESET_B(net1788),
    .D(_00015_),
    .Q(\i_latch_mem.data_out[12] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _18111_ (.RESET_B(net1789),
    .D(_00016_),
    .Q(\i_latch_mem.data_out[13] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18112_ (.RESET_B(net1790),
    .D(_00017_),
    .Q(\i_latch_mem.data_out[14] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _18113_ (.RESET_B(net1791),
    .D(_00018_),
    .Q(\i_latch_mem.data_out[15] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _18114_ (.RESET_B(net1792),
    .D(net3915),
    .Q(\i_latch_mem.data_out[16] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _18115_ (.RESET_B(net2675),
    .D(_00020_),
    .Q(\i_latch_mem.data_out[17] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18116_ (.RESET_B(net2676),
    .D(_00021_),
    .Q(\i_latch_mem.data_out[18] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18117_ (.RESET_B(net2677),
    .D(_00022_),
    .Q(\i_latch_mem.data_out[19] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _18118_ (.RESET_B(net2678),
    .D(_00024_),
    .Q(\i_latch_mem.data_out[20] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _18119_ (.RESET_B(net2679),
    .D(_00025_),
    .Q(\i_latch_mem.data_out[21] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18120_ (.RESET_B(net2680),
    .D(_00026_),
    .Q(\i_latch_mem.data_out[22] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18121_ (.RESET_B(net2681),
    .D(_00027_),
    .Q(\i_latch_mem.data_out[23] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18122_ (.RESET_B(net2682),
    .D(net3491),
    .Q(\i_latch_mem.data_out[24] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _18123_ (.RESET_B(net2683),
    .D(_00029_),
    .Q(\i_latch_mem.data_out[25] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _18124_ (.RESET_B(net2684),
    .D(_00030_),
    .Q(\i_latch_mem.data_out[26] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _18125_ (.RESET_B(net2685),
    .D(_00031_),
    .Q(\i_latch_mem.data_out[27] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _18126_ (.RESET_B(net2686),
    .D(net3642),
    .Q(\i_latch_mem.data_out[28] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _18127_ (.RESET_B(net2687),
    .D(net3624),
    .Q(\i_latch_mem.data_out[29] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _18128_ (.RESET_B(net1448),
    .D(net3663),
    .Q(\i_latch_mem.data_out[30] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _18129_ (.RESET_B(net1322),
    .D(_00036_),
    .Q(\i_latch_mem.data_out[31] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_2 _18130_ (.RESET_B(net1289),
    .D(_01641_),
    .Q(\i_i2c_peri.i_i2c.missed_ack_reg ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _18131_ (.RESET_B(net1257),
    .D(net5026),
    .Q(\i_latch_mem.cycle[1] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _18132_ (.RESET_B(net1180),
    .D(net3610),
    .Q(\i_i2c_peri.i_i2c.data_reg[7] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _18133_ (.RESET_B(net1076),
    .D(net4442),
    .Q(\i_i2c_peri.i_i2c.data_reg[6] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _18134_ (.RESET_B(net1004),
    .D(net4478),
    .Q(\i_i2c_peri.i_i2c.data_reg[5] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _18135_ (.RESET_B(net940),
    .D(net4368),
    .Q(\i_i2c_peri.i_i2c.data_reg[4] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _18136_ (.RESET_B(net870),
    .D(net4375),
    .Q(\i_i2c_peri.i_i2c.data_reg[3] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _18137_ (.RESET_B(net336),
    .D(net4536),
    .Q(\i_i2c_peri.i_i2c.data_reg[2] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _18138_ (.RESET_B(net200),
    .D(net4641),
    .Q(\i_i2c_peri.i_i2c.data_reg[1] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _18139_ (.RESET_B(net1575),
    .D(_01650_),
    .Q(\i_i2c_peri.i_i2c.data_reg[0] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _18140_ (.RESET_B(net1355),
    .D(_01651_),
    .Q(\i_i2c_peri.i_i2c.s_axis_cmd_ready_reg ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _18141_ (.RESET_B(net1213),
    .D(_01652_),
    .Q(\i_i2c_peri.i_i2c.s_axis_data_tready_reg ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _18142_ (.RESET_B(net1148),
    .D(net3578),
    .Q(\i_tinyqv.cpu.i_core.mie[4] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _18143_ (.RESET_B(net972),
    .D(net3557),
    .Q(\i_tinyqv.cpu.i_core.mie[3] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_2 _18144_ (.RESET_B(net368),
    .D(net4178),
    .Q(\i_tinyqv.cpu.i_core.mie[2] ),
    .CLK(clknet_leaf_181_clk_regs));
 sg13g2_dfrbpq_2 _18145_ (.RESET_B(net1687),
    .D(net4123),
    .Q(\i_tinyqv.cpu.i_core.mie[1] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_2 _18146_ (.RESET_B(net1040),
    .D(_01657_),
    .Q(\i_tinyqv.cpu.i_core.mie[0] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_2 _18147_ (.RESET_B(net303),
    .D(_01658_),
    .Q(\i_tinyqv.cpu.i_core.mip[1] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_2 _18148_ (.RESET_B(net903),
    .D(net4358),
    .Q(\i_tinyqv.cpu.i_core.mip[0] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_tiehi _16472__15 (.L_HI(net15));
 sg13g2_tiehi _16471__16 (.L_HI(net16));
 sg13g2_tiehi _16470__17 (.L_HI(net17));
 sg13g2_tiehi _16469__18 (.L_HI(net18));
 sg13g2_tiehi _16468__19 (.L_HI(net19));
 sg13g2_tiehi _16467__20 (.L_HI(net20));
 sg13g2_tiehi _16466__21 (.L_HI(net21));
 sg13g2_tiehi _16465__22 (.L_HI(net22));
 sg13g2_tiehi _16464__23 (.L_HI(net23));
 sg13g2_tiehi _16463__24 (.L_HI(net24));
 sg13g2_tiehi _16462__25 (.L_HI(net25));
 sg13g2_tiehi _16461__26 (.L_HI(net26));
 sg13g2_tiehi _16460__27 (.L_HI(net27));
 sg13g2_tiehi _16459__28 (.L_HI(net28));
 sg13g2_tiehi _16458__29 (.L_HI(net29));
 sg13g2_tiehi _16457__30 (.L_HI(net30));
 sg13g2_tiehi _16456__31 (.L_HI(net31));
 sg13g2_tiehi _16455__32 (.L_HI(net32));
 sg13g2_tiehi _16454__33 (.L_HI(net33));
 sg13g2_tiehi _16453__34 (.L_HI(net34));
 sg13g2_tiehi _16452__35 (.L_HI(net35));
 sg13g2_tiehi _17666__36 (.L_HI(net36));
 sg13g2_tiehi _16451__37 (.L_HI(net37));
 sg13g2_tiehi _17665__38 (.L_HI(net38));
 sg13g2_tiehi _16450__39 (.L_HI(net39));
 sg13g2_tiehi _16449__40 (.L_HI(net40));
 sg13g2_tiehi _16448__41 (.L_HI(net41));
 sg13g2_tiehi _16447__42 (.L_HI(net42));
 sg13g2_tiehi _16446__43 (.L_HI(net43));
 sg13g2_tiehi _17664__44 (.L_HI(net44));
 sg13g2_tiehi _16445__45 (.L_HI(net45));
 sg13g2_tiehi _16443__46 (.L_HI(net46));
 sg13g2_tiehi _16442__47 (.L_HI(net47));
 sg13g2_tiehi _16441__48 (.L_HI(net48));
 sg13g2_tiehi _16440__49 (.L_HI(net49));
 sg13g2_tiehi _16439__50 (.L_HI(net50));
 sg13g2_tiehi _16438__51 (.L_HI(net51));
 sg13g2_tiehi _16437__52 (.L_HI(net52));
 sg13g2_tiehi _16436__53 (.L_HI(net53));
 sg13g2_tiehi _16435__54 (.L_HI(net54));
 sg13g2_tiehi _16434__55 (.L_HI(net55));
 sg13g2_tiehi _16433__56 (.L_HI(net56));
 sg13g2_tiehi _16432__57 (.L_HI(net57));
 sg13g2_tiehi _16431__58 (.L_HI(net58));
 sg13g2_tiehi _16430__59 (.L_HI(net59));
 sg13g2_tiehi _16429__60 (.L_HI(net60));
 sg13g2_tiehi _16428__61 (.L_HI(net61));
 sg13g2_tiehi _16427__62 (.L_HI(net62));
 sg13g2_tiehi _16426__63 (.L_HI(net63));
 sg13g2_tiehi _16425__64 (.L_HI(net64));
 sg13g2_tiehi _17663__65 (.L_HI(net65));
 sg13g2_tiehi _16424__66 (.L_HI(net66));
 sg13g2_tiehi _17662__67 (.L_HI(net67));
 sg13g2_tiehi _16423__68 (.L_HI(net68));
 sg13g2_tiehi _17661__69 (.L_HI(net69));
 sg13g2_tiehi _16422__70 (.L_HI(net70));
 sg13g2_tiehi _18019__71 (.L_HI(net71));
 sg13g2_tiehi _16421__72 (.L_HI(net72));
 sg13g2_tiehi _17660__73 (.L_HI(net73));
 sg13g2_tiehi _16420__74 (.L_HI(net74));
 sg13g2_tiehi _17920__75 (.L_HI(net75));
 sg13g2_tiehi _16419__76 (.L_HI(net76));
 sg13g2_tiehi _17658__77 (.L_HI(net77));
 sg13g2_tiehi _16418__78 (.L_HI(net78));
 sg13g2_tiehi _17657__79 (.L_HI(net79));
 sg13g2_tiehi _16417__80 (.L_HI(net80));
 sg13g2_tiehi _17656__81 (.L_HI(net81));
 sg13g2_tiehi _16416__82 (.L_HI(net82));
 sg13g2_tiehi _17655__83 (.L_HI(net83));
 sg13g2_tiehi _16415__84 (.L_HI(net84));
 sg13g2_tiehi _16414__85 (.L_HI(net85));
 sg13g2_tiehi _17654__86 (.L_HI(net86));
 sg13g2_tiehi _16412__87 (.L_HI(net87));
 sg13g2_tiehi _17653__88 (.L_HI(net88));
 sg13g2_tiehi _16411__89 (.L_HI(net89));
 sg13g2_tiehi _16324__90 (.L_HI(net90));
 sg13g2_tiehi _17652__91 (.L_HI(net91));
 sg13g2_tiehi _16410__92 (.L_HI(net92));
 sg13g2_tiehi _17651__93 (.L_HI(net93));
 sg13g2_tiehi _16409__94 (.L_HI(net94));
 sg13g2_tiehi _17650__95 (.L_HI(net95));
 sg13g2_tiehi _16408__96 (.L_HI(net96));
 sg13g2_tiehi _17649__97 (.L_HI(net97));
 sg13g2_tiehi _16407__98 (.L_HI(net98));
 sg13g2_tiehi _17648__99 (.L_HI(net99));
 sg13g2_tiehi _16406__100 (.L_HI(net100));
 sg13g2_tiehi _17647__101 (.L_HI(net101));
 sg13g2_tiehi _16405__102 (.L_HI(net102));
 sg13g2_tiehi _17646__103 (.L_HI(net103));
 sg13g2_tiehi _16404__104 (.L_HI(net104));
 sg13g2_tiehi _17645__105 (.L_HI(net105));
 sg13g2_tiehi _16403__106 (.L_HI(net106));
 sg13g2_tiehi _17644__107 (.L_HI(net107));
 sg13g2_tiehi _16402__108 (.L_HI(net108));
 sg13g2_tiehi _17643__109 (.L_HI(net109));
 sg13g2_tiehi _16401__110 (.L_HI(net110));
 sg13g2_tiehi _17642__111 (.L_HI(net111));
 sg13g2_tiehi _16400__112 (.L_HI(net112));
 sg13g2_tiehi _17641__113 (.L_HI(net113));
 sg13g2_tiehi _16399__114 (.L_HI(net114));
 sg13g2_tiehi _18068__115 (.L_HI(net115));
 sg13g2_tiehi _16398__116 (.L_HI(net116));
 sg13g2_tiehi _17640__117 (.L_HI(net117));
 sg13g2_tiehi _16397__118 (.L_HI(net118));
 sg13g2_tiehi _17639__119 (.L_HI(net119));
 sg13g2_tiehi _16396__120 (.L_HI(net120));
 sg13g2_tiehi _16413__121 (.L_HI(net121));
 sg13g2_tiehi _17638__122 (.L_HI(net122));
 sg13g2_tiehi _16395__123 (.L_HI(net123));
 sg13g2_tiehi _17637__124 (.L_HI(net124));
 sg13g2_tiehi _16394__125 (.L_HI(net125));
 sg13g2_tiehi _17636__126 (.L_HI(net126));
 sg13g2_tiehi _16393__127 (.L_HI(net127));
 sg13g2_tiehi _17635__128 (.L_HI(net128));
 sg13g2_tiehi _16392__129 (.L_HI(net129));
 sg13g2_tiehi _17634__130 (.L_HI(net130));
 sg13g2_tiehi _16391__131 (.L_HI(net131));
 sg13g2_tiehi _17633__132 (.L_HI(net132));
 sg13g2_tiehi _16390__133 (.L_HI(net133));
 sg13g2_tiehi _17632__134 (.L_HI(net134));
 sg13g2_tiehi _16389__135 (.L_HI(net135));
 sg13g2_tiehi _17631__136 (.L_HI(net136));
 sg13g2_tiehi _16388__137 (.L_HI(net137));
 sg13g2_tiehi _17630__138 (.L_HI(net138));
 sg13g2_tiehi _16387__139 (.L_HI(net139));
 sg13g2_tiehi _17629__140 (.L_HI(net140));
 sg13g2_tiehi _16386__141 (.L_HI(net141));
 sg13g2_tiehi _17628__142 (.L_HI(net142));
 sg13g2_tiehi _16385__143 (.L_HI(net143));
 sg13g2_tiehi _17627__144 (.L_HI(net144));
 sg13g2_tiehi _16384__145 (.L_HI(net145));
 sg13g2_tiehi _17626__146 (.L_HI(net146));
 sg13g2_tiehi _16383__147 (.L_HI(net147));
 sg13g2_tiehi _17625__148 (.L_HI(net148));
 sg13g2_tiehi _16382__149 (.L_HI(net149));
 sg13g2_tiehi _17624__150 (.L_HI(net150));
 sg13g2_tiehi _16381__151 (.L_HI(net151));
 sg13g2_tiehi _17623__152 (.L_HI(net152));
 sg13g2_tiehi _16380__153 (.L_HI(net153));
 sg13g2_tiehi _16379__154 (.L_HI(net154));
 sg13g2_tiehi _16378__155 (.L_HI(net155));
 sg13g2_tiehi _16377__156 (.L_HI(net156));
 sg13g2_tiehi _16376__157 (.L_HI(net157));
 sg13g2_tiehi _17622__158 (.L_HI(net158));
 sg13g2_tiehi _16375__159 (.L_HI(net159));
 sg13g2_tiehi _17621__160 (.L_HI(net160));
 sg13g2_tiehi _16374__161 (.L_HI(net161));
 sg13g2_tiehi _17620__162 (.L_HI(net162));
 sg13g2_tiehi _16373__163 (.L_HI(net163));
 sg13g2_tiehi _17619__164 (.L_HI(net164));
 sg13g2_tiehi _16372__165 (.L_HI(net165));
 sg13g2_tiehi _17618__166 (.L_HI(net166));
 sg13g2_tiehi _16371__167 (.L_HI(net167));
 sg13g2_tiehi _17617__168 (.L_HI(net168));
 sg13g2_tiehi _16370__169 (.L_HI(net169));
 sg13g2_tiehi _17616__170 (.L_HI(net170));
 sg13g2_tiehi _16369__171 (.L_HI(net171));
 sg13g2_tiehi _17615__172 (.L_HI(net172));
 sg13g2_tiehi _16368__173 (.L_HI(net173));
 sg13g2_tiehi _17614__174 (.L_HI(net174));
 sg13g2_tiehi _16367__175 (.L_HI(net175));
 sg13g2_tiehi _17613__176 (.L_HI(net176));
 sg13g2_tiehi _16366__177 (.L_HI(net177));
 sg13g2_tiehi _17612__178 (.L_HI(net178));
 sg13g2_tiehi _16365__179 (.L_HI(net179));
 sg13g2_tiehi _17611__180 (.L_HI(net180));
 sg13g2_tiehi _16364__181 (.L_HI(net181));
 sg13g2_tiehi _17610__182 (.L_HI(net182));
 sg13g2_tiehi _16363__183 (.L_HI(net183));
 sg13g2_tiehi _17609__184 (.L_HI(net184));
 sg13g2_tiehi _16362__185 (.L_HI(net185));
 sg13g2_tiehi _17608__186 (.L_HI(net186));
 sg13g2_tiehi _16361__187 (.L_HI(net187));
 sg13g2_tiehi _17919__188 (.L_HI(net188));
 sg13g2_tiehi _16360__189 (.L_HI(net189));
 sg13g2_tiehi _17607__190 (.L_HI(net190));
 sg13g2_tiehi _16359__191 (.L_HI(net191));
 sg13g2_tiehi _18018__192 (.L_HI(net192));
 sg13g2_tiehi _16358__193 (.L_HI(net193));
 sg13g2_tiehi _17606__194 (.L_HI(net194));
 sg13g2_tiehi _16357__195 (.L_HI(net195));
 sg13g2_tiehi _17918__196 (.L_HI(net196));
 sg13g2_tiehi _16356__197 (.L_HI(net197));
 sg13g2_tiehi _17605__198 (.L_HI(net198));
 sg13g2_tiehi _16355__199 (.L_HI(net199));
 sg13g2_tiehi _18138__200 (.L_HI(net200));
 sg13g2_tiehi _16354__201 (.L_HI(net201));
 sg13g2_tiehi _17604__202 (.L_HI(net202));
 sg13g2_tiehi _16353__203 (.L_HI(net203));
 sg13g2_tiehi _17603__204 (.L_HI(net204));
 sg13g2_tiehi _16352__205 (.L_HI(net205));
 sg13g2_tiehi _17602__206 (.L_HI(net206));
 sg13g2_tiehi _16351__207 (.L_HI(net207));
 sg13g2_tiehi _17601__208 (.L_HI(net208));
 sg13g2_tiehi _16350__209 (.L_HI(net209));
 sg13g2_tiehi _17600__210 (.L_HI(net210));
 sg13g2_tiehi _16349__211 (.L_HI(net211));
 sg13g2_tiehi _17599__212 (.L_HI(net212));
 sg13g2_tiehi _16348__213 (.L_HI(net213));
 sg13g2_tiehi _17598__214 (.L_HI(net214));
 sg13g2_tiehi _16347__215 (.L_HI(net215));
 sg13g2_tiehi _17597__216 (.L_HI(net216));
 sg13g2_tiehi _16346__217 (.L_HI(net217));
 sg13g2_tiehi _17596__218 (.L_HI(net218));
 sg13g2_tiehi _16345__219 (.L_HI(net219));
 sg13g2_tiehi _17595__220 (.L_HI(net220));
 sg13g2_tiehi _16344__221 (.L_HI(net221));
 sg13g2_tiehi _17594__222 (.L_HI(net222));
 sg13g2_tiehi _16343__223 (.L_HI(net223));
 sg13g2_tiehi _17593__224 (.L_HI(net224));
 sg13g2_tiehi _16342__225 (.L_HI(net225));
 sg13g2_tiehi _16341__226 (.L_HI(net226));
 sg13g2_tiehi _17592__227 (.L_HI(net227));
 sg13g2_tiehi _16340__228 (.L_HI(net228));
 sg13g2_tiehi _17591__229 (.L_HI(net229));
 sg13g2_tiehi _16339__230 (.L_HI(net230));
 sg13g2_tiehi _17590__231 (.L_HI(net231));
 sg13g2_tiehi _16338__232 (.L_HI(net232));
 sg13g2_tiehi _17589__233 (.L_HI(net233));
 sg13g2_tiehi _16337__234 (.L_HI(net234));
 sg13g2_tiehi _17588__235 (.L_HI(net235));
 sg13g2_tiehi _16336__236 (.L_HI(net236));
 sg13g2_tiehi _17587__237 (.L_HI(net237));
 sg13g2_tiehi _16335__238 (.L_HI(net238));
 sg13g2_tiehi _17586__239 (.L_HI(net239));
 sg13g2_tiehi _16334__240 (.L_HI(net240));
 sg13g2_tiehi _17585__241 (.L_HI(net241));
 sg13g2_tiehi _16333__242 (.L_HI(net242));
 sg13g2_tiehi _17584__243 (.L_HI(net243));
 sg13g2_tiehi _16332__244 (.L_HI(net244));
 sg13g2_tiehi _17583__245 (.L_HI(net245));
 sg13g2_tiehi _16331__246 (.L_HI(net246));
 sg13g2_tiehi _17582__247 (.L_HI(net247));
 sg13g2_tiehi _16330__248 (.L_HI(net248));
 sg13g2_tiehi _17581__249 (.L_HI(net249));
 sg13g2_tiehi _16329__250 (.L_HI(net250));
 sg13g2_tiehi _17580__251 (.L_HI(net251));
 sg13g2_tiehi _16328__252 (.L_HI(net252));
 sg13g2_tiehi _17579__253 (.L_HI(net253));
 sg13g2_tiehi _16327__254 (.L_HI(net254));
 sg13g2_tiehi _17578__255 (.L_HI(net255));
 sg13g2_tiehi _16326__256 (.L_HI(net256));
 sg13g2_tiehi _17577__257 (.L_HI(net257));
 sg13g2_tiehi _16325__258 (.L_HI(net258));
 sg13g2_tiehi _17576__259 (.L_HI(net259));
 sg13g2_tiehi _17575__260 (.L_HI(net260));
 sg13g2_tiehi _17574__261 (.L_HI(net261));
 sg13g2_tiehi _17573__262 (.L_HI(net262));
 sg13g2_tiehi _17572__263 (.L_HI(net263));
 sg13g2_tiehi _17571__264 (.L_HI(net264));
 sg13g2_tiehi _17570__265 (.L_HI(net265));
 sg13g2_tiehi _17569__266 (.L_HI(net266));
 sg13g2_tiehi _17568__267 (.L_HI(net267));
 sg13g2_tiehi _17567__268 (.L_HI(net268));
 sg13g2_tiehi _17566__269 (.L_HI(net269));
 sg13g2_tiehi _17565__270 (.L_HI(net270));
 sg13g2_tiehi _17564__271 (.L_HI(net271));
 sg13g2_tiehi _17917__272 (.L_HI(net272));
 sg13g2_tiehi _17563__273 (.L_HI(net273));
 sg13g2_tiehi _18017__274 (.L_HI(net274));
 sg13g2_tiehi _17550__275 (.L_HI(net275));
 sg13g2_tiehi _17916__276 (.L_HI(net276));
 sg13g2_tiehi _17549__277 (.L_HI(net277));
 sg13g2_tiehi _18067__278 (.L_HI(net278));
 sg13g2_tiehi _17548__279 (.L_HI(net279));
 sg13g2_tiehi _17915__280 (.L_HI(net280));
 sg13g2_tiehi _17547__281 (.L_HI(net281));
 sg13g2_tiehi _18016__282 (.L_HI(net282));
 sg13g2_tiehi _17546__283 (.L_HI(net283));
 sg13g2_tiehi _17914__284 (.L_HI(net284));
 sg13g2_tiehi _17545__285 (.L_HI(net285));
 sg13g2_tiehi _18092__286 (.L_HI(net286));
 sg13g2_tiehi _17544__287 (.L_HI(net287));
 sg13g2_tiehi _17913__288 (.L_HI(net288));
 sg13g2_tiehi _17543__289 (.L_HI(net289));
 sg13g2_tiehi _18015__290 (.L_HI(net290));
 sg13g2_tiehi _17542__291 (.L_HI(net291));
 sg13g2_tiehi _17912__292 (.L_HI(net292));
 sg13g2_tiehi _17541__293 (.L_HI(net293));
 sg13g2_tiehi _18066__294 (.L_HI(net294));
 sg13g2_tiehi _17540__295 (.L_HI(net295));
 sg13g2_tiehi _17911__296 (.L_HI(net296));
 sg13g2_tiehi _16444__297 (.L_HI(net297));
 sg13g2_tiehi _17539__298 (.L_HI(net298));
 sg13g2_tiehi _18014__299 (.L_HI(net299));
 sg13g2_tiehi _17538__300 (.L_HI(net300));
 sg13g2_tiehi _17910__301 (.L_HI(net301));
 sg13g2_tiehi _17537__302 (.L_HI(net302));
 sg13g2_tiehi _18147__303 (.L_HI(net303));
 sg13g2_tiehi _17536__304 (.L_HI(net304));
 sg13g2_tiehi _17909__305 (.L_HI(net305));
 sg13g2_tiehi _17535__306 (.L_HI(net306));
 sg13g2_tiehi _18013__307 (.L_HI(net307));
 sg13g2_tiehi _17534__308 (.L_HI(net308));
 sg13g2_tiehi _17533__309 (.L_HI(net309));
 sg13g2_tiehi _17908__310 (.L_HI(net310));
 sg13g2_tiehi _17532__311 (.L_HI(net311));
 sg13g2_tiehi _18065__312 (.L_HI(net312));
 sg13g2_tiehi _17531__313 (.L_HI(net313));
 sg13g2_tiehi _17907__314 (.L_HI(net314));
 sg13g2_tiehi _17530__315 (.L_HI(net315));
 sg13g2_tiehi _18012__316 (.L_HI(net316));
 sg13g2_tiehi _17529__317 (.L_HI(net317));
 sg13g2_tiehi _17906__318 (.L_HI(net318));
 sg13g2_tiehi _17528__319 (.L_HI(net319));
 sg13g2_tiehi _18091__320 (.L_HI(net320));
 sg13g2_tiehi _17527__321 (.L_HI(net321));
 sg13g2_tiehi _17905__322 (.L_HI(net322));
 sg13g2_tiehi _17526__323 (.L_HI(net323));
 sg13g2_tiehi _18011__324 (.L_HI(net324));
 sg13g2_tiehi _17525__325 (.L_HI(net325));
 sg13g2_tiehi _17904__326 (.L_HI(net326));
 sg13g2_tiehi _17524__327 (.L_HI(net327));
 sg13g2_tiehi _18064__328 (.L_HI(net328));
 sg13g2_tiehi _17523__329 (.L_HI(net329));
 sg13g2_tiehi _17903__330 (.L_HI(net330));
 sg13g2_tiehi _17522__331 (.L_HI(net331));
 sg13g2_tiehi _18010__332 (.L_HI(net332));
 sg13g2_tiehi _17521__333 (.L_HI(net333));
 sg13g2_tiehi _17902__334 (.L_HI(net334));
 sg13g2_tiehi _17520__335 (.L_HI(net335));
 sg13g2_tiehi _18137__336 (.L_HI(net336));
 sg13g2_tiehi _17519__337 (.L_HI(net337));
 sg13g2_tiehi _17901__338 (.L_HI(net338));
 sg13g2_tiehi _17518__339 (.L_HI(net339));
 sg13g2_tiehi _18009__340 (.L_HI(net340));
 sg13g2_tiehi _17517__341 (.L_HI(net341));
 sg13g2_tiehi _17900__342 (.L_HI(net342));
 sg13g2_tiehi _17516__343 (.L_HI(net343));
 sg13g2_tiehi _18063__344 (.L_HI(net344));
 sg13g2_tiehi _17515__345 (.L_HI(net345));
 sg13g2_tiehi _17899__346 (.L_HI(net346));
 sg13g2_tiehi _17514__347 (.L_HI(net347));
 sg13g2_tiehi _18008__348 (.L_HI(net348));
 sg13g2_tiehi _17513__349 (.L_HI(net349));
 sg13g2_tiehi _17898__350 (.L_HI(net350));
 sg13g2_tiehi _17512__351 (.L_HI(net351));
 sg13g2_tiehi _18090__352 (.L_HI(net352));
 sg13g2_tiehi _17511__353 (.L_HI(net353));
 sg13g2_tiehi _17897__354 (.L_HI(net354));
 sg13g2_tiehi _17510__355 (.L_HI(net355));
 sg13g2_tiehi _18007__356 (.L_HI(net356));
 sg13g2_tiehi _17509__357 (.L_HI(net357));
 sg13g2_tiehi _17896__358 (.L_HI(net358));
 sg13g2_tiehi _17508__359 (.L_HI(net359));
 sg13g2_tiehi _18062__360 (.L_HI(net360));
 sg13g2_tiehi _17507__361 (.L_HI(net361));
 sg13g2_tiehi _17895__362 (.L_HI(net362));
 sg13g2_tiehi _17506__363 (.L_HI(net363));
 sg13g2_tiehi _18006__364 (.L_HI(net364));
 sg13g2_tiehi _17505__365 (.L_HI(net365));
 sg13g2_tiehi _17894__366 (.L_HI(net366));
 sg13g2_tiehi _17504__367 (.L_HI(net367));
 sg13g2_tiehi _18144__368 (.L_HI(net368));
 sg13g2_tiehi _17503__369 (.L_HI(net369));
 sg13g2_tiehi _17893__370 (.L_HI(net370));
 sg13g2_tiehi _17502__371 (.L_HI(net371));
 sg13g2_tiehi _18005__372 (.L_HI(net372));
 sg13g2_tiehi _17501__373 (.L_HI(net373));
 sg13g2_tiehi _17892__374 (.L_HI(net374));
 sg13g2_tiehi _16620__375 (.L_HI(net375));
 sg13g2_tiehi _16698__376 (.L_HI(net376));
 sg13g2_tiehi _16699__377 (.L_HI(net377));
 sg13g2_tiehi _16700__378 (.L_HI(net378));
 sg13g2_tiehi _16701__379 (.L_HI(net379));
 sg13g2_tiehi _16702__380 (.L_HI(net380));
 sg13g2_tiehi _16703__381 (.L_HI(net381));
 sg13g2_tiehi _16704__382 (.L_HI(net382));
 sg13g2_tiehi _16705__383 (.L_HI(net383));
 sg13g2_tiehi _16706__384 (.L_HI(net384));
 sg13g2_tiehi _16707__385 (.L_HI(net385));
 sg13g2_tiehi _16708__386 (.L_HI(net386));
 sg13g2_tiehi _16709__387 (.L_HI(net387));
 sg13g2_tiehi _16710__388 (.L_HI(net388));
 sg13g2_tiehi _16711__389 (.L_HI(net389));
 sg13g2_tiehi _16712__390 (.L_HI(net390));
 sg13g2_tiehi _16713__391 (.L_HI(net391));
 sg13g2_tiehi _16714__392 (.L_HI(net392));
 sg13g2_tiehi _16715__393 (.L_HI(net393));
 sg13g2_tiehi _16716__394 (.L_HI(net394));
 sg13g2_tiehi _16717__395 (.L_HI(net395));
 sg13g2_tiehi _16718__396 (.L_HI(net396));
 sg13g2_tiehi _16719__397 (.L_HI(net397));
 sg13g2_tiehi _16720__398 (.L_HI(net398));
 sg13g2_tiehi _16721__399 (.L_HI(net399));
 sg13g2_tiehi _16722__400 (.L_HI(net400));
 sg13g2_tiehi _16723__401 (.L_HI(net401));
 sg13g2_tiehi _16724__402 (.L_HI(net402));
 sg13g2_tiehi _17500__403 (.L_HI(net403));
 sg13g2_tiehi _18061__404 (.L_HI(net404));
 sg13g2_tiehi _17499__405 (.L_HI(net405));
 sg13g2_tiehi _17891__406 (.L_HI(net406));
 sg13g2_tiehi _17498__407 (.L_HI(net407));
 sg13g2_tiehi _16725__408 (.L_HI(net408));
 sg13g2_tiehi _16731__409 (.L_HI(net409));
 sg13g2_tiehi _16732__410 (.L_HI(net410));
 sg13g2_tiehi _16733__411 (.L_HI(net411));
 sg13g2_tiehi _16734__412 (.L_HI(net412));
 sg13g2_tiehi _16735__413 (.L_HI(net413));
 sg13g2_tiehi _16736__414 (.L_HI(net414));
 sg13g2_tiehi _16737__415 (.L_HI(net415));
 sg13g2_tiehi _16738__416 (.L_HI(net416));
 sg13g2_tiehi _16739__417 (.L_HI(net417));
 sg13g2_tiehi _16740__418 (.L_HI(net418));
 sg13g2_tiehi _16741__419 (.L_HI(net419));
 sg13g2_tiehi _16742__420 (.L_HI(net420));
 sg13g2_tiehi _16743__421 (.L_HI(net421));
 sg13g2_tiehi _16744__422 (.L_HI(net422));
 sg13g2_tiehi _16745__423 (.L_HI(net423));
 sg13g2_tiehi _16746__424 (.L_HI(net424));
 sg13g2_tiehi _16747__425 (.L_HI(net425));
 sg13g2_tiehi _16748__426 (.L_HI(net426));
 sg13g2_tiehi _16749__427 (.L_HI(net427));
 sg13g2_tiehi _16750__428 (.L_HI(net428));
 sg13g2_tiehi _16751__429 (.L_HI(net429));
 sg13g2_tiehi _16752__430 (.L_HI(net430));
 sg13g2_tiehi _16753__431 (.L_HI(net431));
 sg13g2_tiehi _16754__432 (.L_HI(net432));
 sg13g2_tiehi _16755__433 (.L_HI(net433));
 sg13g2_tiehi _16756__434 (.L_HI(net434));
 sg13g2_tiehi _16757__435 (.L_HI(net435));
 sg13g2_tiehi _18004__436 (.L_HI(net436));
 sg13g2_tiehi _17497__437 (.L_HI(net437));
 sg13g2_tiehi _17890__438 (.L_HI(net438));
 sg13g2_tiehi _17496__439 (.L_HI(net439));
 sg13g2_tiehi _18089__440 (.L_HI(net440));
 sg13g2_tiehi _17495__441 (.L_HI(net441));
 sg13g2_tiehi _16758__442 (.L_HI(net442));
 sg13g2_tiehi _16765__443 (.L_HI(net443));
 sg13g2_tiehi _16766__444 (.L_HI(net444));
 sg13g2_tiehi _16767__445 (.L_HI(net445));
 sg13g2_tiehi _16768__446 (.L_HI(net446));
 sg13g2_tiehi _16769__447 (.L_HI(net447));
 sg13g2_tiehi _16770__448 (.L_HI(net448));
 sg13g2_tiehi _16771__449 (.L_HI(net449));
 sg13g2_tiehi _16772__450 (.L_HI(net450));
 sg13g2_tiehi _16773__451 (.L_HI(net451));
 sg13g2_tiehi _16774__452 (.L_HI(net452));
 sg13g2_tiehi _16775__453 (.L_HI(net453));
 sg13g2_tiehi _16776__454 (.L_HI(net454));
 sg13g2_tiehi _16777__455 (.L_HI(net455));
 sg13g2_tiehi _16778__456 (.L_HI(net456));
 sg13g2_tiehi _16779__457 (.L_HI(net457));
 sg13g2_tiehi _16780__458 (.L_HI(net458));
 sg13g2_tiehi _16781__459 (.L_HI(net459));
 sg13g2_tiehi _16782__460 (.L_HI(net460));
 sg13g2_tiehi _16783__461 (.L_HI(net461));
 sg13g2_tiehi _16784__462 (.L_HI(net462));
 sg13g2_tiehi _16785__463 (.L_HI(net463));
 sg13g2_tiehi _16786__464 (.L_HI(net464));
 sg13g2_tiehi _16787__465 (.L_HI(net465));
 sg13g2_tiehi _16788__466 (.L_HI(net466));
 sg13g2_tiehi _16789__467 (.L_HI(net467));
 sg13g2_tiehi _16790__468 (.L_HI(net468));
 sg13g2_tiehi _16791__469 (.L_HI(net469));
 sg13g2_tiehi _16792__470 (.L_HI(net470));
 sg13g2_tiehi _16793__471 (.L_HI(net471));
 sg13g2_tiehi _16794__472 (.L_HI(net472));
 sg13g2_tiehi _16795__473 (.L_HI(net473));
 sg13g2_tiehi _16796__474 (.L_HI(net474));
 sg13g2_tiehi _16797__475 (.L_HI(net475));
 sg13g2_tiehi _16798__476 (.L_HI(net476));
 sg13g2_tiehi _16799__477 (.L_HI(net477));
 sg13g2_tiehi _16800__478 (.L_HI(net478));
 sg13g2_tiehi _16801__479 (.L_HI(net479));
 sg13g2_tiehi _16802__480 (.L_HI(net480));
 sg13g2_tiehi _16803__481 (.L_HI(net481));
 sg13g2_tiehi _16804__482 (.L_HI(net482));
 sg13g2_tiehi _16805__483 (.L_HI(net483));
 sg13g2_tiehi _16806__484 (.L_HI(net484));
 sg13g2_tiehi _16807__485 (.L_HI(net485));
 sg13g2_tiehi _16808__486 (.L_HI(net486));
 sg13g2_tiehi _16809__487 (.L_HI(net487));
 sg13g2_tiehi _16810__488 (.L_HI(net488));
 sg13g2_tiehi _16811__489 (.L_HI(net489));
 sg13g2_tiehi _16812__490 (.L_HI(net490));
 sg13g2_tiehi _16813__491 (.L_HI(net491));
 sg13g2_tiehi _16814__492 (.L_HI(net492));
 sg13g2_tiehi _16815__493 (.L_HI(net493));
 sg13g2_tiehi _16816__494 (.L_HI(net494));
 sg13g2_tiehi _16817__495 (.L_HI(net495));
 sg13g2_tiehi _16818__496 (.L_HI(net496));
 sg13g2_tiehi _16819__497 (.L_HI(net497));
 sg13g2_tiehi _16820__498 (.L_HI(net498));
 sg13g2_tiehi _16821__499 (.L_HI(net499));
 sg13g2_tiehi _16822__500 (.L_HI(net500));
 sg13g2_tiehi _16823__501 (.L_HI(net501));
 sg13g2_tiehi _16824__502 (.L_HI(net502));
 sg13g2_tiehi _16825__503 (.L_HI(net503));
 sg13g2_tiehi _16826__504 (.L_HI(net504));
 sg13g2_tiehi _16827__505 (.L_HI(net505));
 sg13g2_tiehi _16828__506 (.L_HI(net506));
 sg13g2_tiehi _16829__507 (.L_HI(net507));
 sg13g2_tiehi _16830__508 (.L_HI(net508));
 sg13g2_tiehi _16831__509 (.L_HI(net509));
 sg13g2_tiehi _16832__510 (.L_HI(net510));
 sg13g2_tiehi _16833__511 (.L_HI(net511));
 sg13g2_tiehi _16834__512 (.L_HI(net512));
 sg13g2_tiehi _16835__513 (.L_HI(net513));
 sg13g2_tiehi _16836__514 (.L_HI(net514));
 sg13g2_tiehi _16837__515 (.L_HI(net515));
 sg13g2_tiehi _16838__516 (.L_HI(net516));
 sg13g2_tiehi _16839__517 (.L_HI(net517));
 sg13g2_tiehi _16840__518 (.L_HI(net518));
 sg13g2_tiehi _16841__519 (.L_HI(net519));
 sg13g2_tiehi _16842__520 (.L_HI(net520));
 sg13g2_tiehi _16843__521 (.L_HI(net521));
 sg13g2_tiehi _16844__522 (.L_HI(net522));
 sg13g2_tiehi _16845__523 (.L_HI(net523));
 sg13g2_tiehi _16846__524 (.L_HI(net524));
 sg13g2_tiehi _16847__525 (.L_HI(net525));
 sg13g2_tiehi _16848__526 (.L_HI(net526));
 sg13g2_tiehi _16849__527 (.L_HI(net527));
 sg13g2_tiehi _16850__528 (.L_HI(net528));
 sg13g2_tiehi _16851__529 (.L_HI(net529));
 sg13g2_tiehi _16852__530 (.L_HI(net530));
 sg13g2_tiehi _16853__531 (.L_HI(net531));
 sg13g2_tiehi _16854__532 (.L_HI(net532));
 sg13g2_tiehi _16855__533 (.L_HI(net533));
 sg13g2_tiehi _16856__534 (.L_HI(net534));
 sg13g2_tiehi _16857__535 (.L_HI(net535));
 sg13g2_tiehi _16858__536 (.L_HI(net536));
 sg13g2_tiehi _16859__537 (.L_HI(net537));
 sg13g2_tiehi _16860__538 (.L_HI(net538));
 sg13g2_tiehi _16861__539 (.L_HI(net539));
 sg13g2_tiehi _16862__540 (.L_HI(net540));
 sg13g2_tiehi _16863__541 (.L_HI(net541));
 sg13g2_tiehi _16864__542 (.L_HI(net542));
 sg13g2_tiehi _16865__543 (.L_HI(net543));
 sg13g2_tiehi _16866__544 (.L_HI(net544));
 sg13g2_tiehi _16867__545 (.L_HI(net545));
 sg13g2_tiehi _16868__546 (.L_HI(net546));
 sg13g2_tiehi _16869__547 (.L_HI(net547));
 sg13g2_tiehi _16870__548 (.L_HI(net548));
 sg13g2_tiehi _16871__549 (.L_HI(net549));
 sg13g2_tiehi _16872__550 (.L_HI(net550));
 sg13g2_tiehi _16873__551 (.L_HI(net551));
 sg13g2_tiehi _16874__552 (.L_HI(net552));
 sg13g2_tiehi _16875__553 (.L_HI(net553));
 sg13g2_tiehi _16876__554 (.L_HI(net554));
 sg13g2_tiehi _16877__555 (.L_HI(net555));
 sg13g2_tiehi _16878__556 (.L_HI(net556));
 sg13g2_tiehi _16879__557 (.L_HI(net557));
 sg13g2_tiehi _16880__558 (.L_HI(net558));
 sg13g2_tiehi _16881__559 (.L_HI(net559));
 sg13g2_tiehi _16882__560 (.L_HI(net560));
 sg13g2_tiehi _16883__561 (.L_HI(net561));
 sg13g2_tiehi _16884__562 (.L_HI(net562));
 sg13g2_tiehi _16885__563 (.L_HI(net563));
 sg13g2_tiehi _16886__564 (.L_HI(net564));
 sg13g2_tiehi _16887__565 (.L_HI(net565));
 sg13g2_tiehi _16888__566 (.L_HI(net566));
 sg13g2_tiehi _16889__567 (.L_HI(net567));
 sg13g2_tiehi _16890__568 (.L_HI(net568));
 sg13g2_tiehi _16891__569 (.L_HI(net569));
 sg13g2_tiehi _16892__570 (.L_HI(net570));
 sg13g2_tiehi _16893__571 (.L_HI(net571));
 sg13g2_tiehi _16894__572 (.L_HI(net572));
 sg13g2_tiehi _16895__573 (.L_HI(net573));
 sg13g2_tiehi _16896__574 (.L_HI(net574));
 sg13g2_tiehi _16897__575 (.L_HI(net575));
 sg13g2_tiehi _16898__576 (.L_HI(net576));
 sg13g2_tiehi _16899__577 (.L_HI(net577));
 sg13g2_tiehi _16900__578 (.L_HI(net578));
 sg13g2_tiehi _16901__579 (.L_HI(net579));
 sg13g2_tiehi _16902__580 (.L_HI(net580));
 sg13g2_tiehi _16903__581 (.L_HI(net581));
 sg13g2_tiehi _16904__582 (.L_HI(net582));
 sg13g2_tiehi _16905__583 (.L_HI(net583));
 sg13g2_tiehi _16906__584 (.L_HI(net584));
 sg13g2_tiehi _16907__585 (.L_HI(net585));
 sg13g2_tiehi _16908__586 (.L_HI(net586));
 sg13g2_tiehi _16909__587 (.L_HI(net587));
 sg13g2_tiehi _16910__588 (.L_HI(net588));
 sg13g2_tiehi _16911__589 (.L_HI(net589));
 sg13g2_tiehi _16912__590 (.L_HI(net590));
 sg13g2_tiehi _16913__591 (.L_HI(net591));
 sg13g2_tiehi _16914__592 (.L_HI(net592));
 sg13g2_tiehi _16915__593 (.L_HI(net593));
 sg13g2_tiehi _16916__594 (.L_HI(net594));
 sg13g2_tiehi _16917__595 (.L_HI(net595));
 sg13g2_tiehi _16918__596 (.L_HI(net596));
 sg13g2_tiehi _16919__597 (.L_HI(net597));
 sg13g2_tiehi _16920__598 (.L_HI(net598));
 sg13g2_tiehi _16921__599 (.L_HI(net599));
 sg13g2_tiehi _16922__600 (.L_HI(net600));
 sg13g2_tiehi _16923__601 (.L_HI(net601));
 sg13g2_tiehi _16924__602 (.L_HI(net602));
 sg13g2_tiehi _16925__603 (.L_HI(net603));
 sg13g2_tiehi _16926__604 (.L_HI(net604));
 sg13g2_tiehi _16927__605 (.L_HI(net605));
 sg13g2_tiehi _16928__606 (.L_HI(net606));
 sg13g2_tiehi _16929__607 (.L_HI(net607));
 sg13g2_tiehi _16930__608 (.L_HI(net608));
 sg13g2_tiehi _16931__609 (.L_HI(net609));
 sg13g2_tiehi _16932__610 (.L_HI(net610));
 sg13g2_tiehi _16933__611 (.L_HI(net611));
 sg13g2_tiehi _16934__612 (.L_HI(net612));
 sg13g2_tiehi _16935__613 (.L_HI(net613));
 sg13g2_tiehi _16936__614 (.L_HI(net614));
 sg13g2_tiehi _16937__615 (.L_HI(net615));
 sg13g2_tiehi _16938__616 (.L_HI(net616));
 sg13g2_tiehi _16939__617 (.L_HI(net617));
 sg13g2_tiehi _16940__618 (.L_HI(net618));
 sg13g2_tiehi _16941__619 (.L_HI(net619));
 sg13g2_tiehi _16942__620 (.L_HI(net620));
 sg13g2_tiehi _16943__621 (.L_HI(net621));
 sg13g2_tiehi _16944__622 (.L_HI(net622));
 sg13g2_tiehi _16945__623 (.L_HI(net623));
 sg13g2_tiehi _16946__624 (.L_HI(net624));
 sg13g2_tiehi _16947__625 (.L_HI(net625));
 sg13g2_tiehi _16948__626 (.L_HI(net626));
 sg13g2_tiehi _16949__627 (.L_HI(net627));
 sg13g2_tiehi _16950__628 (.L_HI(net628));
 sg13g2_tiehi _16951__629 (.L_HI(net629));
 sg13g2_tiehi _16952__630 (.L_HI(net630));
 sg13g2_tiehi _16953__631 (.L_HI(net631));
 sg13g2_tiehi _16954__632 (.L_HI(net632));
 sg13g2_tiehi _16955__633 (.L_HI(net633));
 sg13g2_tiehi _16956__634 (.L_HI(net634));
 sg13g2_tiehi _16957__635 (.L_HI(net635));
 sg13g2_tiehi _16958__636 (.L_HI(net636));
 sg13g2_tiehi _16959__637 (.L_HI(net637));
 sg13g2_tiehi _16960__638 (.L_HI(net638));
 sg13g2_tiehi _16961__639 (.L_HI(net639));
 sg13g2_tiehi _16962__640 (.L_HI(net640));
 sg13g2_tiehi _16963__641 (.L_HI(net641));
 sg13g2_tiehi _16964__642 (.L_HI(net642));
 sg13g2_tiehi _16965__643 (.L_HI(net643));
 sg13g2_tiehi _16966__644 (.L_HI(net644));
 sg13g2_tiehi _16967__645 (.L_HI(net645));
 sg13g2_tiehi _16968__646 (.L_HI(net646));
 sg13g2_tiehi _16969__647 (.L_HI(net647));
 sg13g2_tiehi _16970__648 (.L_HI(net648));
 sg13g2_tiehi _16971__649 (.L_HI(net649));
 sg13g2_tiehi _16972__650 (.L_HI(net650));
 sg13g2_tiehi _16973__651 (.L_HI(net651));
 sg13g2_tiehi _16974__652 (.L_HI(net652));
 sg13g2_tiehi _16975__653 (.L_HI(net653));
 sg13g2_tiehi _16976__654 (.L_HI(net654));
 sg13g2_tiehi _16977__655 (.L_HI(net655));
 sg13g2_tiehi _16978__656 (.L_HI(net656));
 sg13g2_tiehi _16979__657 (.L_HI(net657));
 sg13g2_tiehi _16980__658 (.L_HI(net658));
 sg13g2_tiehi _16981__659 (.L_HI(net659));
 sg13g2_tiehi _16982__660 (.L_HI(net660));
 sg13g2_tiehi _16983__661 (.L_HI(net661));
 sg13g2_tiehi _16984__662 (.L_HI(net662));
 sg13g2_tiehi _16985__663 (.L_HI(net663));
 sg13g2_tiehi _16986__664 (.L_HI(net664));
 sg13g2_tiehi _16987__665 (.L_HI(net665));
 sg13g2_tiehi _16988__666 (.L_HI(net666));
 sg13g2_tiehi _16989__667 (.L_HI(net667));
 sg13g2_tiehi _16990__668 (.L_HI(net668));
 sg13g2_tiehi _16991__669 (.L_HI(net669));
 sg13g2_tiehi _16992__670 (.L_HI(net670));
 sg13g2_tiehi _16993__671 (.L_HI(net671));
 sg13g2_tiehi _16994__672 (.L_HI(net672));
 sg13g2_tiehi _16995__673 (.L_HI(net673));
 sg13g2_tiehi _16996__674 (.L_HI(net674));
 sg13g2_tiehi _16997__675 (.L_HI(net675));
 sg13g2_tiehi _16998__676 (.L_HI(net676));
 sg13g2_tiehi _16999__677 (.L_HI(net677));
 sg13g2_tiehi _17000__678 (.L_HI(net678));
 sg13g2_tiehi _17001__679 (.L_HI(net679));
 sg13g2_tiehi _17002__680 (.L_HI(net680));
 sg13g2_tiehi _17003__681 (.L_HI(net681));
 sg13g2_tiehi _17004__682 (.L_HI(net682));
 sg13g2_tiehi _17005__683 (.L_HI(net683));
 sg13g2_tiehi _17006__684 (.L_HI(net684));
 sg13g2_tiehi _17007__685 (.L_HI(net685));
 sg13g2_tiehi _17008__686 (.L_HI(net686));
 sg13g2_tiehi _17009__687 (.L_HI(net687));
 sg13g2_tiehi _17010__688 (.L_HI(net688));
 sg13g2_tiehi _17011__689 (.L_HI(net689));
 sg13g2_tiehi _17012__690 (.L_HI(net690));
 sg13g2_tiehi _17013__691 (.L_HI(net691));
 sg13g2_tiehi _17014__692 (.L_HI(net692));
 sg13g2_tiehi _17015__693 (.L_HI(net693));
 sg13g2_tiehi _17016__694 (.L_HI(net694));
 sg13g2_tiehi _17017__695 (.L_HI(net695));
 sg13g2_tiehi _17018__696 (.L_HI(net696));
 sg13g2_tiehi _17019__697 (.L_HI(net697));
 sg13g2_tiehi _17020__698 (.L_HI(net698));
 sg13g2_tiehi _17021__699 (.L_HI(net699));
 sg13g2_tiehi _17022__700 (.L_HI(net700));
 sg13g2_tiehi _17023__701 (.L_HI(net701));
 sg13g2_tiehi _17024__702 (.L_HI(net702));
 sg13g2_tiehi _17025__703 (.L_HI(net703));
 sg13g2_tiehi _17026__704 (.L_HI(net704));
 sg13g2_tiehi _17027__705 (.L_HI(net705));
 sg13g2_tiehi _17028__706 (.L_HI(net706));
 sg13g2_tiehi _17029__707 (.L_HI(net707));
 sg13g2_tiehi _17030__708 (.L_HI(net708));
 sg13g2_tiehi _17031__709 (.L_HI(net709));
 sg13g2_tiehi _17032__710 (.L_HI(net710));
 sg13g2_tiehi _17033__711 (.L_HI(net711));
 sg13g2_tiehi _17034__712 (.L_HI(net712));
 sg13g2_tiehi _17035__713 (.L_HI(net713));
 sg13g2_tiehi _17036__714 (.L_HI(net714));
 sg13g2_tiehi _17037__715 (.L_HI(net715));
 sg13g2_tiehi _17038__716 (.L_HI(net716));
 sg13g2_tiehi _17039__717 (.L_HI(net717));
 sg13g2_tiehi _17040__718 (.L_HI(net718));
 sg13g2_tiehi _17041__719 (.L_HI(net719));
 sg13g2_tiehi _17042__720 (.L_HI(net720));
 sg13g2_tiehi _17043__721 (.L_HI(net721));
 sg13g2_tiehi _17044__722 (.L_HI(net722));
 sg13g2_tiehi _17045__723 (.L_HI(net723));
 sg13g2_tiehi _17046__724 (.L_HI(net724));
 sg13g2_tiehi _17047__725 (.L_HI(net725));
 sg13g2_tiehi _17048__726 (.L_HI(net726));
 sg13g2_tiehi _17049__727 (.L_HI(net727));
 sg13g2_tiehi _17050__728 (.L_HI(net728));
 sg13g2_tiehi _17051__729 (.L_HI(net729));
 sg13g2_tiehi _17052__730 (.L_HI(net730));
 sg13g2_tiehi _17053__731 (.L_HI(net731));
 sg13g2_tiehi _17054__732 (.L_HI(net732));
 sg13g2_tiehi _17055__733 (.L_HI(net733));
 sg13g2_tiehi _17056__734 (.L_HI(net734));
 sg13g2_tiehi _17057__735 (.L_HI(net735));
 sg13g2_tiehi _17058__736 (.L_HI(net736));
 sg13g2_tiehi _17059__737 (.L_HI(net737));
 sg13g2_tiehi _17060__738 (.L_HI(net738));
 sg13g2_tiehi _17061__739 (.L_HI(net739));
 sg13g2_tiehi _17062__740 (.L_HI(net740));
 sg13g2_tiehi _17063__741 (.L_HI(net741));
 sg13g2_tiehi _17064__742 (.L_HI(net742));
 sg13g2_tiehi _17065__743 (.L_HI(net743));
 sg13g2_tiehi _17066__744 (.L_HI(net744));
 sg13g2_tiehi _17067__745 (.L_HI(net745));
 sg13g2_tiehi _17068__746 (.L_HI(net746));
 sg13g2_tiehi _17069__747 (.L_HI(net747));
 sg13g2_tiehi _17070__748 (.L_HI(net748));
 sg13g2_tiehi _17071__749 (.L_HI(net749));
 sg13g2_tiehi _17072__750 (.L_HI(net750));
 sg13g2_tiehi _17073__751 (.L_HI(net751));
 sg13g2_tiehi _17074__752 (.L_HI(net752));
 sg13g2_tiehi _17075__753 (.L_HI(net753));
 sg13g2_tiehi _17076__754 (.L_HI(net754));
 sg13g2_tiehi _17077__755 (.L_HI(net755));
 sg13g2_tiehi _17078__756 (.L_HI(net756));
 sg13g2_tiehi _17079__757 (.L_HI(net757));
 sg13g2_tiehi _17080__758 (.L_HI(net758));
 sg13g2_tiehi _17081__759 (.L_HI(net759));
 sg13g2_tiehi _17082__760 (.L_HI(net760));
 sg13g2_tiehi _17083__761 (.L_HI(net761));
 sg13g2_tiehi _17084__762 (.L_HI(net762));
 sg13g2_tiehi _17085__763 (.L_HI(net763));
 sg13g2_tiehi _17086__764 (.L_HI(net764));
 sg13g2_tiehi _17087__765 (.L_HI(net765));
 sg13g2_tiehi _17088__766 (.L_HI(net766));
 sg13g2_tiehi _17089__767 (.L_HI(net767));
 sg13g2_tiehi _17090__768 (.L_HI(net768));
 sg13g2_tiehi _17091__769 (.L_HI(net769));
 sg13g2_tiehi _17092__770 (.L_HI(net770));
 sg13g2_tiehi _17093__771 (.L_HI(net771));
 sg13g2_tiehi _17094__772 (.L_HI(net772));
 sg13g2_tiehi _17095__773 (.L_HI(net773));
 sg13g2_tiehi _17096__774 (.L_HI(net774));
 sg13g2_tiehi _17097__775 (.L_HI(net775));
 sg13g2_tiehi _17098__776 (.L_HI(net776));
 sg13g2_tiehi _17099__777 (.L_HI(net777));
 sg13g2_tiehi _17100__778 (.L_HI(net778));
 sg13g2_tiehi _17101__779 (.L_HI(net779));
 sg13g2_tiehi _17102__780 (.L_HI(net780));
 sg13g2_tiehi _17103__781 (.L_HI(net781));
 sg13g2_tiehi _17104__782 (.L_HI(net782));
 sg13g2_tiehi _17105__783 (.L_HI(net783));
 sg13g2_tiehi _17106__784 (.L_HI(net784));
 sg13g2_tiehi _17107__785 (.L_HI(net785));
 sg13g2_tiehi _17108__786 (.L_HI(net786));
 sg13g2_tiehi _17109__787 (.L_HI(net787));
 sg13g2_tiehi _17110__788 (.L_HI(net788));
 sg13g2_tiehi _17111__789 (.L_HI(net789));
 sg13g2_tiehi _17112__790 (.L_HI(net790));
 sg13g2_tiehi _17113__791 (.L_HI(net791));
 sg13g2_tiehi _17114__792 (.L_HI(net792));
 sg13g2_tiehi _17115__793 (.L_HI(net793));
 sg13g2_tiehi _17116__794 (.L_HI(net794));
 sg13g2_tiehi _17117__795 (.L_HI(net795));
 sg13g2_tiehi _17118__796 (.L_HI(net796));
 sg13g2_tiehi _17119__797 (.L_HI(net797));
 sg13g2_tiehi _17120__798 (.L_HI(net798));
 sg13g2_tiehi _17121__799 (.L_HI(net799));
 sg13g2_tiehi _17122__800 (.L_HI(net800));
 sg13g2_tiehi _17123__801 (.L_HI(net801));
 sg13g2_tiehi _17124__802 (.L_HI(net802));
 sg13g2_tiehi _17125__803 (.L_HI(net803));
 sg13g2_tiehi _17126__804 (.L_HI(net804));
 sg13g2_tiehi _17127__805 (.L_HI(net805));
 sg13g2_tiehi _17128__806 (.L_HI(net806));
 sg13g2_tiehi _17129__807 (.L_HI(net807));
 sg13g2_tiehi _17130__808 (.L_HI(net808));
 sg13g2_tiehi _17131__809 (.L_HI(net809));
 sg13g2_tiehi _17132__810 (.L_HI(net810));
 sg13g2_tiehi _17133__811 (.L_HI(net811));
 sg13g2_tiehi _17134__812 (.L_HI(net812));
 sg13g2_tiehi _17135__813 (.L_HI(net813));
 sg13g2_tiehi _17136__814 (.L_HI(net814));
 sg13g2_tiehi _17137__815 (.L_HI(net815));
 sg13g2_tiehi _17138__816 (.L_HI(net816));
 sg13g2_tiehi _17139__817 (.L_HI(net817));
 sg13g2_tiehi _17140__818 (.L_HI(net818));
 sg13g2_tiehi _17141__819 (.L_HI(net819));
 sg13g2_tiehi _17142__820 (.L_HI(net820));
 sg13g2_tiehi _17143__821 (.L_HI(net821));
 sg13g2_tiehi _17144__822 (.L_HI(net822));
 sg13g2_tiehi _17145__823 (.L_HI(net823));
 sg13g2_tiehi _17146__824 (.L_HI(net824));
 sg13g2_tiehi _17147__825 (.L_HI(net825));
 sg13g2_tiehi _17148__826 (.L_HI(net826));
 sg13g2_tiehi _17149__827 (.L_HI(net827));
 sg13g2_tiehi _17150__828 (.L_HI(net828));
 sg13g2_tiehi _17151__829 (.L_HI(net829));
 sg13g2_tiehi _17152__830 (.L_HI(net830));
 sg13g2_tiehi _17153__831 (.L_HI(net831));
 sg13g2_tiehi _17154__832 (.L_HI(net832));
 sg13g2_tiehi _17155__833 (.L_HI(net833));
 sg13g2_tiehi _17156__834 (.L_HI(net834));
 sg13g2_tiehi _17157__835 (.L_HI(net835));
 sg13g2_tiehi _17158__836 (.L_HI(net836));
 sg13g2_tiehi _17159__837 (.L_HI(net837));
 sg13g2_tiehi _17160__838 (.L_HI(net838));
 sg13g2_tiehi _17161__839 (.L_HI(net839));
 sg13g2_tiehi _17162__840 (.L_HI(net840));
 sg13g2_tiehi _17163__841 (.L_HI(net841));
 sg13g2_tiehi _17164__842 (.L_HI(net842));
 sg13g2_tiehi _17165__843 (.L_HI(net843));
 sg13g2_tiehi _17166__844 (.L_HI(net844));
 sg13g2_tiehi _17167__845 (.L_HI(net845));
 sg13g2_tiehi _17168__846 (.L_HI(net846));
 sg13g2_tiehi _17169__847 (.L_HI(net847));
 sg13g2_tiehi _17170__848 (.L_HI(net848));
 sg13g2_tiehi _17171__849 (.L_HI(net849));
 sg13g2_tiehi _17172__850 (.L_HI(net850));
 sg13g2_tiehi _17173__851 (.L_HI(net851));
 sg13g2_tiehi _17174__852 (.L_HI(net852));
 sg13g2_tiehi _17175__853 (.L_HI(net853));
 sg13g2_tiehi _17176__854 (.L_HI(net854));
 sg13g2_tiehi _17177__855 (.L_HI(net855));
 sg13g2_tiehi _17889__856 (.L_HI(net856));
 sg13g2_tiehi _17494__857 (.L_HI(net857));
 sg13g2_tiehi _18003__858 (.L_HI(net858));
 sg13g2_tiehi _17493__859 (.L_HI(net859));
 sg13g2_tiehi _17888__860 (.L_HI(net860));
 sg13g2_tiehi _17492__861 (.L_HI(net861));
 sg13g2_tiehi _18060__862 (.L_HI(net862));
 sg13g2_tiehi _17491__863 (.L_HI(net863));
 sg13g2_tiehi _17887__864 (.L_HI(net864));
 sg13g2_tiehi _17490__865 (.L_HI(net865));
 sg13g2_tiehi _18002__866 (.L_HI(net866));
 sg13g2_tiehi _17489__867 (.L_HI(net867));
 sg13g2_tiehi _17886__868 (.L_HI(net868));
 sg13g2_tiehi _17488__869 (.L_HI(net869));
 sg13g2_tiehi _18136__870 (.L_HI(net870));
 sg13g2_tiehi _17487__871 (.L_HI(net871));
 sg13g2_tiehi _17885__872 (.L_HI(net872));
 sg13g2_tiehi _17486__873 (.L_HI(net873));
 sg13g2_tiehi _18001__874 (.L_HI(net874));
 sg13g2_tiehi _17178__875 (.L_HI(net875));
 sg13g2_tiehi _17485__876 (.L_HI(net876));
 sg13g2_tiehi _17884__877 (.L_HI(net877));
 sg13g2_tiehi _17484__878 (.L_HI(net878));
 sg13g2_tiehi _18059__879 (.L_HI(net879));
 sg13g2_tiehi _17483__880 (.L_HI(net880));
 sg13g2_tiehi _17883__881 (.L_HI(net881));
 sg13g2_tiehi _17482__882 (.L_HI(net882));
 sg13g2_tiehi _18000__883 (.L_HI(net883));
 sg13g2_tiehi _17481__884 (.L_HI(net884));
 sg13g2_tiehi _17882__885 (.L_HI(net885));
 sg13g2_tiehi _17480__886 (.L_HI(net886));
 sg13g2_tiehi _18088__887 (.L_HI(net887));
 sg13g2_tiehi _17479__888 (.L_HI(net888));
 sg13g2_tiehi _17881__889 (.L_HI(net889));
 sg13g2_tiehi _17478__890 (.L_HI(net890));
 sg13g2_tiehi _17999__891 (.L_HI(net891));
 sg13g2_tiehi _17477__892 (.L_HI(net892));
 sg13g2_tiehi _17880__893 (.L_HI(net893));
 sg13g2_tiehi _17476__894 (.L_HI(net894));
 sg13g2_tiehi _18058__895 (.L_HI(net895));
 sg13g2_tiehi _17475__896 (.L_HI(net896));
 sg13g2_tiehi _17879__897 (.L_HI(net897));
 sg13g2_tiehi _17474__898 (.L_HI(net898));
 sg13g2_tiehi _17998__899 (.L_HI(net899));
 sg13g2_tiehi _17473__900 (.L_HI(net900));
 sg13g2_tiehi _17878__901 (.L_HI(net901));
 sg13g2_tiehi _17472__902 (.L_HI(net902));
 sg13g2_tiehi _18148__903 (.L_HI(net903));
 sg13g2_tiehi _17471__904 (.L_HI(net904));
 sg13g2_tiehi _17877__905 (.L_HI(net905));
 sg13g2_tiehi _17470__906 (.L_HI(net906));
 sg13g2_tiehi _17997__907 (.L_HI(net907));
 sg13g2_tiehi _17469__908 (.L_HI(net908));
 sg13g2_tiehi _17876__909 (.L_HI(net909));
 sg13g2_tiehi _17468__910 (.L_HI(net910));
 sg13g2_tiehi _18057__911 (.L_HI(net911));
 sg13g2_tiehi _17467__912 (.L_HI(net912));
 sg13g2_tiehi _17875__913 (.L_HI(net913));
 sg13g2_tiehi _17198__914 (.L_HI(net914));
 sg13g2_tiehi _17237__915 (.L_HI(net915));
 sg13g2_tiehi _17238__916 (.L_HI(net916));
 sg13g2_tiehi _17239__917 (.L_HI(net917));
 sg13g2_tiehi _17240__918 (.L_HI(net918));
 sg13g2_tiehi _17466__919 (.L_HI(net919));
 sg13g2_tiehi _17996__920 (.L_HI(net920));
 sg13g2_tiehi _17465__921 (.L_HI(net921));
 sg13g2_tiehi _17874__922 (.L_HI(net922));
 sg13g2_tiehi _17464__923 (.L_HI(net923));
 sg13g2_tiehi _18087__924 (.L_HI(net924));
 sg13g2_tiehi _17463__925 (.L_HI(net925));
 sg13g2_tiehi _17873__926 (.L_HI(net926));
 sg13g2_tiehi _17462__927 (.L_HI(net927));
 sg13g2_tiehi _17995__928 (.L_HI(net928));
 sg13g2_tiehi _17461__929 (.L_HI(net929));
 sg13g2_tiehi _17872__930 (.L_HI(net930));
 sg13g2_tiehi _17460__931 (.L_HI(net931));
 sg13g2_tiehi _18056__932 (.L_HI(net932));
 sg13g2_tiehi _17459__933 (.L_HI(net933));
 sg13g2_tiehi _17871__934 (.L_HI(net934));
 sg13g2_tiehi _17458__935 (.L_HI(net935));
 sg13g2_tiehi _17994__936 (.L_HI(net936));
 sg13g2_tiehi _17457__937 (.L_HI(net937));
 sg13g2_tiehi _17870__938 (.L_HI(net938));
 sg13g2_tiehi _17456__939 (.L_HI(net939));
 sg13g2_tiehi _18135__940 (.L_HI(net940));
 sg13g2_tiehi _17455__941 (.L_HI(net941));
 sg13g2_tiehi _17869__942 (.L_HI(net942));
 sg13g2_tiehi _17454__943 (.L_HI(net943));
 sg13g2_tiehi _17993__944 (.L_HI(net944));
 sg13g2_tiehi _17453__945 (.L_HI(net945));
 sg13g2_tiehi _17868__946 (.L_HI(net946));
 sg13g2_tiehi _17452__947 (.L_HI(net947));
 sg13g2_tiehi _18055__948 (.L_HI(net948));
 sg13g2_tiehi _17451__949 (.L_HI(net949));
 sg13g2_tiehi _17867__950 (.L_HI(net950));
 sg13g2_tiehi _17450__951 (.L_HI(net951));
 sg13g2_tiehi _17992__952 (.L_HI(net952));
 sg13g2_tiehi _17449__953 (.L_HI(net953));
 sg13g2_tiehi _17866__954 (.L_HI(net954));
 sg13g2_tiehi _17448__955 (.L_HI(net955));
 sg13g2_tiehi _18086__956 (.L_HI(net956));
 sg13g2_tiehi _17447__957 (.L_HI(net957));
 sg13g2_tiehi _17865__958 (.L_HI(net958));
 sg13g2_tiehi _17446__959 (.L_HI(net959));
 sg13g2_tiehi _17991__960 (.L_HI(net960));
 sg13g2_tiehi _17445__961 (.L_HI(net961));
 sg13g2_tiehi _17864__962 (.L_HI(net962));
 sg13g2_tiehi _17444__963 (.L_HI(net963));
 sg13g2_tiehi _18054__964 (.L_HI(net964));
 sg13g2_tiehi _17443__965 (.L_HI(net965));
 sg13g2_tiehi _17863__966 (.L_HI(net966));
 sg13g2_tiehi _17442__967 (.L_HI(net967));
 sg13g2_tiehi _17990__968 (.L_HI(net968));
 sg13g2_tiehi _17441__969 (.L_HI(net969));
 sg13g2_tiehi _17862__970 (.L_HI(net970));
 sg13g2_tiehi _17440__971 (.L_HI(net971));
 sg13g2_tiehi _18143__972 (.L_HI(net972));
 sg13g2_tiehi _17439__973 (.L_HI(net973));
 sg13g2_tiehi _17861__974 (.L_HI(net974));
 sg13g2_tiehi _17438__975 (.L_HI(net975));
 sg13g2_tiehi _17989__976 (.L_HI(net976));
 sg13g2_tiehi _17437__977 (.L_HI(net977));
 sg13g2_tiehi _17860__978 (.L_HI(net978));
 sg13g2_tiehi _17436__979 (.L_HI(net979));
 sg13g2_tiehi _18053__980 (.L_HI(net980));
 sg13g2_tiehi _17435__981 (.L_HI(net981));
 sg13g2_tiehi _17859__982 (.L_HI(net982));
 sg13g2_tiehi _17434__983 (.L_HI(net983));
 sg13g2_tiehi _17988__984 (.L_HI(net984));
 sg13g2_tiehi _17433__985 (.L_HI(net985));
 sg13g2_tiehi _17858__986 (.L_HI(net986));
 sg13g2_tiehi _17432__987 (.L_HI(net987));
 sg13g2_tiehi _18085__988 (.L_HI(net988));
 sg13g2_tiehi _17431__989 (.L_HI(net989));
 sg13g2_tiehi _17857__990 (.L_HI(net990));
 sg13g2_tiehi _17430__991 (.L_HI(net991));
 sg13g2_tiehi _17987__992 (.L_HI(net992));
 sg13g2_tiehi _17429__993 (.L_HI(net993));
 sg13g2_tiehi _17856__994 (.L_HI(net994));
 sg13g2_tiehi _17428__995 (.L_HI(net995));
 sg13g2_tiehi _18052__996 (.L_HI(net996));
 sg13g2_tiehi _17427__997 (.L_HI(net997));
 sg13g2_tiehi _17855__998 (.L_HI(net998));
 sg13g2_tiehi _17426__999 (.L_HI(net999));
 sg13g2_tiehi _17986__1000 (.L_HI(net1000));
 sg13g2_tiehi _17425__1001 (.L_HI(net1001));
 sg13g2_tiehi _17854__1002 (.L_HI(net1002));
 sg13g2_tiehi _17424__1003 (.L_HI(net1003));
 sg13g2_tiehi _18134__1004 (.L_HI(net1004));
 sg13g2_tiehi _17423__1005 (.L_HI(net1005));
 sg13g2_tiehi _17853__1006 (.L_HI(net1006));
 sg13g2_tiehi _17422__1007 (.L_HI(net1007));
 sg13g2_tiehi _17985__1008 (.L_HI(net1008));
 sg13g2_tiehi _17421__1009 (.L_HI(net1009));
 sg13g2_tiehi _17852__1010 (.L_HI(net1010));
 sg13g2_tiehi _17420__1011 (.L_HI(net1011));
 sg13g2_tiehi _18051__1012 (.L_HI(net1012));
 sg13g2_tiehi _17419__1013 (.L_HI(net1013));
 sg13g2_tiehi _17851__1014 (.L_HI(net1014));
 sg13g2_tiehi _17418__1015 (.L_HI(net1015));
 sg13g2_tiehi _17984__1016 (.L_HI(net1016));
 sg13g2_tiehi _17417__1017 (.L_HI(net1017));
 sg13g2_tiehi _17850__1018 (.L_HI(net1018));
 sg13g2_tiehi _17416__1019 (.L_HI(net1019));
 sg13g2_tiehi _18084__1020 (.L_HI(net1020));
 sg13g2_tiehi _17415__1021 (.L_HI(net1021));
 sg13g2_tiehi _17849__1022 (.L_HI(net1022));
 sg13g2_tiehi _17414__1023 (.L_HI(net1023));
 sg13g2_tiehi _17983__1024 (.L_HI(net1024));
 sg13g2_tiehi _17413__1025 (.L_HI(net1025));
 sg13g2_tiehi _17848__1026 (.L_HI(net1026));
 sg13g2_tiehi _17412__1027 (.L_HI(net1027));
 sg13g2_tiehi _17847__1028 (.L_HI(net1028));
 sg13g2_tiehi _17411__1029 (.L_HI(net1029));
 sg13g2_tiehi _18050__1030 (.L_HI(net1030));
 sg13g2_tiehi _17410__1031 (.L_HI(net1031));
 sg13g2_tiehi _17846__1032 (.L_HI(net1032));
 sg13g2_tiehi _17409__1033 (.L_HI(net1033));
 sg13g2_tiehi _17845__1034 (.L_HI(net1034));
 sg13g2_tiehi _17408__1035 (.L_HI(net1035));
 sg13g2_tiehi _17982__1036 (.L_HI(net1036));
 sg13g2_tiehi _17407__1037 (.L_HI(net1037));
 sg13g2_tiehi _17844__1038 (.L_HI(net1038));
 sg13g2_tiehi _17406__1039 (.L_HI(net1039));
 sg13g2_tiehi _18146__1040 (.L_HI(net1040));
 sg13g2_tiehi _17405__1041 (.L_HI(net1041));
 sg13g2_tiehi _17843__1042 (.L_HI(net1042));
 sg13g2_tiehi _17404__1043 (.L_HI(net1043));
 sg13g2_tiehi _17981__1044 (.L_HI(net1044));
 sg13g2_tiehi _17403__1045 (.L_HI(net1045));
 sg13g2_tiehi _17842__1046 (.L_HI(net1046));
 sg13g2_tiehi _17402__1047 (.L_HI(net1047));
 sg13g2_tiehi _18049__1048 (.L_HI(net1048));
 sg13g2_tiehi _17401__1049 (.L_HI(net1049));
 sg13g2_tiehi _17841__1050 (.L_HI(net1050));
 sg13g2_tiehi _17400__1051 (.L_HI(net1051));
 sg13g2_tiehi _17840__1052 (.L_HI(net1052));
 sg13g2_tiehi _17399__1053 (.L_HI(net1053));
 sg13g2_tiehi _17980__1054 (.L_HI(net1054));
 sg13g2_tiehi _17398__1055 (.L_HI(net1055));
 sg13g2_tiehi _17839__1056 (.L_HI(net1056));
 sg13g2_tiehi _17397__1057 (.L_HI(net1057));
 sg13g2_tiehi _18083__1058 (.L_HI(net1058));
 sg13g2_tiehi _17396__1059 (.L_HI(net1059));
 sg13g2_tiehi _17838__1060 (.L_HI(net1060));
 sg13g2_tiehi _17395__1061 (.L_HI(net1061));
 sg13g2_tiehi _17979__1062 (.L_HI(net1062));
 sg13g2_tiehi _17394__1063 (.L_HI(net1063));
 sg13g2_tiehi _17837__1064 (.L_HI(net1064));
 sg13g2_tiehi _17393__1065 (.L_HI(net1065));
 sg13g2_tiehi _18048__1066 (.L_HI(net1066));
 sg13g2_tiehi _17392__1067 (.L_HI(net1067));
 sg13g2_tiehi _17836__1068 (.L_HI(net1068));
 sg13g2_tiehi _17391__1069 (.L_HI(net1069));
 sg13g2_tiehi _17835__1070 (.L_HI(net1070));
 sg13g2_tiehi _17390__1071 (.L_HI(net1071));
 sg13g2_tiehi _17978__1072 (.L_HI(net1072));
 sg13g2_tiehi _17389__1073 (.L_HI(net1073));
 sg13g2_tiehi _17834__1074 (.L_HI(net1074));
 sg13g2_tiehi _17388__1075 (.L_HI(net1075));
 sg13g2_tiehi _18133__1076 (.L_HI(net1076));
 sg13g2_tiehi _17387__1077 (.L_HI(net1077));
 sg13g2_tiehi _17833__1078 (.L_HI(net1078));
 sg13g2_tiehi _17386__1079 (.L_HI(net1079));
 sg13g2_tiehi _17832__1080 (.L_HI(net1080));
 sg13g2_tiehi _17385__1081 (.L_HI(net1081));
 sg13g2_tiehi _17977__1082 (.L_HI(net1082));
 sg13g2_tiehi _17384__1083 (.L_HI(net1083));
 sg13g2_tiehi _17831__1084 (.L_HI(net1084));
 sg13g2_tiehi _17383__1085 (.L_HI(net1085));
 sg13g2_tiehi _18047__1086 (.L_HI(net1086));
 sg13g2_tiehi _17382__1087 (.L_HI(net1087));
 sg13g2_tiehi _17830__1088 (.L_HI(net1088));
 sg13g2_tiehi _17381__1089 (.L_HI(net1089));
 sg13g2_tiehi _17976__1090 (.L_HI(net1090));
 sg13g2_tiehi _17380__1091 (.L_HI(net1091));
 sg13g2_tiehi _17829__1092 (.L_HI(net1092));
 sg13g2_tiehi _17379__1093 (.L_HI(net1093));
 sg13g2_tiehi _18082__1094 (.L_HI(net1094));
 sg13g2_tiehi _17378__1095 (.L_HI(net1095));
 sg13g2_tiehi _17828__1096 (.L_HI(net1096));
 sg13g2_tiehi _17377__1097 (.L_HI(net1097));
 sg13g2_tiehi _17827__1098 (.L_HI(net1098));
 sg13g2_tiehi _17376__1099 (.L_HI(net1099));
 sg13g2_tiehi _17826__1100 (.L_HI(net1100));
 sg13g2_tiehi _17375__1101 (.L_HI(net1101));
 sg13g2_tiehi _17975__1102 (.L_HI(net1102));
 sg13g2_tiehi _17374__1103 (.L_HI(net1103));
 sg13g2_tiehi _17825__1104 (.L_HI(net1104));
 sg13g2_tiehi _17373__1105 (.L_HI(net1105));
 sg13g2_tiehi _17824__1106 (.L_HI(net1106));
 sg13g2_tiehi _17372__1107 (.L_HI(net1107));
 sg13g2_tiehi _17823__1108 (.L_HI(net1108));
 sg13g2_tiehi _17371__1109 (.L_HI(net1109));
 sg13g2_tiehi _17822__1110 (.L_HI(net1110));
 sg13g2_tiehi _17370__1111 (.L_HI(net1111));
 sg13g2_tiehi _17821__1112 (.L_HI(net1112));
 sg13g2_tiehi _17369__1113 (.L_HI(net1113));
 sg13g2_tiehi _17820__1114 (.L_HI(net1114));
 sg13g2_tiehi _17368__1115 (.L_HI(net1115));
 sg13g2_tiehi _17819__1116 (.L_HI(net1116));
 sg13g2_tiehi _17367__1117 (.L_HI(net1117));
 sg13g2_tiehi _17818__1118 (.L_HI(net1118));
 sg13g2_tiehi _17366__1119 (.L_HI(net1119));
 sg13g2_tiehi _17817__1120 (.L_HI(net1120));
 sg13g2_tiehi _17365__1121 (.L_HI(net1121));
 sg13g2_tiehi _17816__1122 (.L_HI(net1122));
 sg13g2_tiehi _17364__1123 (.L_HI(net1123));
 sg13g2_tiehi _17815__1124 (.L_HI(net1124));
 sg13g2_tiehi _17363__1125 (.L_HI(net1125));
 sg13g2_tiehi _17814__1126 (.L_HI(net1126));
 sg13g2_tiehi _17362__1127 (.L_HI(net1127));
 sg13g2_tiehi _17813__1128 (.L_HI(net1128));
 sg13g2_tiehi _17361__1129 (.L_HI(net1129));
 sg13g2_tiehi _17812__1130 (.L_HI(net1130));
 sg13g2_tiehi _17360__1131 (.L_HI(net1131));
 sg13g2_tiehi _17811__1132 (.L_HI(net1132));
 sg13g2_tiehi _17359__1133 (.L_HI(net1133));
 sg13g2_tiehi _17810__1134 (.L_HI(net1134));
 sg13g2_tiehi _17358__1135 (.L_HI(net1135));
 sg13g2_tiehi _17809__1136 (.L_HI(net1136));
 sg13g2_tiehi _17357__1137 (.L_HI(net1137));
 sg13g2_tiehi _17808__1138 (.L_HI(net1138));
 sg13g2_tiehi _17356__1139 (.L_HI(net1139));
 sg13g2_tiehi _18046__1140 (.L_HI(net1140));
 sg13g2_tiehi _17355__1141 (.L_HI(net1141));
 sg13g2_tiehi _17807__1142 (.L_HI(net1142));
 sg13g2_tiehi _17354__1143 (.L_HI(net1143));
 sg13g2_tiehi _17974__1144 (.L_HI(net1144));
 sg13g2_tiehi _17353__1145 (.L_HI(net1145));
 sg13g2_tiehi _17806__1146 (.L_HI(net1146));
 sg13g2_tiehi _17352__1147 (.L_HI(net1147));
 sg13g2_tiehi _18142__1148 (.L_HI(net1148));
 sg13g2_tiehi _17351__1149 (.L_HI(net1149));
 sg13g2_tiehi _17805__1150 (.L_HI(net1150));
 sg13g2_tiehi _17350__1151 (.L_HI(net1151));
 sg13g2_tiehi _17973__1152 (.L_HI(net1152));
 sg13g2_tiehi _17349__1153 (.L_HI(net1153));
 sg13g2_tiehi _17804__1154 (.L_HI(net1154));
 sg13g2_tiehi _17348__1155 (.L_HI(net1155));
 sg13g2_tiehi _18045__1156 (.L_HI(net1156));
 sg13g2_tiehi _17347__1157 (.L_HI(net1157));
 sg13g2_tiehi _17803__1158 (.L_HI(net1158));
 sg13g2_tiehi _17346__1159 (.L_HI(net1159));
 sg13g2_tiehi _17972__1160 (.L_HI(net1160));
 sg13g2_tiehi _17345__1161 (.L_HI(net1161));
 sg13g2_tiehi _17802__1162 (.L_HI(net1162));
 sg13g2_tiehi _17344__1163 (.L_HI(net1163));
 sg13g2_tiehi _18081__1164 (.L_HI(net1164));
 sg13g2_tiehi _17343__1165 (.L_HI(net1165));
 sg13g2_tiehi _17801__1166 (.L_HI(net1166));
 sg13g2_tiehi _17342__1167 (.L_HI(net1167));
 sg13g2_tiehi _17971__1168 (.L_HI(net1168));
 sg13g2_tiehi _17341__1169 (.L_HI(net1169));
 sg13g2_tiehi _17800__1170 (.L_HI(net1170));
 sg13g2_tiehi _17340__1171 (.L_HI(net1171));
 sg13g2_tiehi _18044__1172 (.L_HI(net1172));
 sg13g2_tiehi _17339__1173 (.L_HI(net1173));
 sg13g2_tiehi _17799__1174 (.L_HI(net1174));
 sg13g2_tiehi _17338__1175 (.L_HI(net1175));
 sg13g2_tiehi _17970__1176 (.L_HI(net1176));
 sg13g2_tiehi _17337__1177 (.L_HI(net1177));
 sg13g2_tiehi _17798__1178 (.L_HI(net1178));
 sg13g2_tiehi _17336__1179 (.L_HI(net1179));
 sg13g2_tiehi _18132__1180 (.L_HI(net1180));
 sg13g2_tiehi _17335__1181 (.L_HI(net1181));
 sg13g2_tiehi _17797__1182 (.L_HI(net1182));
 sg13g2_tiehi _17334__1183 (.L_HI(net1183));
 sg13g2_tiehi _17969__1184 (.L_HI(net1184));
 sg13g2_tiehi _17333__1185 (.L_HI(net1185));
 sg13g2_tiehi _17332__1186 (.L_HI(net1186));
 sg13g2_tiehi _17796__1187 (.L_HI(net1187));
 sg13g2_tiehi _17331__1188 (.L_HI(net1188));
 sg13g2_tiehi _18043__1189 (.L_HI(net1189));
 sg13g2_tiehi _17330__1190 (.L_HI(net1190));
 sg13g2_tiehi _17795__1191 (.L_HI(net1191));
 sg13g2_tiehi _17329__1192 (.L_HI(net1192));
 sg13g2_tiehi _17968__1193 (.L_HI(net1193));
 sg13g2_tiehi _17328__1194 (.L_HI(net1194));
 sg13g2_tiehi _17794__1195 (.L_HI(net1195));
 sg13g2_tiehi _17327__1196 (.L_HI(net1196));
 sg13g2_tiehi _18080__1197 (.L_HI(net1197));
 sg13g2_tiehi _17326__1198 (.L_HI(net1198));
 sg13g2_tiehi _17793__1199 (.L_HI(net1199));
 sg13g2_tiehi _17325__1200 (.L_HI(net1200));
 sg13g2_tiehi _17967__1201 (.L_HI(net1201));
 sg13g2_tiehi _17324__1202 (.L_HI(net1202));
 sg13g2_tiehi _17792__1203 (.L_HI(net1203));
 sg13g2_tiehi _17323__1204 (.L_HI(net1204));
 sg13g2_tiehi _18042__1205 (.L_HI(net1205));
 sg13g2_tiehi _17322__1206 (.L_HI(net1206));
 sg13g2_tiehi _17791__1207 (.L_HI(net1207));
 sg13g2_tiehi _17321__1208 (.L_HI(net1208));
 sg13g2_tiehi _17966__1209 (.L_HI(net1209));
 sg13g2_tiehi _17320__1210 (.L_HI(net1210));
 sg13g2_tiehi _17790__1211 (.L_HI(net1211));
 sg13g2_tiehi _17319__1212 (.L_HI(net1212));
 sg13g2_tiehi _18141__1213 (.L_HI(net1213));
 sg13g2_tiehi _17318__1214 (.L_HI(net1214));
 sg13g2_tiehi _17789__1215 (.L_HI(net1215));
 sg13g2_tiehi _17317__1216 (.L_HI(net1216));
 sg13g2_tiehi _17965__1217 (.L_HI(net1217));
 sg13g2_tiehi _17316__1218 (.L_HI(net1218));
 sg13g2_tiehi _17788__1219 (.L_HI(net1219));
 sg13g2_tiehi _17315__1220 (.L_HI(net1220));
 sg13g2_tiehi _18041__1221 (.L_HI(net1221));
 sg13g2_tiehi _17314__1222 (.L_HI(net1222));
 sg13g2_tiehi _17787__1223 (.L_HI(net1223));
 sg13g2_tiehi _17313__1224 (.L_HI(net1224));
 sg13g2_tiehi _17964__1225 (.L_HI(net1225));
 sg13g2_tiehi _17312__1226 (.L_HI(net1226));
 sg13g2_tiehi _17786__1227 (.L_HI(net1227));
 sg13g2_tiehi _17241__1228 (.L_HI(net1228));
 sg13g2_tiehi _17551__1229 (.L_HI(net1229));
 sg13g2_tiehi _17552__1230 (.L_HI(net1230));
 sg13g2_tiehi _17553__1231 (.L_HI(net1231));
 sg13g2_tiehi _17554__1232 (.L_HI(net1232));
 sg13g2_tiehi _17555__1233 (.L_HI(net1233));
 sg13g2_tiehi _17556__1234 (.L_HI(net1234));
 sg13g2_tiehi _17557__1235 (.L_HI(net1235));
 sg13g2_tiehi _17558__1236 (.L_HI(net1236));
 sg13g2_tiehi _17559__1237 (.L_HI(net1237));
 sg13g2_tiehi _17560__1238 (.L_HI(net1238));
 sg13g2_tiehi _17561__1239 (.L_HI(net1239));
 sg13g2_tiehi _17311__1240 (.L_HI(net1240));
 sg13g2_tiehi _18079__1241 (.L_HI(net1241));
 sg13g2_tiehi _17310__1242 (.L_HI(net1242));
 sg13g2_tiehi _17785__1243 (.L_HI(net1243));
 sg13g2_tiehi _17309__1244 (.L_HI(net1244));
 sg13g2_tiehi _17963__1245 (.L_HI(net1245));
 sg13g2_tiehi _17308__1246 (.L_HI(net1246));
 sg13g2_tiehi _17784__1247 (.L_HI(net1247));
 sg13g2_tiehi _17307__1248 (.L_HI(net1248));
 sg13g2_tiehi _18040__1249 (.L_HI(net1249));
 sg13g2_tiehi _17306__1250 (.L_HI(net1250));
 sg13g2_tiehi _17783__1251 (.L_HI(net1251));
 sg13g2_tiehi _17305__1252 (.L_HI(net1252));
 sg13g2_tiehi _17962__1253 (.L_HI(net1253));
 sg13g2_tiehi _17304__1254 (.L_HI(net1254));
 sg13g2_tiehi _17782__1255 (.L_HI(net1255));
 sg13g2_tiehi _17303__1256 (.L_HI(net1256));
 sg13g2_tiehi _18131__1257 (.L_HI(net1257));
 sg13g2_tiehi _17302__1258 (.L_HI(net1258));
 sg13g2_tiehi _17781__1259 (.L_HI(net1259));
 sg13g2_tiehi _17301__1260 (.L_HI(net1260));
 sg13g2_tiehi _17961__1261 (.L_HI(net1261));
 sg13g2_tiehi _17300__1262 (.L_HI(net1262));
 sg13g2_tiehi _17780__1263 (.L_HI(net1263));
 sg13g2_tiehi _17299__1264 (.L_HI(net1264));
 sg13g2_tiehi _18039__1265 (.L_HI(net1265));
 sg13g2_tiehi _17298__1266 (.L_HI(net1266));
 sg13g2_tiehi _17779__1267 (.L_HI(net1267));
 sg13g2_tiehi _17297__1268 (.L_HI(net1268));
 sg13g2_tiehi _17960__1269 (.L_HI(net1269));
 sg13g2_tiehi _17296__1270 (.L_HI(net1270));
 sg13g2_tiehi _17778__1271 (.L_HI(net1271));
 sg13g2_tiehi _17295__1272 (.L_HI(net1272));
 sg13g2_tiehi _18078__1273 (.L_HI(net1273));
 sg13g2_tiehi _17294__1274 (.L_HI(net1274));
 sg13g2_tiehi _17777__1275 (.L_HI(net1275));
 sg13g2_tiehi _17293__1276 (.L_HI(net1276));
 sg13g2_tiehi _17959__1277 (.L_HI(net1277));
 sg13g2_tiehi _17292__1278 (.L_HI(net1278));
 sg13g2_tiehi _17776__1279 (.L_HI(net1279));
 sg13g2_tiehi _17291__1280 (.L_HI(net1280));
 sg13g2_tiehi _18038__1281 (.L_HI(net1281));
 sg13g2_tiehi _17290__1282 (.L_HI(net1282));
 sg13g2_tiehi _17775__1283 (.L_HI(net1283));
 sg13g2_tiehi _17289__1284 (.L_HI(net1284));
 sg13g2_tiehi _17958__1285 (.L_HI(net1285));
 sg13g2_tiehi _17288__1286 (.L_HI(net1286));
 sg13g2_tiehi _17774__1287 (.L_HI(net1287));
 sg13g2_tiehi _17287__1288 (.L_HI(net1288));
 sg13g2_tiehi _18130__1289 (.L_HI(net1289));
 sg13g2_tiehi _17286__1290 (.L_HI(net1290));
 sg13g2_tiehi _17773__1291 (.L_HI(net1291));
 sg13g2_tiehi _17285__1292 (.L_HI(net1292));
 sg13g2_tiehi _17957__1293 (.L_HI(net1293));
 sg13g2_tiehi _17284__1294 (.L_HI(net1294));
 sg13g2_tiehi _17772__1295 (.L_HI(net1295));
 sg13g2_tiehi _17283__1296 (.L_HI(net1296));
 sg13g2_tiehi _18037__1297 (.L_HI(net1297));
 sg13g2_tiehi _17282__1298 (.L_HI(net1298));
 sg13g2_tiehi _17771__1299 (.L_HI(net1299));
 sg13g2_tiehi _17281__1300 (.L_HI(net1300));
 sg13g2_tiehi _17956__1301 (.L_HI(net1301));
 sg13g2_tiehi _17280__1302 (.L_HI(net1302));
 sg13g2_tiehi _17279__1303 (.L_HI(net1303));
 sg13g2_tiehi _17770__1304 (.L_HI(net1304));
 sg13g2_tiehi _17278__1305 (.L_HI(net1305));
 sg13g2_tiehi _18077__1306 (.L_HI(net1306));
 sg13g2_tiehi _17277__1307 (.L_HI(net1307));
 sg13g2_tiehi _17769__1308 (.L_HI(net1308));
 sg13g2_tiehi _17276__1309 (.L_HI(net1309));
 sg13g2_tiehi _17955__1310 (.L_HI(net1310));
 sg13g2_tiehi _17275__1311 (.L_HI(net1311));
 sg13g2_tiehi _17768__1312 (.L_HI(net1312));
 sg13g2_tiehi _17274__1313 (.L_HI(net1313));
 sg13g2_tiehi _18036__1314 (.L_HI(net1314));
 sg13g2_tiehi _17273__1315 (.L_HI(net1315));
 sg13g2_tiehi _17767__1316 (.L_HI(net1316));
 sg13g2_tiehi _17272__1317 (.L_HI(net1317));
 sg13g2_tiehi _17954__1318 (.L_HI(net1318));
 sg13g2_tiehi _17271__1319 (.L_HI(net1319));
 sg13g2_tiehi _17766__1320 (.L_HI(net1320));
 sg13g2_tiehi _17270__1321 (.L_HI(net1321));
 sg13g2_tiehi _18129__1322 (.L_HI(net1322));
 sg13g2_tiehi _17269__1323 (.L_HI(net1323));
 sg13g2_tiehi _17765__1324 (.L_HI(net1324));
 sg13g2_tiehi _17268__1325 (.L_HI(net1325));
 sg13g2_tiehi _17953__1326 (.L_HI(net1326));
 sg13g2_tiehi _17267__1327 (.L_HI(net1327));
 sg13g2_tiehi _17764__1328 (.L_HI(net1328));
 sg13g2_tiehi _17266__1329 (.L_HI(net1329));
 sg13g2_tiehi _18035__1330 (.L_HI(net1330));
 sg13g2_tiehi _17265__1331 (.L_HI(net1331));
 sg13g2_tiehi _17763__1332 (.L_HI(net1332));
 sg13g2_tiehi _17264__1333 (.L_HI(net1333));
 sg13g2_tiehi _17952__1334 (.L_HI(net1334));
 sg13g2_tiehi _17263__1335 (.L_HI(net1335));
 sg13g2_tiehi _17562__1336 (.L_HI(net1336));
 sg13g2_tiehi _17762__1337 (.L_HI(net1337));
 sg13g2_tiehi _17262__1338 (.L_HI(net1338));
 sg13g2_tiehi _18076__1339 (.L_HI(net1339));
 sg13g2_tiehi _17261__1340 (.L_HI(net1340));
 sg13g2_tiehi _17761__1341 (.L_HI(net1341));
 sg13g2_tiehi _17260__1342 (.L_HI(net1342));
 sg13g2_tiehi _17951__1343 (.L_HI(net1343));
 sg13g2_tiehi _17259__1344 (.L_HI(net1344));
 sg13g2_tiehi _17760__1345 (.L_HI(net1345));
 sg13g2_tiehi _17258__1346 (.L_HI(net1346));
 sg13g2_tiehi _18034__1347 (.L_HI(net1347));
 sg13g2_tiehi _17257__1348 (.L_HI(net1348));
 sg13g2_tiehi _17759__1349 (.L_HI(net1349));
 sg13g2_tiehi _17256__1350 (.L_HI(net1350));
 sg13g2_tiehi _17950__1351 (.L_HI(net1351));
 sg13g2_tiehi _17255__1352 (.L_HI(net1352));
 sg13g2_tiehi _17758__1353 (.L_HI(net1353));
 sg13g2_tiehi _17254__1354 (.L_HI(net1354));
 sg13g2_tiehi _18140__1355 (.L_HI(net1355));
 sg13g2_tiehi _17253__1356 (.L_HI(net1356));
 sg13g2_tiehi _17757__1357 (.L_HI(net1357));
 sg13g2_tiehi _17252__1358 (.L_HI(net1358));
 sg13g2_tiehi _17949__1359 (.L_HI(net1359));
 sg13g2_tiehi _17251__1360 (.L_HI(net1360));
 sg13g2_tiehi _17756__1361 (.L_HI(net1361));
 sg13g2_tiehi _17250__1362 (.L_HI(net1362));
 sg13g2_tiehi _18033__1363 (.L_HI(net1363));
 sg13g2_tiehi _17249__1364 (.L_HI(net1364));
 sg13g2_tiehi _17755__1365 (.L_HI(net1365));
 sg13g2_tiehi _17248__1366 (.L_HI(net1366));
 sg13g2_tiehi _17948__1367 (.L_HI(net1367));
 sg13g2_tiehi _17247__1368 (.L_HI(net1368));
 sg13g2_tiehi _17754__1369 (.L_HI(net1369));
 sg13g2_tiehi _17246__1370 (.L_HI(net1370));
 sg13g2_tiehi _18075__1371 (.L_HI(net1371));
 sg13g2_tiehi _17245__1372 (.L_HI(net1372));
 sg13g2_tiehi _17753__1373 (.L_HI(net1373));
 sg13g2_tiehi _17659__1374 (.L_HI(net1374));
 sg13g2_tiehi _17244__1375 (.L_HI(net1375));
 sg13g2_tiehi _17947__1376 (.L_HI(net1376));
 sg13g2_tiehi _17243__1377 (.L_HI(net1377));
 sg13g2_tiehi _17752__1378 (.L_HI(net1378));
 sg13g2_tiehi _17242__1379 (.L_HI(net1379));
 sg13g2_tiehi _18032__1380 (.L_HI(net1380));
 sg13g2_tiehi _17236__1381 (.L_HI(net1381));
 sg13g2_tiehi _17751__1382 (.L_HI(net1382));
 sg13g2_tiehi _17235__1383 (.L_HI(net1383));
 sg13g2_tiehi _17946__1384 (.L_HI(net1384));
 sg13g2_tiehi _17234__1385 (.L_HI(net1385));
 sg13g2_tiehi _17750__1386 (.L_HI(net1386));
 sg13g2_tiehi _17233__1387 (.L_HI(net1387));
 sg13g2_tiehi _17232__1388 (.L_HI(net1388));
 sg13g2_tiehi _17231__1389 (.L_HI(net1389));
 sg13g2_tiehi _17230__1390 (.L_HI(net1390));
 sg13g2_tiehi _17229__1391 (.L_HI(net1391));
 sg13g2_tiehi _17228__1392 (.L_HI(net1392));
 sg13g2_tiehi _17227__1393 (.L_HI(net1393));
 sg13g2_tiehi _17226__1394 (.L_HI(net1394));
 sg13g2_tiehi _17225__1395 (.L_HI(net1395));
 sg13g2_tiehi _17224__1396 (.L_HI(net1396));
 sg13g2_tiehi _17223__1397 (.L_HI(net1397));
 sg13g2_tiehi _17222__1398 (.L_HI(net1398));
 sg13g2_tiehi _17221__1399 (.L_HI(net1399));
 sg13g2_tiehi _17220__1400 (.L_HI(net1400));
 sg13g2_tiehi _17219__1401 (.L_HI(net1401));
 sg13g2_tiehi _17218__1402 (.L_HI(net1402));
 sg13g2_tiehi _17217__1403 (.L_HI(net1403));
 sg13g2_tiehi _17216__1404 (.L_HI(net1404));
 sg13g2_tiehi _17215__1405 (.L_HI(net1405));
 sg13g2_tiehi _17214__1406 (.L_HI(net1406));
 sg13g2_tiehi _17213__1407 (.L_HI(net1407));
 sg13g2_tiehi _17212__1408 (.L_HI(net1408));
 sg13g2_tiehi _17211__1409 (.L_HI(net1409));
 sg13g2_tiehi _17210__1410 (.L_HI(net1410));
 sg13g2_tiehi _17209__1411 (.L_HI(net1411));
 sg13g2_tiehi _18096__1412 (.L_HI(net1412));
 sg13g2_tiehi _17208__1413 (.L_HI(net1413));
 sg13g2_tiehi _17749__1414 (.L_HI(net1414));
 sg13g2_tiehi _17207__1415 (.L_HI(net1415));
 sg13g2_tiehi _17945__1416 (.L_HI(net1416));
 sg13g2_tiehi _17206__1417 (.L_HI(net1417));
 sg13g2_tiehi _17748__1418 (.L_HI(net1418));
 sg13g2_tiehi _17205__1419 (.L_HI(net1419));
 sg13g2_tiehi _18031__1420 (.L_HI(net1420));
 sg13g2_tiehi _17204__1421 (.L_HI(net1421));
 sg13g2_tiehi _17747__1422 (.L_HI(net1422));
 sg13g2_tiehi _17203__1423 (.L_HI(net1423));
 sg13g2_tiehi _17944__1424 (.L_HI(net1424));
 sg13g2_tiehi _17202__1425 (.L_HI(net1425));
 sg13g2_tiehi _17201__1426 (.L_HI(net1426));
 sg13g2_tiehi _17200__1427 (.L_HI(net1427));
 sg13g2_tiehi _17746__1428 (.L_HI(net1428));
 sg13g2_tiehi _17199__1429 (.L_HI(net1429));
 sg13g2_tiehi _18074__1430 (.L_HI(net1430));
 sg13g2_tiehi _17197__1431 (.L_HI(net1431));
 sg13g2_tiehi _17745__1432 (.L_HI(net1432));
 sg13g2_tiehi _17196__1433 (.L_HI(net1433));
 sg13g2_tiehi _17195__1434 (.L_HI(net1434));
 sg13g2_tiehi _17943__1435 (.L_HI(net1435));
 sg13g2_tiehi _17194__1436 (.L_HI(net1436));
 sg13g2_tiehi _17744__1437 (.L_HI(net1437));
 sg13g2_tiehi _17193__1438 (.L_HI(net1438));
 sg13g2_tiehi _18030__1439 (.L_HI(net1439));
 sg13g2_tiehi _17192__1440 (.L_HI(net1440));
 sg13g2_tiehi _17743__1441 (.L_HI(net1441));
 sg13g2_tiehi _17191__1442 (.L_HI(net1442));
 sg13g2_tiehi _17942__1443 (.L_HI(net1443));
 sg13g2_tiehi _17190__1444 (.L_HI(net1444));
 sg13g2_tiehi _17742__1445 (.L_HI(net1445));
 sg13g2_tiehi _17189__1446 (.L_HI(net1446));
 sg13g2_tiehi _17188__1447 (.L_HI(net1447));
 sg13g2_tiehi _18128__1448 (.L_HI(net1448));
 sg13g2_tiehi _17187__1449 (.L_HI(net1449));
 sg13g2_tiehi _17741__1450 (.L_HI(net1450));
 sg13g2_tiehi _17186__1451 (.L_HI(net1451));
 sg13g2_tiehi _17941__1452 (.L_HI(net1452));
 sg13g2_tiehi _17185__1453 (.L_HI(net1453));
 sg13g2_tiehi _17740__1454 (.L_HI(net1454));
 sg13g2_tiehi _17184__1455 (.L_HI(net1455));
 sg13g2_tiehi _18029__1456 (.L_HI(net1456));
 sg13g2_tiehi _17183__1457 (.L_HI(net1457));
 sg13g2_tiehi _17739__1458 (.L_HI(net1458));
 sg13g2_tiehi _17182__1459 (.L_HI(net1459));
 sg13g2_tiehi _17940__1460 (.L_HI(net1460));
 sg13g2_tiehi _17181__1461 (.L_HI(net1461));
 sg13g2_tiehi _17738__1462 (.L_HI(net1462));
 sg13g2_tiehi _17180__1463 (.L_HI(net1463));
 sg13g2_tiehi _17179__1464 (.L_HI(net1464));
 sg13g2_tiehi _16764__1465 (.L_HI(net1465));
 sg13g2_tiehi _16763__1466 (.L_HI(net1466));
 sg13g2_tiehi _16762__1467 (.L_HI(net1467));
 sg13g2_tiehi _16761__1468 (.L_HI(net1468));
 sg13g2_tiehi _16760__1469 (.L_HI(net1469));
 sg13g2_tiehi _16759__1470 (.L_HI(net1470));
 sg13g2_tiehi _16730__1471 (.L_HI(net1471));
 sg13g2_tiehi _16729__1472 (.L_HI(net1472));
 sg13g2_tiehi _16728__1473 (.L_HI(net1473));
 sg13g2_tiehi _16727__1474 (.L_HI(net1474));
 sg13g2_tiehi _16726__1475 (.L_HI(net1475));
 sg13g2_tiehi _18073__1476 (.L_HI(net1476));
 sg13g2_tiehi _16697__1477 (.L_HI(net1477));
 sg13g2_tiehi _17737__1478 (.L_HI(net1478));
 sg13g2_tiehi _16696__1479 (.L_HI(net1479));
 sg13g2_tiehi _17939__1480 (.L_HI(net1480));
 sg13g2_tiehi _16695__1481 (.L_HI(net1481));
 sg13g2_tiehi _17736__1482 (.L_HI(net1482));
 sg13g2_tiehi _16694__1483 (.L_HI(net1483));
 sg13g2_tiehi _18028__1484 (.L_HI(net1484));
 sg13g2_tiehi _16693__1485 (.L_HI(net1485));
 sg13g2_tiehi _17735__1486 (.L_HI(net1486));
 sg13g2_tiehi _16692__1487 (.L_HI(net1487));
 sg13g2_tiehi _16691__1488 (.L_HI(net1488));
 sg13g2_tiehi _16690__1489 (.L_HI(net1489));
 sg13g2_tiehi _16689__1490 (.L_HI(net1490));
 sg13g2_tiehi _16688__1491 (.L_HI(net1491));
 sg13g2_tiehi _16687__1492 (.L_HI(net1492));
 sg13g2_tiehi _16686__1493 (.L_HI(net1493));
 sg13g2_tiehi _16685__1494 (.L_HI(net1494));
 sg13g2_tiehi _16684__1495 (.L_HI(net1495));
 sg13g2_tiehi _16683__1496 (.L_HI(net1496));
 sg13g2_tiehi _16682__1497 (.L_HI(net1497));
 sg13g2_tiehi _16681__1498 (.L_HI(net1498));
 sg13g2_tiehi _16680__1499 (.L_HI(net1499));
 sg13g2_tiehi _16679__1500 (.L_HI(net1500));
 sg13g2_tiehi _16678__1501 (.L_HI(net1501));
 sg13g2_tiehi _16677__1502 (.L_HI(net1502));
 sg13g2_tiehi _16676__1503 (.L_HI(net1503));
 sg13g2_tiehi _16675__1504 (.L_HI(net1504));
 sg13g2_tiehi _16674__1505 (.L_HI(net1505));
 sg13g2_tiehi _16673__1506 (.L_HI(net1506));
 sg13g2_tiehi _16672__1507 (.L_HI(net1507));
 sg13g2_tiehi _16671__1508 (.L_HI(net1508));
 sg13g2_tiehi _16670__1509 (.L_HI(net1509));
 sg13g2_tiehi _16669__1510 (.L_HI(net1510));
 sg13g2_tiehi _16668__1511 (.L_HI(net1511));
 sg13g2_tiehi _16667__1512 (.L_HI(net1512));
 sg13g2_tiehi _16666__1513 (.L_HI(net1513));
 sg13g2_tiehi _16665__1514 (.L_HI(net1514));
 sg13g2_tiehi _16664__1515 (.L_HI(net1515));
 sg13g2_tiehi _16663__1516 (.L_HI(net1516));
 sg13g2_tiehi _16662__1517 (.L_HI(net1517));
 sg13g2_tiehi _16661__1518 (.L_HI(net1518));
 sg13g2_tiehi _16660__1519 (.L_HI(net1519));
 sg13g2_tiehi _16659__1520 (.L_HI(net1520));
 sg13g2_tiehi _16658__1521 (.L_HI(net1521));
 sg13g2_tiehi _16657__1522 (.L_HI(net1522));
 sg13g2_tiehi _16656__1523 (.L_HI(net1523));
 sg13g2_tiehi _16655__1524 (.L_HI(net1524));
 sg13g2_tiehi _16654__1525 (.L_HI(net1525));
 sg13g2_tiehi _16653__1526 (.L_HI(net1526));
 sg13g2_tiehi _16652__1527 (.L_HI(net1527));
 sg13g2_tiehi _16651__1528 (.L_HI(net1528));
 sg13g2_tiehi _16650__1529 (.L_HI(net1529));
 sg13g2_tiehi _16649__1530 (.L_HI(net1530));
 sg13g2_tiehi _16648__1531 (.L_HI(net1531));
 sg13g2_tiehi _16647__1532 (.L_HI(net1532));
 sg13g2_tiehi _16646__1533 (.L_HI(net1533));
 sg13g2_tiehi _16645__1534 (.L_HI(net1534));
 sg13g2_tiehi _17938__1535 (.L_HI(net1535));
 sg13g2_tiehi _16644__1536 (.L_HI(net1536));
 sg13g2_tiehi _17734__1537 (.L_HI(net1537));
 sg13g2_tiehi _16643__1538 (.L_HI(net1538));
 sg13g2_tiehi _18095__1539 (.L_HI(net1539));
 sg13g2_tiehi _16642__1540 (.L_HI(net1540));
 sg13g2_tiehi _17733__1541 (.L_HI(net1541));
 sg13g2_tiehi _16641__1542 (.L_HI(net1542));
 sg13g2_tiehi _17937__1543 (.L_HI(net1543));
 sg13g2_tiehi _16640__1544 (.L_HI(net1544));
 sg13g2_tiehi _17732__1545 (.L_HI(net1545));
 sg13g2_tiehi _16639__1546 (.L_HI(net1546));
 sg13g2_tiehi _18027__1547 (.L_HI(net1547));
 sg13g2_tiehi _16638__1548 (.L_HI(net1548));
 sg13g2_tiehi _17731__1549 (.L_HI(net1549));
 sg13g2_tiehi _16637__1550 (.L_HI(net1550));
 sg13g2_tiehi _17936__1551 (.L_HI(net1551));
 sg13g2_tiehi _16636__1552 (.L_HI(net1552));
 sg13g2_tiehi _17730__1553 (.L_HI(net1553));
 sg13g2_tiehi _16635__1554 (.L_HI(net1554));
 sg13g2_tiehi _18072__1555 (.L_HI(net1555));
 sg13g2_tiehi _16634__1556 (.L_HI(net1556));
 sg13g2_tiehi _17729__1557 (.L_HI(net1557));
 sg13g2_tiehi _16633__1558 (.L_HI(net1558));
 sg13g2_tiehi _16632__1559 (.L_HI(net1559));
 sg13g2_tiehi _17935__1560 (.L_HI(net1560));
 sg13g2_tiehi _16631__1561 (.L_HI(net1561));
 sg13g2_tiehi _16630__1562 (.L_HI(net1562));
 sg13g2_tiehi _16629__1563 (.L_HI(net1563));
 sg13g2_tiehi _16628__1564 (.L_HI(net1564));
 sg13g2_tiehi _17728__1565 (.L_HI(net1565));
 sg13g2_tiehi _16627__1566 (.L_HI(net1566));
 sg13g2_tiehi _18026__1567 (.L_HI(net1567));
 sg13g2_tiehi _16626__1568 (.L_HI(net1568));
 sg13g2_tiehi _17727__1569 (.L_HI(net1569));
 sg13g2_tiehi _16625__1570 (.L_HI(net1570));
 sg13g2_tiehi _17934__1571 (.L_HI(net1571));
 sg13g2_tiehi _16624__1572 (.L_HI(net1572));
 sg13g2_tiehi _17726__1573 (.L_HI(net1573));
 sg13g2_tiehi _16623__1574 (.L_HI(net1574));
 sg13g2_tiehi _18139__1575 (.L_HI(net1575));
 sg13g2_tiehi _16622__1576 (.L_HI(net1576));
 sg13g2_tiehi _17725__1577 (.L_HI(net1577));
 sg13g2_tiehi _16621__1578 (.L_HI(net1578));
 sg13g2_tiehi _17933__1579 (.L_HI(net1579));
 sg13g2_tiehi _16619__1580 (.L_HI(net1580));
 sg13g2_tiehi _17724__1581 (.L_HI(net1581));
 sg13g2_tiehi _16618__1582 (.L_HI(net1582));
 sg13g2_tiehi _17723__1583 (.L_HI(net1583));
 sg13g2_tiehi _16617__1584 (.L_HI(net1584));
 sg13g2_tiehi _17722__1585 (.L_HI(net1585));
 sg13g2_tiehi _16616__1586 (.L_HI(net1586));
 sg13g2_tiehi _17721__1587 (.L_HI(net1587));
 sg13g2_tiehi _16615__1588 (.L_HI(net1588));
 sg13g2_tiehi _17720__1589 (.L_HI(net1589));
 sg13g2_tiehi _16614__1590 (.L_HI(net1590));
 sg13g2_tiehi _17719__1591 (.L_HI(net1591));
 sg13g2_tiehi _16613__1592 (.L_HI(net1592));
 sg13g2_tiehi _17718__1593 (.L_HI(net1593));
 sg13g2_tiehi _16612__1594 (.L_HI(net1594));
 sg13g2_tiehi _17717__1595 (.L_HI(net1595));
 sg13g2_tiehi _16611__1596 (.L_HI(net1596));
 sg13g2_tiehi _17716__1597 (.L_HI(net1597));
 sg13g2_tiehi _16610__1598 (.L_HI(net1598));
 sg13g2_tiehi _17715__1599 (.L_HI(net1599));
 sg13g2_tiehi _16609__1600 (.L_HI(net1600));
 sg13g2_tiehi _17714__1601 (.L_HI(net1601));
 sg13g2_tiehi _16608__1602 (.L_HI(net1602));
 sg13g2_tiehi _17713__1603 (.L_HI(net1603));
 sg13g2_tiehi _16607__1604 (.L_HI(net1604));
 sg13g2_tiehi _17712__1605 (.L_HI(net1605));
 sg13g2_tiehi _16606__1606 (.L_HI(net1606));
 sg13g2_tiehi _17711__1607 (.L_HI(net1607));
 sg13g2_tiehi _16605__1608 (.L_HI(net1608));
 sg13g2_tiehi _17710__1609 (.L_HI(net1609));
 sg13g2_tiehi _16604__1610 (.L_HI(net1610));
 sg13g2_tiehi _18025__1611 (.L_HI(net1611));
 sg13g2_tiehi _16603__1612 (.L_HI(net1612));
 sg13g2_tiehi _17709__1613 (.L_HI(net1613));
 sg13g2_tiehi _16602__1614 (.L_HI(net1614));
 sg13g2_tiehi _17708__1615 (.L_HI(net1615));
 sg13g2_tiehi _16601__1616 (.L_HI(net1616));
 sg13g2_tiehi _17707__1617 (.L_HI(net1617));
 sg13g2_tiehi _16600__1618 (.L_HI(net1618));
 sg13g2_tiehi _17706__1619 (.L_HI(net1619));
 sg13g2_tiehi _16599__1620 (.L_HI(net1620));
 sg13g2_tiehi _17705__1621 (.L_HI(net1621));
 sg13g2_tiehi _16598__1622 (.L_HI(net1622));
 sg13g2_tiehi _17704__1623 (.L_HI(net1623));
 sg13g2_tiehi _16597__1624 (.L_HI(net1624));
 sg13g2_tiehi _17703__1625 (.L_HI(net1625));
 sg13g2_tiehi _16596__1626 (.L_HI(net1626));
 sg13g2_tiehi _17702__1627 (.L_HI(net1627));
 sg13g2_tiehi _16595__1628 (.L_HI(net1628));
 sg13g2_tiehi _17701__1629 (.L_HI(net1629));
 sg13g2_tiehi _16594__1630 (.L_HI(net1630));
 sg13g2_tiehi _17700__1631 (.L_HI(net1631));
 sg13g2_tiehi _16593__1632 (.L_HI(net1632));
 sg13g2_tiehi _17699__1633 (.L_HI(net1633));
 sg13g2_tiehi _16592__1634 (.L_HI(net1634));
 sg13g2_tiehi _17932__1635 (.L_HI(net1635));
 sg13g2_tiehi _16591__1636 (.L_HI(net1636));
 sg13g2_tiehi _17698__1637 (.L_HI(net1637));
 sg13g2_tiehi _16590__1638 (.L_HI(net1638));
 sg13g2_tiehi _18071__1639 (.L_HI(net1639));
 sg13g2_tiehi _16589__1640 (.L_HI(net1640));
 sg13g2_tiehi _17696__1641 (.L_HI(net1641));
 sg13g2_tiehi _16588__1642 (.L_HI(net1642));
 sg13g2_tiehi _17931__1643 (.L_HI(net1643));
 sg13g2_tiehi _16587__1644 (.L_HI(net1644));
 sg13g2_tiehi _17695__1645 (.L_HI(net1645));
 sg13g2_tiehi _16586__1646 (.L_HI(net1646));
 sg13g2_tiehi _18024__1647 (.L_HI(net1647));
 sg13g2_tiehi _16585__1648 (.L_HI(net1648));
 sg13g2_tiehi _17694__1649 (.L_HI(net1649));
 sg13g2_tiehi _16584__1650 (.L_HI(net1650));
 sg13g2_tiehi _17930__1651 (.L_HI(net1651));
 sg13g2_tiehi _16583__1652 (.L_HI(net1652));
 sg13g2_tiehi _17693__1653 (.L_HI(net1653));
 sg13g2_tiehi _16582__1654 (.L_HI(net1654));
 sg13g2_tiehi _18094__1655 (.L_HI(net1655));
 sg13g2_tiehi _16581__1656 (.L_HI(net1656));
 sg13g2_tiehi _17692__1657 (.L_HI(net1657));
 sg13g2_tiehi _16580__1658 (.L_HI(net1658));
 sg13g2_tiehi _17929__1659 (.L_HI(net1659));
 sg13g2_tiehi _16579__1660 (.L_HI(net1660));
 sg13g2_tiehi _17691__1661 (.L_HI(net1661));
 sg13g2_tiehi _16578__1662 (.L_HI(net1662));
 sg13g2_tiehi _18023__1663 (.L_HI(net1663));
 sg13g2_tiehi _16577__1664 (.L_HI(net1664));
 sg13g2_tiehi _17690__1665 (.L_HI(net1665));
 sg13g2_tiehi _16576__1666 (.L_HI(net1666));
 sg13g2_tiehi _17928__1667 (.L_HI(net1667));
 sg13g2_tiehi _16575__1668 (.L_HI(net1668));
 sg13g2_tiehi _17689__1669 (.L_HI(net1669));
 sg13g2_tiehi _16574__1670 (.L_HI(net1670));
 sg13g2_tiehi _18070__1671 (.L_HI(net1671));
 sg13g2_tiehi _16573__1672 (.L_HI(net1672));
 sg13g2_tiehi _17688__1673 (.L_HI(net1673));
 sg13g2_tiehi _16572__1674 (.L_HI(net1674));
 sg13g2_tiehi _17927__1675 (.L_HI(net1675));
 sg13g2_tiehi _16571__1676 (.L_HI(net1676));
 sg13g2_tiehi _17687__1677 (.L_HI(net1677));
 sg13g2_tiehi _16570__1678 (.L_HI(net1678));
 sg13g2_tiehi _18022__1679 (.L_HI(net1679));
 sg13g2_tiehi _16569__1680 (.L_HI(net1680));
 sg13g2_tiehi _17686__1681 (.L_HI(net1681));
 sg13g2_tiehi _16568__1682 (.L_HI(net1682));
 sg13g2_tiehi _17926__1683 (.L_HI(net1683));
 sg13g2_tiehi _16567__1684 (.L_HI(net1684));
 sg13g2_tiehi _17685__1685 (.L_HI(net1685));
 sg13g2_tiehi _16566__1686 (.L_HI(net1686));
 sg13g2_tiehi _18145__1687 (.L_HI(net1687));
 sg13g2_tiehi _16565__1688 (.L_HI(net1688));
 sg13g2_tiehi _17684__1689 (.L_HI(net1689));
 sg13g2_tiehi _16564__1690 (.L_HI(net1690));
 sg13g2_tiehi _17925__1691 (.L_HI(net1691));
 sg13g2_tiehi _16563__1692 (.L_HI(net1692));
 sg13g2_tiehi _17683__1693 (.L_HI(net1693));
 sg13g2_tiehi _16562__1694 (.L_HI(net1694));
 sg13g2_tiehi _18021__1695 (.L_HI(net1695));
 sg13g2_tiehi _16561__1696 (.L_HI(net1696));
 sg13g2_tiehi _17682__1697 (.L_HI(net1697));
 sg13g2_tiehi _16560__1698 (.L_HI(net1698));
 sg13g2_tiehi _17924__1699 (.L_HI(net1699));
 sg13g2_tiehi _16559__1700 (.L_HI(net1700));
 sg13g2_tiehi _17681__1701 (.L_HI(net1701));
 sg13g2_tiehi _16558__1702 (.L_HI(net1702));
 sg13g2_tiehi _18069__1703 (.L_HI(net1703));
 sg13g2_tiehi _16557__1704 (.L_HI(net1704));
 sg13g2_tiehi _17680__1705 (.L_HI(net1705));
 sg13g2_tiehi _16556__1706 (.L_HI(net1706));
 sg13g2_tiehi _17923__1707 (.L_HI(net1707));
 sg13g2_tiehi _16555__1708 (.L_HI(net1708));
 sg13g2_tiehi _16554__1709 (.L_HI(net1709));
 sg13g2_tiehi _16553__1710 (.L_HI(net1710));
 sg13g2_tiehi _16552__1711 (.L_HI(net1711));
 sg13g2_tiehi _16551__1712 (.L_HI(net1712));
 sg13g2_tiehi _16550__1713 (.L_HI(net1713));
 sg13g2_tiehi _16549__1714 (.L_HI(net1714));
 sg13g2_tiehi _16548__1715 (.L_HI(net1715));
 sg13g2_tiehi _16547__1716 (.L_HI(net1716));
 sg13g2_tiehi _16546__1717 (.L_HI(net1717));
 sg13g2_tiehi _16545__1718 (.L_HI(net1718));
 sg13g2_tiehi _16544__1719 (.L_HI(net1719));
 sg13g2_tiehi _16543__1720 (.L_HI(net1720));
 sg13g2_tiehi _16542__1721 (.L_HI(net1721));
 sg13g2_tiehi _16541__1722 (.L_HI(net1722));
 sg13g2_tiehi _16540__1723 (.L_HI(net1723));
 sg13g2_tiehi _16539__1724 (.L_HI(net1724));
 sg13g2_tiehi _16538__1725 (.L_HI(net1725));
 sg13g2_tiehi _16537__1726 (.L_HI(net1726));
 sg13g2_tiehi _16536__1727 (.L_HI(net1727));
 sg13g2_tiehi _16535__1728 (.L_HI(net1728));
 sg13g2_tiehi _16534__1729 (.L_HI(net1729));
 sg13g2_tiehi _16533__1730 (.L_HI(net1730));
 sg13g2_tiehi _16532__1731 (.L_HI(net1731));
 sg13g2_tiehi _16531__1732 (.L_HI(net1732));
 sg13g2_tiehi _16530__1733 (.L_HI(net1733));
 sg13g2_tiehi _16529__1734 (.L_HI(net1734));
 sg13g2_tiehi _16528__1735 (.L_HI(net1735));
 sg13g2_tiehi _16527__1736 (.L_HI(net1736));
 sg13g2_tiehi _16526__1737 (.L_HI(net1737));
 sg13g2_tiehi _16525__1738 (.L_HI(net1738));
 sg13g2_tiehi _16524__1739 (.L_HI(net1739));
 sg13g2_tiehi _17679__1740 (.L_HI(net1740));
 sg13g2_tiehi _16523__1741 (.L_HI(net1741));
 sg13g2_tiehi _18020__1742 (.L_HI(net1742));
 sg13g2_tiehi _16522__1743 (.L_HI(net1743));
 sg13g2_tiehi _16521__1744 (.L_HI(net1744));
 sg13g2_tiehi _16520__1745 (.L_HI(net1745));
 sg13g2_tiehi _16519__1746 (.L_HI(net1746));
 sg13g2_tiehi _16518__1747 (.L_HI(net1747));
 sg13g2_tiehi _16517__1748 (.L_HI(net1748));
 sg13g2_tiehi _16516__1749 (.L_HI(net1749));
 sg13g2_tiehi _16515__1750 (.L_HI(net1750));
 sg13g2_tiehi _16514__1751 (.L_HI(net1751));
 sg13g2_tiehi _16513__1752 (.L_HI(net1752));
 sg13g2_tiehi _16512__1753 (.L_HI(net1753));
 sg13g2_tiehi _16511__1754 (.L_HI(net1754));
 sg13g2_tiehi _16510__1755 (.L_HI(net1755));
 sg13g2_tiehi _16509__1756 (.L_HI(net1756));
 sg13g2_tiehi _16508__1757 (.L_HI(net1757));
 sg13g2_tiehi _16507__1758 (.L_HI(net1758));
 sg13g2_tiehi _16506__1759 (.L_HI(net1759));
 sg13g2_tiehi _17678__1760 (.L_HI(net1760));
 sg13g2_tiehi _16505__1761 (.L_HI(net1761));
 sg13g2_tiehi _17922__1762 (.L_HI(net1762));
 sg13g2_tiehi _16504__1763 (.L_HI(net1763));
 sg13g2_tiehi _17677__1764 (.L_HI(net1764));
 sg13g2_tiehi _16503__1765 (.L_HI(net1765));
 sg13g2_tiehi _17676__1766 (.L_HI(net1766));
 sg13g2_tiehi _16502__1767 (.L_HI(net1767));
 sg13g2_tiehi _17675__1768 (.L_HI(net1768));
 sg13g2_tiehi _16501__1769 (.L_HI(net1769));
 sg13g2_tiehi _17674__1770 (.L_HI(net1770));
 sg13g2_tiehi _16500__1771 (.L_HI(net1771));
 sg13g2_tiehi _17673__1772 (.L_HI(net1772));
 sg13g2_tiehi _16499__1773 (.L_HI(net1773));
 sg13g2_tiehi _17697__1774 (.L_HI(net1774));
 sg13g2_tiehi _18097__1775 (.L_HI(net1775));
 sg13g2_tiehi _18098__1776 (.L_HI(net1776));
 sg13g2_tiehi _18099__1777 (.L_HI(net1777));
 sg13g2_tiehi _18100__1778 (.L_HI(net1778));
 sg13g2_tiehi _18101__1779 (.L_HI(net1779));
 sg13g2_tiehi _18102__1780 (.L_HI(net1780));
 sg13g2_tiehi _18103__1781 (.L_HI(net1781));
 sg13g2_tiehi _18104__1782 (.L_HI(net1782));
 sg13g2_tiehi _18105__1783 (.L_HI(net1783));
 sg13g2_tiehi _18106__1784 (.L_HI(net1784));
 sg13g2_tiehi _18107__1785 (.L_HI(net1785));
 sg13g2_tiehi _18108__1786 (.L_HI(net1786));
 sg13g2_tiehi _18109__1787 (.L_HI(net1787));
 sg13g2_tiehi _18110__1788 (.L_HI(net1788));
 sg13g2_tiehi _18111__1789 (.L_HI(net1789));
 sg13g2_tiehi _18112__1790 (.L_HI(net1790));
 sg13g2_tiehi _18113__1791 (.L_HI(net1791));
 sg13g2_tiehi _18114__1792 (.L_HI(net1792));
 sg13g2_tiehi _18115__1793 (.L_HI(net2675));
 sg13g2_tiehi _18116__1794 (.L_HI(net2676));
 sg13g2_tiehi _18117__1795 (.L_HI(net2677));
 sg13g2_tiehi _18118__1796 (.L_HI(net2678));
 sg13g2_tiehi _18119__1797 (.L_HI(net2679));
 sg13g2_tiehi _18120__1798 (.L_HI(net2680));
 sg13g2_tiehi _18121__1799 (.L_HI(net2681));
 sg13g2_tiehi _18122__1800 (.L_HI(net2682));
 sg13g2_tiehi _18123__1801 (.L_HI(net2683));
 sg13g2_tiehi _18124__1802 (.L_HI(net2684));
 sg13g2_tiehi _18125__1803 (.L_HI(net2685));
 sg13g2_tiehi _18126__1804 (.L_HI(net2686));
 sg13g2_tiehi _18127__1805 (.L_HI(net2687));
 sg13g2_tiehi _17672__1806 (.L_HI(net2688));
 sg13g2_tiehi _16498__1807 (.L_HI(net2689));
 sg13g2_tiehi _18093__1808 (.L_HI(net2690));
 sg13g2_tiehi _16497__1809 (.L_HI(net2691));
 sg13g2_tiehi _16496__1810 (.L_HI(net2692));
 sg13g2_tiehi _17671__1811 (.L_HI(net2693));
 sg13g2_tiehi _16495__1812 (.L_HI(net2694));
 sg13g2_tiehi _17670__1813 (.L_HI(net2695));
 sg13g2_tiehi _16494__1814 (.L_HI(net2696));
 sg13g2_tiehi _17921__1815 (.L_HI(net2697));
 sg13g2_tiehi _16493__1816 (.L_HI(net2698));
 sg13g2_tiehi _17669__1817 (.L_HI(net2699));
 sg13g2_tiehi _16492__1818 (.L_HI(net2700));
 sg13g2_tiehi _17668__1819 (.L_HI(net2701));
 sg13g2_tiehi _16491__1820 (.L_HI(net2702));
 sg13g2_tiehi _16490__1821 (.L_HI(net2703));
 sg13g2_tiehi _16489__1822 (.L_HI(net2704));
 sg13g2_tiehi _16488__1823 (.L_HI(net2705));
 sg13g2_tiehi _16487__1824 (.L_HI(net2706));
 sg13g2_tiehi _16486__1825 (.L_HI(net2707));
 sg13g2_tiehi _17667__1826 (.L_HI(net2708));
 sg13g2_tiehi _16485__1827 (.L_HI(net2709));
 sg13g2_tiehi _16484__1828 (.L_HI(net2710));
 sg13g2_tiehi _16483__1829 (.L_HI(net2711));
 sg13g2_tiehi _16482__1830 (.L_HI(net2712));
 sg13g2_tiehi _16481__1831 (.L_HI(net2713));
 sg13g2_tiehi _16480__1832 (.L_HI(net2714));
 sg13g2_tiehi _16479__1833 (.L_HI(net2715));
 sg13g2_tiehi _16478__1834 (.L_HI(net2716));
 sg13g2_tiehi _16477__1835 (.L_HI(net2717));
 sg13g2_tiehi _16476__1836 (.L_HI(net2718));
 sg13g2_tiehi _16475__1837 (.L_HI(net2719));
 sg13g2_tiehi _16474__1838 (.L_HI(net2720));
 sg13g2_inv_1 _09414__1 (.Y(net2721),
    .A(clknet_leaf_65_clk));
 sg13g2_buf_1 _19974_ (.A(net2617),
    .X(uio_oe[0]));
 sg13g2_buf_1 _19975_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _19976_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _19977_ (.A(net2617),
    .X(uio_oe[3]));
 sg13g2_buf_1 _19978_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _19979_ (.A(net2617),
    .X(uio_oe[6]));
 sg13g2_buf_1 _19980_ (.A(net2617),
    .X(uio_oe[7]));
 sg13g2_buf_1 _19981_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .X(uio_out[0]));
 sg13g2_buf_8 _19982_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .X(uio_out[3]));
 sg13g2_buf_1 _19983_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .X(uio_out[6]));
 sg13g2_buf_2 _19984_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .X(uio_out[7]));
 sg13g2_buf_8 fanout1793 (.A(net1794),
    .X(net1793));
 sg13g2_buf_2 fanout1794 (.A(net1795),
    .X(net1794));
 sg13g2_buf_2 fanout1795 (.A(_04784_),
    .X(net1795));
 sg13g2_buf_8 fanout1796 (.A(net1797),
    .X(net1796));
 sg13g2_buf_8 fanout1797 (.A(_04012_),
    .X(net1797));
 sg13g2_buf_8 fanout1798 (.A(_03880_),
    .X(net1798));
 sg13g2_buf_8 fanout1799 (.A(_03880_),
    .X(net1799));
 sg13g2_buf_8 fanout1800 (.A(net1802),
    .X(net1800));
 sg13g2_buf_8 fanout1801 (.A(net1802),
    .X(net1801));
 sg13g2_buf_8 fanout1802 (.A(_06716_),
    .X(net1802));
 sg13g2_buf_8 fanout1803 (.A(net1805),
    .X(net1803));
 sg13g2_buf_8 fanout1804 (.A(net1805),
    .X(net1804));
 sg13g2_buf_8 fanout1805 (.A(_06117_),
    .X(net1805));
 sg13g2_buf_8 fanout1806 (.A(_05974_),
    .X(net1806));
 sg13g2_buf_8 fanout1807 (.A(_05974_),
    .X(net1807));
 sg13g2_buf_8 fanout1808 (.A(net1809),
    .X(net1808));
 sg13g2_buf_8 fanout1809 (.A(_05780_),
    .X(net1809));
 sg13g2_buf_8 fanout1810 (.A(_04826_),
    .X(net1810));
 sg13g2_buf_8 fanout1811 (.A(net1813),
    .X(net1811));
 sg13g2_buf_8 fanout1812 (.A(net1813),
    .X(net1812));
 sg13g2_buf_8 fanout1813 (.A(_04654_),
    .X(net1813));
 sg13g2_buf_8 fanout1814 (.A(_03749_),
    .X(net1814));
 sg13g2_buf_8 fanout1815 (.A(_03749_),
    .X(net1815));
 sg13g2_buf_8 fanout1816 (.A(_03564_),
    .X(net1816));
 sg13g2_buf_8 fanout1817 (.A(_03564_),
    .X(net1817));
 sg13g2_buf_8 fanout1818 (.A(net1819),
    .X(net1818));
 sg13g2_buf_8 fanout1819 (.A(net1822),
    .X(net1819));
 sg13g2_buf_8 fanout1820 (.A(net1821),
    .X(net1820));
 sg13g2_buf_8 fanout1821 (.A(net1822),
    .X(net1821));
 sg13g2_buf_2 fanout1822 (.A(net1823),
    .X(net1822));
 sg13g2_buf_8 fanout1823 (.A(net1830),
    .X(net1823));
 sg13g2_buf_8 fanout1824 (.A(net1828),
    .X(net1824));
 sg13g2_buf_8 fanout1825 (.A(net1827),
    .X(net1825));
 sg13g2_buf_8 fanout1826 (.A(net1827),
    .X(net1826));
 sg13g2_buf_2 fanout1827 (.A(net1828),
    .X(net1827));
 sg13g2_buf_1 fanout1828 (.A(net1830),
    .X(net1828));
 sg13g2_buf_8 fanout1829 (.A(net1830),
    .X(net1829));
 sg13g2_buf_8 fanout1830 (.A(_05508_),
    .X(net1830));
 sg13g2_buf_8 fanout1831 (.A(net1832),
    .X(net1831));
 sg13g2_buf_1 fanout1832 (.A(net1834),
    .X(net1832));
 sg13g2_buf_8 fanout1833 (.A(net1834),
    .X(net1833));
 sg13g2_buf_1 fanout1834 (.A(_04740_),
    .X(net1834));
 sg13g2_buf_8 fanout1835 (.A(_04739_),
    .X(net1835));
 sg13g2_buf_1 fanout1836 (.A(_04739_),
    .X(net1836));
 sg13g2_buf_8 fanout1837 (.A(net1839),
    .X(net1837));
 sg13g2_buf_8 fanout1838 (.A(net1839),
    .X(net1838));
 sg13g2_buf_8 fanout1839 (.A(_06797_),
    .X(net1839));
 sg13g2_buf_8 fanout1840 (.A(net1841),
    .X(net1840));
 sg13g2_buf_8 fanout1841 (.A(_05454_),
    .X(net1841));
 sg13g2_buf_8 fanout1842 (.A(_05453_),
    .X(net1842));
 sg13g2_buf_1 fanout1843 (.A(_05453_),
    .X(net1843));
 sg13g2_buf_8 fanout1844 (.A(net1845),
    .X(net1844));
 sg13g2_buf_8 fanout1845 (.A(net1846),
    .X(net1845));
 sg13g2_buf_8 fanout1846 (.A(net1847),
    .X(net1846));
 sg13g2_buf_8 fanout1847 (.A(_04994_),
    .X(net1847));
 sg13g2_buf_8 fanout1848 (.A(net1851),
    .X(net1848));
 sg13g2_buf_1 fanout1849 (.A(net1851),
    .X(net1849));
 sg13g2_buf_8 fanout1850 (.A(net1851),
    .X(net1850));
 sg13g2_buf_8 fanout1851 (.A(_04993_),
    .X(net1851));
 sg13g2_buf_8 fanout1852 (.A(net1853),
    .X(net1852));
 sg13g2_buf_1 fanout1853 (.A(net1854),
    .X(net1853));
 sg13g2_buf_8 fanout1854 (.A(_04733_),
    .X(net1854));
 sg13g2_buf_8 fanout1855 (.A(net1856),
    .X(net1855));
 sg13g2_buf_1 fanout1856 (.A(_04733_),
    .X(net1856));
 sg13g2_buf_8 fanout1857 (.A(net1861),
    .X(net1857));
 sg13g2_buf_8 fanout1858 (.A(net1861),
    .X(net1858));
 sg13g2_buf_8 fanout1859 (.A(net1861),
    .X(net1859));
 sg13g2_buf_1 fanout1860 (.A(net1861),
    .X(net1860));
 sg13g2_buf_8 fanout1861 (.A(_04732_),
    .X(net1861));
 sg13g2_buf_8 fanout1862 (.A(net1863),
    .X(net1862));
 sg13g2_buf_8 fanout1863 (.A(_07078_),
    .X(net1863));
 sg13g2_buf_8 fanout1864 (.A(_04648_),
    .X(net1864));
 sg13g2_buf_8 fanout1865 (.A(net1866),
    .X(net1865));
 sg13g2_buf_8 fanout1866 (.A(_04648_),
    .X(net1866));
 sg13g2_buf_8 fanout1867 (.A(net1868),
    .X(net1867));
 sg13g2_buf_2 fanout1868 (.A(_04647_),
    .X(net1868));
 sg13g2_buf_8 fanout1869 (.A(net1870),
    .X(net1869));
 sg13g2_buf_8 fanout1870 (.A(_04647_),
    .X(net1870));
 sg13g2_buf_8 fanout1871 (.A(net1872),
    .X(net1871));
 sg13g2_buf_8 fanout1872 (.A(_06126_),
    .X(net1872));
 sg13g2_buf_8 fanout1873 (.A(net1874),
    .X(net1873));
 sg13g2_buf_8 fanout1874 (.A(_04603_),
    .X(net1874));
 sg13g2_buf_8 fanout1875 (.A(_04603_),
    .X(net1875));
 sg13g2_buf_8 fanout1876 (.A(net1877),
    .X(net1876));
 sg13g2_buf_8 fanout1877 (.A(net1878),
    .X(net1877));
 sg13g2_buf_8 fanout1878 (.A(net1879),
    .X(net1878));
 sg13g2_buf_8 fanout1879 (.A(net1884),
    .X(net1879));
 sg13g2_buf_8 fanout1880 (.A(net1884),
    .X(net1880));
 sg13g2_buf_1 fanout1881 (.A(net1884),
    .X(net1881));
 sg13g2_buf_8 fanout1882 (.A(net1883),
    .X(net1882));
 sg13g2_buf_8 fanout1883 (.A(net1884),
    .X(net1883));
 sg13g2_buf_8 fanout1884 (.A(_04574_),
    .X(net1884));
 sg13g2_buf_8 fanout1885 (.A(net1886),
    .X(net1885));
 sg13g2_buf_2 fanout1886 (.A(_04323_),
    .X(net1886));
 sg13g2_buf_8 fanout1887 (.A(net1888),
    .X(net1887));
 sg13g2_buf_8 fanout1888 (.A(_06763_),
    .X(net1888));
 sg13g2_buf_2 fanout1889 (.A(_03147_),
    .X(net1889));
 sg13g2_buf_8 fanout1890 (.A(net1892),
    .X(net1890));
 sg13g2_buf_2 fanout1891 (.A(net1892),
    .X(net1891));
 sg13g2_buf_2 fanout1892 (.A(_07048_),
    .X(net1892));
 sg13g2_buf_8 fanout1893 (.A(net1896),
    .X(net1893));
 sg13g2_buf_8 fanout1894 (.A(net1896),
    .X(net1894));
 sg13g2_buf_1 fanout1895 (.A(net1896),
    .X(net1895));
 sg13g2_buf_8 fanout1896 (.A(_06903_),
    .X(net1896));
 sg13g2_buf_8 fanout1897 (.A(net1898),
    .X(net1897));
 sg13g2_buf_1 fanout1898 (.A(net1899),
    .X(net1898));
 sg13g2_buf_1 fanout1899 (.A(_06840_),
    .X(net1899));
 sg13g2_buf_8 fanout1900 (.A(net1901),
    .X(net1900));
 sg13g2_buf_2 fanout1901 (.A(net1902),
    .X(net1901));
 sg13g2_buf_1 fanout1902 (.A(net1903),
    .X(net1902));
 sg13g2_buf_1 fanout1903 (.A(_07067_),
    .X(net1903));
 sg13g2_buf_8 fanout1904 (.A(_07029_),
    .X(net1904));
 sg13g2_buf_1 fanout1905 (.A(_07029_),
    .X(net1905));
 sg13g2_buf_8 fanout1906 (.A(_03421_),
    .X(net1906));
 sg13g2_buf_8 fanout1907 (.A(_03421_),
    .X(net1907));
 sg13g2_buf_8 fanout1908 (.A(_03417_),
    .X(net1908));
 sg13g2_buf_8 fanout1909 (.A(net1910),
    .X(net1909));
 sg13g2_buf_8 fanout1910 (.A(_02441_),
    .X(net1910));
 sg13g2_buf_8 fanout1911 (.A(_02331_),
    .X(net1911));
 sg13g2_buf_8 fanout1912 (.A(_02331_),
    .X(net1912));
 sg13g2_buf_8 fanout1913 (.A(net1914),
    .X(net1913));
 sg13g2_buf_8 fanout1914 (.A(_02309_),
    .X(net1914));
 sg13g2_buf_8 fanout1915 (.A(_02237_),
    .X(net1915));
 sg13g2_buf_8 fanout1916 (.A(_02237_),
    .X(net1916));
 sg13g2_buf_8 fanout1917 (.A(_02169_),
    .X(net1917));
 sg13g2_buf_8 fanout1918 (.A(_02169_),
    .X(net1918));
 sg13g2_buf_8 fanout1919 (.A(net1920),
    .X(net1919));
 sg13g2_buf_8 fanout1920 (.A(_02108_),
    .X(net1920));
 sg13g2_buf_8 fanout1921 (.A(net1922),
    .X(net1921));
 sg13g2_buf_8 fanout1922 (.A(_01698_),
    .X(net1922));
 sg13g2_buf_8 fanout1923 (.A(_06791_),
    .X(net1923));
 sg13g2_buf_8 fanout1924 (.A(_06599_),
    .X(net1924));
 sg13g2_buf_1 fanout1925 (.A(_06599_),
    .X(net1925));
 sg13g2_buf_8 fanout1926 (.A(net1928),
    .X(net1926));
 sg13g2_buf_8 fanout1927 (.A(net1928),
    .X(net1927));
 sg13g2_buf_8 fanout1928 (.A(net1930),
    .X(net1928));
 sg13g2_buf_1 fanout1929 (.A(net1930),
    .X(net1929));
 sg13g2_buf_8 fanout1930 (.A(net1933),
    .X(net1930));
 sg13g2_buf_8 fanout1931 (.A(net1932),
    .X(net1931));
 sg13g2_buf_8 fanout1932 (.A(net1933),
    .X(net1932));
 sg13g2_buf_8 fanout1933 (.A(_06599_),
    .X(net1933));
 sg13g2_buf_8 fanout1934 (.A(net1937),
    .X(net1934));
 sg13g2_buf_2 fanout1935 (.A(net1937),
    .X(net1935));
 sg13g2_buf_8 fanout1936 (.A(net1937),
    .X(net1936));
 sg13g2_buf_8 fanout1937 (.A(_06395_),
    .X(net1937));
 sg13g2_buf_8 fanout1938 (.A(net1943),
    .X(net1938));
 sg13g2_buf_8 fanout1939 (.A(net1942),
    .X(net1939));
 sg13g2_buf_2 fanout1940 (.A(net1942),
    .X(net1940));
 sg13g2_buf_8 fanout1941 (.A(net1942),
    .X(net1941));
 sg13g2_buf_2 fanout1942 (.A(net1943),
    .X(net1942));
 sg13g2_buf_1 fanout1943 (.A(net1944),
    .X(net1943));
 sg13g2_buf_8 fanout1944 (.A(_06395_),
    .X(net1944));
 sg13g2_buf_8 fanout1945 (.A(net1946),
    .X(net1945));
 sg13g2_buf_1 fanout1946 (.A(net1949),
    .X(net1946));
 sg13g2_buf_8 fanout1947 (.A(net1949),
    .X(net1947));
 sg13g2_buf_1 fanout1948 (.A(net1949),
    .X(net1948));
 sg13g2_buf_8 fanout1949 (.A(_06282_),
    .X(net1949));
 sg13g2_buf_8 fanout1950 (.A(net1951),
    .X(net1950));
 sg13g2_buf_8 fanout1951 (.A(net1952),
    .X(net1951));
 sg13g2_buf_8 fanout1952 (.A(_06226_),
    .X(net1952));
 sg13g2_buf_8 fanout1953 (.A(net1954),
    .X(net1953));
 sg13g2_buf_1 fanout1954 (.A(net1955),
    .X(net1954));
 sg13g2_buf_1 fanout1955 (.A(_06226_),
    .X(net1955));
 sg13g2_buf_8 fanout1956 (.A(_05852_),
    .X(net1956));
 sg13g2_buf_1 fanout1957 (.A(_05852_),
    .X(net1957));
 sg13g2_buf_8 fanout1958 (.A(_05546_),
    .X(net1958));
 sg13g2_buf_8 fanout1959 (.A(_02461_),
    .X(net1959));
 sg13g2_buf_8 fanout1960 (.A(_02461_),
    .X(net1960));
 sg13g2_buf_8 fanout1961 (.A(net1962),
    .X(net1961));
 sg13g2_buf_8 fanout1962 (.A(_02451_),
    .X(net1962));
 sg13g2_buf_8 fanout1963 (.A(_02440_),
    .X(net1963));
 sg13g2_buf_8 fanout1964 (.A(net1965),
    .X(net1964));
 sg13g2_buf_2 fanout1965 (.A(net1966),
    .X(net1965));
 sg13g2_buf_1 fanout1966 (.A(_02431_),
    .X(net1966));
 sg13g2_buf_8 fanout1967 (.A(_02421_),
    .X(net1967));
 sg13g2_buf_8 fanout1968 (.A(_02421_),
    .X(net1968));
 sg13g2_buf_8 fanout1969 (.A(net1970),
    .X(net1969));
 sg13g2_buf_8 fanout1970 (.A(_02411_),
    .X(net1970));
 sg13g2_buf_8 fanout1971 (.A(_02401_),
    .X(net1971));
 sg13g2_buf_8 fanout1972 (.A(_02401_),
    .X(net1972));
 sg13g2_buf_8 fanout1973 (.A(_02391_),
    .X(net1973));
 sg13g2_buf_8 fanout1974 (.A(_02391_),
    .X(net1974));
 sg13g2_buf_8 fanout1975 (.A(_02341_),
    .X(net1975));
 sg13g2_buf_8 fanout1976 (.A(_02341_),
    .X(net1976));
 sg13g2_buf_8 fanout1977 (.A(_02330_),
    .X(net1977));
 sg13g2_buf_8 fanout1978 (.A(net1979),
    .X(net1978));
 sg13g2_buf_8 fanout1979 (.A(_02320_),
    .X(net1979));
 sg13g2_buf_8 fanout1980 (.A(_02308_),
    .X(net1980));
 sg13g2_buf_8 fanout1981 (.A(net1982),
    .X(net1981));
 sg13g2_buf_8 fanout1982 (.A(_02289_),
    .X(net1982));
 sg13g2_buf_8 fanout1983 (.A(net1984),
    .X(net1983));
 sg13g2_buf_8 fanout1984 (.A(_02268_),
    .X(net1984));
 sg13g2_buf_8 fanout1985 (.A(_02257_),
    .X(net1985));
 sg13g2_buf_8 fanout1986 (.A(_02257_),
    .X(net1986));
 sg13g2_buf_8 fanout1987 (.A(net1988),
    .X(net1987));
 sg13g2_buf_8 fanout1988 (.A(_02247_),
    .X(net1988));
 sg13g2_buf_8 fanout1989 (.A(_02235_),
    .X(net1989));
 sg13g2_buf_8 fanout1990 (.A(_02225_),
    .X(net1990));
 sg13g2_buf_8 fanout1991 (.A(_02225_),
    .X(net1991));
 sg13g2_buf_8 fanout1992 (.A(_02168_),
    .X(net1992));
 sg13g2_buf_8 fanout1993 (.A(_02107_),
    .X(net1993));
 sg13g2_buf_8 fanout1994 (.A(net1995),
    .X(net1994));
 sg13g2_buf_2 fanout1995 (.A(net1996),
    .X(net1995));
 sg13g2_buf_1 fanout1996 (.A(_07130_),
    .X(net1996));
 sg13g2_buf_8 fanout1997 (.A(net1998),
    .X(net1997));
 sg13g2_buf_8 fanout1998 (.A(_06397_),
    .X(net1998));
 sg13g2_buf_8 fanout1999 (.A(net2000),
    .X(net1999));
 sg13g2_buf_8 fanout2000 (.A(_06225_),
    .X(net2000));
 sg13g2_buf_8 fanout2001 (.A(_06224_),
    .X(net2001));
 sg13g2_buf_8 fanout2002 (.A(net2005),
    .X(net2002));
 sg13g2_buf_8 fanout2003 (.A(net2004),
    .X(net2003));
 sg13g2_buf_2 fanout2004 (.A(net2005),
    .X(net2004));
 sg13g2_buf_8 fanout2005 (.A(_03488_),
    .X(net2005));
 sg13g2_buf_8 fanout2006 (.A(_02490_),
    .X(net2006));
 sg13g2_buf_8 fanout2007 (.A(_02460_),
    .X(net2007));
 sg13g2_buf_8 fanout2008 (.A(_02450_),
    .X(net2008));
 sg13g2_buf_8 fanout2009 (.A(_02430_),
    .X(net2009));
 sg13g2_buf_8 fanout2010 (.A(_02420_),
    .X(net2010));
 sg13g2_buf_8 fanout2011 (.A(_02410_),
    .X(net2011));
 sg13g2_buf_8 fanout2012 (.A(_02400_),
    .X(net2012));
 sg13g2_buf_8 fanout2013 (.A(_02390_),
    .X(net2013));
 sg13g2_buf_8 fanout2014 (.A(net2015),
    .X(net2014));
 sg13g2_buf_8 fanout2015 (.A(_02381_),
    .X(net2015));
 sg13g2_buf_8 fanout2016 (.A(net2017),
    .X(net2016));
 sg13g2_buf_8 fanout2017 (.A(_02371_),
    .X(net2017));
 sg13g2_buf_8 fanout2018 (.A(net2019),
    .X(net2018));
 sg13g2_buf_8 fanout2019 (.A(_02361_),
    .X(net2019));
 sg13g2_buf_8 fanout2020 (.A(_02351_),
    .X(net2020));
 sg13g2_buf_8 fanout2021 (.A(_02351_),
    .X(net2021));
 sg13g2_buf_8 fanout2022 (.A(_02340_),
    .X(net2022));
 sg13g2_buf_8 fanout2023 (.A(_02319_),
    .X(net2023));
 sg13g2_buf_8 fanout2024 (.A(net2025),
    .X(net2024));
 sg13g2_buf_8 fanout2025 (.A(_02299_),
    .X(net2025));
 sg13g2_buf_8 fanout2026 (.A(_02288_),
    .X(net2026));
 sg13g2_buf_8 fanout2027 (.A(net2028),
    .X(net2027));
 sg13g2_buf_8 fanout2028 (.A(_02278_),
    .X(net2028));
 sg13g2_buf_8 fanout2029 (.A(_02267_),
    .X(net2029));
 sg13g2_buf_8 fanout2030 (.A(_02256_),
    .X(net2030));
 sg13g2_buf_8 fanout2031 (.A(_02246_),
    .X(net2031));
 sg13g2_buf_8 fanout2032 (.A(_02224_),
    .X(net2032));
 sg13g2_buf_8 fanout2033 (.A(net2035),
    .X(net2033));
 sg13g2_buf_1 fanout2034 (.A(net2035),
    .X(net2034));
 sg13g2_buf_8 fanout2035 (.A(_02214_),
    .X(net2035));
 sg13g2_buf_8 fanout2036 (.A(net2037),
    .X(net2036));
 sg13g2_buf_8 fanout2037 (.A(_02204_),
    .X(net2037));
 sg13g2_buf_8 fanout2038 (.A(net2039),
    .X(net2038));
 sg13g2_buf_8 fanout2039 (.A(_02193_),
    .X(net2039));
 sg13g2_buf_8 fanout2040 (.A(_02183_),
    .X(net2040));
 sg13g2_buf_8 fanout2041 (.A(_02183_),
    .X(net2041));
 sg13g2_buf_8 fanout2042 (.A(_02159_),
    .X(net2042));
 sg13g2_buf_8 fanout2043 (.A(_02159_),
    .X(net2043));
 sg13g2_buf_8 fanout2044 (.A(net2045),
    .X(net2044));
 sg13g2_buf_1 fanout2045 (.A(net2046),
    .X(net2045));
 sg13g2_buf_1 fanout2046 (.A(_02149_),
    .X(net2046));
 sg13g2_buf_8 fanout2047 (.A(net2049),
    .X(net2047));
 sg13g2_buf_8 fanout2048 (.A(net2049),
    .X(net2048));
 sg13g2_buf_2 fanout2049 (.A(net2050),
    .X(net2049));
 sg13g2_buf_8 fanout2050 (.A(_07010_),
    .X(net2050));
 sg13g2_buf_8 fanout2051 (.A(_05498_),
    .X(net2051));
 sg13g2_buf_8 fanout2052 (.A(net2053),
    .X(net2052));
 sg13g2_buf_8 fanout2053 (.A(_05491_),
    .X(net2053));
 sg13g2_buf_8 fanout2054 (.A(_04903_),
    .X(net2054));
 sg13g2_buf_8 fanout2055 (.A(_04643_),
    .X(net2055));
 sg13g2_buf_8 fanout2056 (.A(_04642_),
    .X(net2056));
 sg13g2_buf_8 fanout2057 (.A(net2058),
    .X(net2057));
 sg13g2_buf_8 fanout2058 (.A(net2059),
    .X(net2058));
 sg13g2_buf_8 fanout2059 (.A(_04424_),
    .X(net2059));
 sg13g2_buf_8 fanout2060 (.A(net2061),
    .X(net2060));
 sg13g2_buf_8 fanout2061 (.A(net2062),
    .X(net2061));
 sg13g2_buf_8 fanout2062 (.A(_04422_),
    .X(net2062));
 sg13g2_buf_8 fanout2063 (.A(net2064),
    .X(net2063));
 sg13g2_buf_8 fanout2064 (.A(net2065),
    .X(net2064));
 sg13g2_buf_2 fanout2065 (.A(net2066),
    .X(net2065));
 sg13g2_buf_8 fanout2066 (.A(_04320_),
    .X(net2066));
 sg13g2_buf_8 fanout2067 (.A(net2068),
    .X(net2067));
 sg13g2_buf_8 fanout2068 (.A(net2069),
    .X(net2068));
 sg13g2_buf_2 fanout2069 (.A(_04320_),
    .X(net2069));
 sg13g2_buf_8 fanout2070 (.A(net2071),
    .X(net2070));
 sg13g2_buf_8 fanout2071 (.A(_04262_),
    .X(net2071));
 sg13g2_buf_2 fanout2072 (.A(net2073),
    .X(net2072));
 sg13g2_buf_8 fanout2073 (.A(net2074),
    .X(net2073));
 sg13g2_buf_8 fanout2074 (.A(_03482_),
    .X(net2074));
 sg13g2_buf_8 fanout2075 (.A(_03478_),
    .X(net2075));
 sg13g2_buf_8 fanout2076 (.A(_03468_),
    .X(net2076));
 sg13g2_buf_8 fanout2077 (.A(net2078),
    .X(net2077));
 sg13g2_buf_2 fanout2078 (.A(net2079),
    .X(net2078));
 sg13g2_buf_8 fanout2079 (.A(_03466_),
    .X(net2079));
 sg13g2_buf_8 fanout2080 (.A(_03455_),
    .X(net2080));
 sg13g2_buf_8 fanout2081 (.A(_03455_),
    .X(net2081));
 sg13g2_buf_8 fanout2082 (.A(_03446_),
    .X(net2082));
 sg13g2_buf_8 fanout2083 (.A(_03443_),
    .X(net2083));
 sg13g2_buf_2 fanout2084 (.A(_03443_),
    .X(net2084));
 sg13g2_buf_8 fanout2085 (.A(net2087),
    .X(net2085));
 sg13g2_buf_8 fanout2086 (.A(net2087),
    .X(net2086));
 sg13g2_buf_8 fanout2087 (.A(_03441_),
    .X(net2087));
 sg13g2_buf_8 fanout2088 (.A(_03441_),
    .X(net2088));
 sg13g2_buf_8 fanout2089 (.A(_03441_),
    .X(net2089));
 sg13g2_buf_8 fanout2090 (.A(_02380_),
    .X(net2090));
 sg13g2_buf_8 fanout2091 (.A(_02370_),
    .X(net2091));
 sg13g2_buf_8 fanout2092 (.A(_02360_),
    .X(net2092));
 sg13g2_buf_8 fanout2093 (.A(_02350_),
    .X(net2093));
 sg13g2_buf_8 fanout2094 (.A(_02298_),
    .X(net2094));
 sg13g2_buf_8 fanout2095 (.A(_02277_),
    .X(net2095));
 sg13g2_buf_8 fanout2096 (.A(_02213_),
    .X(net2096));
 sg13g2_buf_8 fanout2097 (.A(_02203_),
    .X(net2097));
 sg13g2_buf_8 fanout2098 (.A(_02192_),
    .X(net2098));
 sg13g2_buf_8 fanout2099 (.A(_02182_),
    .X(net2099));
 sg13g2_buf_8 fanout2100 (.A(_02158_),
    .X(net2100));
 sg13g2_buf_8 fanout2101 (.A(_02148_),
    .X(net2101));
 sg13g2_buf_8 fanout2102 (.A(_07201_),
    .X(net2102));
 sg13g2_buf_8 fanout2103 (.A(net2106),
    .X(net2103));
 sg13g2_buf_1 fanout2104 (.A(net2106),
    .X(net2104));
 sg13g2_buf_8 fanout2105 (.A(net2106),
    .X(net2105));
 sg13g2_buf_2 fanout2106 (.A(net2107),
    .X(net2106));
 sg13g2_buf_8 fanout2107 (.A(_04588_),
    .X(net2107));
 sg13g2_buf_8 fanout2108 (.A(_04587_),
    .X(net2108));
 sg13g2_buf_8 fanout2109 (.A(_04587_),
    .X(net2109));
 sg13g2_buf_8 fanout2110 (.A(net2112),
    .X(net2110));
 sg13g2_buf_2 fanout2111 (.A(net2112),
    .X(net2111));
 sg13g2_buf_8 fanout2112 (.A(_04421_),
    .X(net2112));
 sg13g2_buf_8 fanout2113 (.A(_04418_),
    .X(net2113));
 sg13g2_buf_8 fanout2114 (.A(_04272_),
    .X(net2114));
 sg13g2_buf_8 fanout2115 (.A(_04272_),
    .X(net2115));
 sg13g2_buf_8 fanout2116 (.A(net2118),
    .X(net2116));
 sg13g2_buf_1 fanout2117 (.A(net2118),
    .X(net2117));
 sg13g2_buf_8 fanout2118 (.A(_03433_),
    .X(net2118));
 sg13g2_buf_8 fanout2119 (.A(net2120),
    .X(net2119));
 sg13g2_buf_8 fanout2120 (.A(_03433_),
    .X(net2120));
 sg13g2_buf_8 fanout2121 (.A(net2122),
    .X(net2121));
 sg13g2_buf_8 fanout2122 (.A(net2123),
    .X(net2122));
 sg13g2_buf_1 fanout2123 (.A(_03432_),
    .X(net2123));
 sg13g2_buf_8 fanout2124 (.A(_03432_),
    .X(net2124));
 sg13g2_buf_8 fanout2125 (.A(_03432_),
    .X(net2125));
 sg13g2_buf_8 fanout2126 (.A(net2127),
    .X(net2126));
 sg13g2_buf_1 fanout2127 (.A(net2128),
    .X(net2127));
 sg13g2_buf_8 fanout2128 (.A(_02833_),
    .X(net2128));
 sg13g2_buf_8 fanout2129 (.A(net2130),
    .X(net2129));
 sg13g2_buf_8 fanout2130 (.A(net2131),
    .X(net2130));
 sg13g2_buf_8 fanout2131 (.A(_02832_),
    .X(net2131));
 sg13g2_buf_8 fanout2132 (.A(net2134),
    .X(net2132));
 sg13g2_buf_8 fanout2133 (.A(net2134),
    .X(net2133));
 sg13g2_buf_8 fanout2134 (.A(_02831_),
    .X(net2134));
 sg13g2_buf_8 fanout2135 (.A(net2136),
    .X(net2135));
 sg13g2_buf_2 fanout2136 (.A(net2137),
    .X(net2136));
 sg13g2_buf_8 fanout2137 (.A(_02830_),
    .X(net2137));
 sg13g2_buf_8 fanout2138 (.A(_02106_),
    .X(net2138));
 sg13g2_buf_8 fanout2139 (.A(_02106_),
    .X(net2139));
 sg13g2_buf_8 fanout2140 (.A(_02105_),
    .X(net2140));
 sg13g2_buf_8 fanout2141 (.A(_02105_),
    .X(net2141));
 sg13g2_buf_8 fanout2142 (.A(net2143),
    .X(net2142));
 sg13g2_buf_1 fanout2143 (.A(_07162_),
    .X(net2143));
 sg13g2_buf_8 fanout2144 (.A(net2146),
    .X(net2144));
 sg13g2_buf_1 fanout2145 (.A(net2146),
    .X(net2145));
 sg13g2_buf_8 fanout2146 (.A(_06905_),
    .X(net2146));
 sg13g2_buf_8 fanout2147 (.A(net2148),
    .X(net2147));
 sg13g2_buf_8 fanout2148 (.A(_06904_),
    .X(net2148));
 sg13g2_buf_8 fanout2149 (.A(net2151),
    .X(net2149));
 sg13g2_buf_1 fanout2150 (.A(net2151),
    .X(net2150));
 sg13g2_buf_8 fanout2151 (.A(net2152),
    .X(net2151));
 sg13g2_buf_8 fanout2152 (.A(net2155),
    .X(net2152));
 sg13g2_buf_8 fanout2153 (.A(net2154),
    .X(net2153));
 sg13g2_buf_8 fanout2154 (.A(net2155),
    .X(net2154));
 sg13g2_buf_8 fanout2155 (.A(_06730_),
    .X(net2155));
 sg13g2_buf_8 fanout2156 (.A(net2158),
    .X(net2156));
 sg13g2_buf_1 fanout2157 (.A(net2158),
    .X(net2157));
 sg13g2_buf_8 fanout2158 (.A(_06497_),
    .X(net2158));
 sg13g2_buf_8 fanout2159 (.A(_04632_),
    .X(net2159));
 sg13g2_buf_1 fanout2160 (.A(_04632_),
    .X(net2160));
 sg13g2_buf_8 fanout2161 (.A(_04626_),
    .X(net2161));
 sg13g2_buf_1 fanout2162 (.A(_04626_),
    .X(net2162));
 sg13g2_buf_8 fanout2163 (.A(_04623_),
    .X(net2163));
 sg13g2_buf_8 fanout2164 (.A(_04621_),
    .X(net2164));
 sg13g2_buf_8 fanout2165 (.A(_04620_),
    .X(net2165));
 sg13g2_buf_8 fanout2166 (.A(_04618_),
    .X(net2166));
 sg13g2_buf_8 fanout2167 (.A(net2168),
    .X(net2167));
 sg13g2_buf_8 fanout2168 (.A(_04608_),
    .X(net2168));
 sg13g2_buf_8 fanout2169 (.A(net2170),
    .X(net2169));
 sg13g2_buf_8 fanout2170 (.A(_04606_),
    .X(net2170));
 sg13g2_buf_8 fanout2171 (.A(net2172),
    .X(net2171));
 sg13g2_buf_2 fanout2172 (.A(net2173),
    .X(net2172));
 sg13g2_buf_1 fanout2173 (.A(_04585_),
    .X(net2173));
 sg13g2_buf_8 fanout2174 (.A(net2175),
    .X(net2174));
 sg13g2_buf_8 fanout2175 (.A(net2177),
    .X(net2175));
 sg13g2_buf_8 fanout2176 (.A(net2177),
    .X(net2176));
 sg13g2_buf_8 fanout2177 (.A(_03435_),
    .X(net2177));
 sg13g2_buf_8 fanout2178 (.A(_03194_),
    .X(net2178));
 sg13g2_buf_8 fanout2179 (.A(net2180),
    .X(net2179));
 sg13g2_buf_8 fanout2180 (.A(net2181),
    .X(net2180));
 sg13g2_buf_8 fanout2181 (.A(_02116_),
    .X(net2181));
 sg13g2_buf_8 fanout2182 (.A(net2184),
    .X(net2182));
 sg13g2_buf_2 fanout2183 (.A(net2184),
    .X(net2183));
 sg13g2_buf_2 fanout2184 (.A(_02116_),
    .X(net2184));
 sg13g2_buf_8 fanout2185 (.A(net2187),
    .X(net2185));
 sg13g2_buf_2 fanout2186 (.A(net2187),
    .X(net2186));
 sg13g2_buf_8 fanout2187 (.A(_06893_),
    .X(net2187));
 sg13g2_buf_8 fanout2188 (.A(net2190),
    .X(net2188));
 sg13g2_buf_1 fanout2189 (.A(net2190),
    .X(net2189));
 sg13g2_buf_1 fanout2190 (.A(_06879_),
    .X(net2190));
 sg13g2_buf_8 fanout2191 (.A(net2194),
    .X(net2191));
 sg13g2_buf_8 fanout2192 (.A(net2194),
    .X(net2192));
 sg13g2_buf_8 fanout2193 (.A(net2194),
    .X(net2193));
 sg13g2_buf_8 fanout2194 (.A(_06415_),
    .X(net2194));
 sg13g2_buf_8 fanout2195 (.A(net2196),
    .X(net2195));
 sg13g2_buf_2 fanout2196 (.A(net2201),
    .X(net2196));
 sg13g2_buf_8 fanout2197 (.A(net2199),
    .X(net2197));
 sg13g2_buf_1 fanout2198 (.A(net2199),
    .X(net2198));
 sg13g2_buf_8 fanout2199 (.A(net2201),
    .X(net2199));
 sg13g2_buf_8 fanout2200 (.A(net2201),
    .X(net2200));
 sg13g2_buf_8 fanout2201 (.A(net2202),
    .X(net2201));
 sg13g2_buf_8 fanout2202 (.A(net2218),
    .X(net2202));
 sg13g2_buf_8 fanout2203 (.A(net2204),
    .X(net2203));
 sg13g2_buf_8 fanout2204 (.A(net2210),
    .X(net2204));
 sg13g2_buf_8 fanout2205 (.A(net2206),
    .X(net2205));
 sg13g2_buf_8 fanout2206 (.A(net2208),
    .X(net2206));
 sg13g2_buf_8 fanout2207 (.A(net2208),
    .X(net2207));
 sg13g2_buf_8 fanout2208 (.A(net2209),
    .X(net2208));
 sg13g2_buf_8 fanout2209 (.A(net2210),
    .X(net2209));
 sg13g2_buf_8 fanout2210 (.A(net2218),
    .X(net2210));
 sg13g2_buf_8 fanout2211 (.A(net2213),
    .X(net2211));
 sg13g2_buf_8 fanout2212 (.A(net2213),
    .X(net2212));
 sg13g2_buf_8 fanout2213 (.A(net2218),
    .X(net2213));
 sg13g2_buf_8 fanout2214 (.A(net2215),
    .X(net2214));
 sg13g2_buf_8 fanout2215 (.A(net2217),
    .X(net2215));
 sg13g2_buf_8 fanout2216 (.A(net2217),
    .X(net2216));
 sg13g2_buf_8 fanout2217 (.A(net2218),
    .X(net2217));
 sg13g2_buf_8 fanout2218 (.A(_06414_),
    .X(net2218));
 sg13g2_buf_8 fanout2219 (.A(_06411_),
    .X(net2219));
 sg13g2_buf_8 fanout2220 (.A(_06385_),
    .X(net2220));
 sg13g2_buf_8 fanout2221 (.A(_05973_),
    .X(net2221));
 sg13g2_buf_8 fanout2222 (.A(_05388_),
    .X(net2222));
 sg13g2_buf_1 fanout2223 (.A(_05388_),
    .X(net2223));
 sg13g2_buf_8 fanout2224 (.A(_05323_),
    .X(net2224));
 sg13g2_buf_1 fanout2225 (.A(_05323_),
    .X(net2225));
 sg13g2_buf_8 fanout2226 (.A(_05290_),
    .X(net2226));
 sg13g2_buf_1 fanout2227 (.A(_05290_),
    .X(net2227));
 sg13g2_buf_8 fanout2228 (.A(_04899_),
    .X(net2228));
 sg13g2_buf_8 fanout2229 (.A(net2232),
    .X(net2229));
 sg13g2_buf_8 fanout2230 (.A(net2231),
    .X(net2230));
 sg13g2_buf_2 fanout2231 (.A(net2232),
    .X(net2231));
 sg13g2_buf_2 fanout2232 (.A(_04876_),
    .X(net2232));
 sg13g2_buf_8 fanout2233 (.A(_04876_),
    .X(net2233));
 sg13g2_buf_8 fanout2234 (.A(_04876_),
    .X(net2234));
 sg13g2_buf_8 fanout2235 (.A(net2237),
    .X(net2235));
 sg13g2_buf_8 fanout2236 (.A(net2237),
    .X(net2236));
 sg13g2_buf_8 fanout2237 (.A(_04584_),
    .X(net2237));
 sg13g2_buf_8 fanout2238 (.A(_04584_),
    .X(net2238));
 sg13g2_buf_8 fanout2239 (.A(_04584_),
    .X(net2239));
 sg13g2_buf_8 fanout2240 (.A(net2242),
    .X(net2240));
 sg13g2_buf_1 fanout2241 (.A(net2242),
    .X(net2241));
 sg13g2_buf_1 fanout2242 (.A(_02820_),
    .X(net2242));
 sg13g2_buf_8 fanout2243 (.A(net2245),
    .X(net2243));
 sg13g2_buf_8 fanout2244 (.A(net2245),
    .X(net2244));
 sg13g2_buf_8 fanout2245 (.A(net2247),
    .X(net2245));
 sg13g2_buf_8 fanout2246 (.A(net2247),
    .X(net2246));
 sg13g2_buf_8 fanout2247 (.A(_02144_),
    .X(net2247));
 sg13g2_buf_8 fanout2248 (.A(net2252),
    .X(net2248));
 sg13g2_buf_8 fanout2249 (.A(net2252),
    .X(net2249));
 sg13g2_buf_8 fanout2250 (.A(net2252),
    .X(net2250));
 sg13g2_buf_8 fanout2251 (.A(net2252),
    .X(net2251));
 sg13g2_buf_8 fanout2252 (.A(_02140_),
    .X(net2252));
 sg13g2_buf_8 fanout2253 (.A(net2254),
    .X(net2253));
 sg13g2_buf_8 fanout2254 (.A(net2257),
    .X(net2254));
 sg13g2_buf_8 fanout2255 (.A(net2256),
    .X(net2255));
 sg13g2_buf_8 fanout2256 (.A(net2257),
    .X(net2256));
 sg13g2_buf_8 fanout2257 (.A(_02136_),
    .X(net2257));
 sg13g2_buf_8 fanout2258 (.A(_02132_),
    .X(net2258));
 sg13g2_buf_2 fanout2259 (.A(_02132_),
    .X(net2259));
 sg13g2_buf_8 fanout2260 (.A(net2262),
    .X(net2260));
 sg13g2_buf_8 fanout2261 (.A(net2262),
    .X(net2261));
 sg13g2_buf_8 fanout2262 (.A(_02132_),
    .X(net2262));
 sg13g2_buf_8 fanout2263 (.A(net2267),
    .X(net2263));
 sg13g2_buf_8 fanout2264 (.A(net2267),
    .X(net2264));
 sg13g2_buf_8 fanout2265 (.A(net2267),
    .X(net2265));
 sg13g2_buf_2 fanout2266 (.A(net2267),
    .X(net2266));
 sg13g2_buf_8 fanout2267 (.A(_02128_),
    .X(net2267));
 sg13g2_buf_8 fanout2268 (.A(net2273),
    .X(net2268));
 sg13g2_buf_8 fanout2269 (.A(net2272),
    .X(net2269));
 sg13g2_buf_8 fanout2270 (.A(net2271),
    .X(net2270));
 sg13g2_buf_8 fanout2271 (.A(net2272),
    .X(net2271));
 sg13g2_buf_8 fanout2272 (.A(net2273),
    .X(net2272));
 sg13g2_buf_8 fanout2273 (.A(_02124_),
    .X(net2273));
 sg13g2_buf_8 fanout2274 (.A(net2275),
    .X(net2274));
 sg13g2_buf_8 fanout2275 (.A(net2279),
    .X(net2275));
 sg13g2_buf_8 fanout2276 (.A(net2278),
    .X(net2276));
 sg13g2_buf_1 fanout2277 (.A(net2278),
    .X(net2277));
 sg13g2_buf_8 fanout2278 (.A(net2279),
    .X(net2278));
 sg13g2_buf_8 fanout2279 (.A(_02120_),
    .X(net2279));
 sg13g2_buf_8 fanout2280 (.A(_06387_),
    .X(net2280));
 sg13g2_buf_8 fanout2281 (.A(net2282),
    .X(net2281));
 sg13g2_buf_8 fanout2282 (.A(_05972_),
    .X(net2282));
 sg13g2_buf_8 fanout2283 (.A(_05372_),
    .X(net2283));
 sg13g2_buf_8 fanout2284 (.A(_04896_),
    .X(net2284));
 sg13g2_buf_8 fanout2285 (.A(_04757_),
    .X(net2285));
 sg13g2_buf_8 fanout2286 (.A(_04745_),
    .X(net2286));
 sg13g2_buf_8 fanout2287 (.A(net2288),
    .X(net2287));
 sg13g2_buf_8 fanout2288 (.A(_04581_),
    .X(net2288));
 sg13g2_buf_8 fanout2289 (.A(net2291),
    .X(net2289));
 sg13g2_buf_8 fanout2290 (.A(net2291),
    .X(net2290));
 sg13g2_buf_8 fanout2291 (.A(_04580_),
    .X(net2291));
 sg13g2_buf_8 fanout2292 (.A(net2293),
    .X(net2292));
 sg13g2_buf_8 fanout2293 (.A(net2295),
    .X(net2293));
 sg13g2_buf_8 fanout2294 (.A(net2295),
    .X(net2294));
 sg13g2_buf_8 fanout2295 (.A(_04571_),
    .X(net2295));
 sg13g2_buf_8 fanout2296 (.A(net2297),
    .X(net2296));
 sg13g2_buf_8 fanout2297 (.A(net2298),
    .X(net2297));
 sg13g2_buf_8 fanout2298 (.A(_04570_),
    .X(net2298));
 sg13g2_buf_8 fanout2299 (.A(net2300),
    .X(net2299));
 sg13g2_buf_8 fanout2300 (.A(_04566_),
    .X(net2300));
 sg13g2_buf_1 fanout2301 (.A(_04566_),
    .X(net2301));
 sg13g2_buf_8 fanout2302 (.A(_04302_),
    .X(net2302));
 sg13g2_buf_1 fanout2303 (.A(_04302_),
    .X(net2303));
 sg13g2_buf_8 fanout2304 (.A(net2305),
    .X(net2304));
 sg13g2_buf_1 fanout2305 (.A(net2306),
    .X(net2305));
 sg13g2_buf_8 fanout2306 (.A(net2307),
    .X(net2306));
 sg13g2_buf_8 fanout2307 (.A(_03538_),
    .X(net2307));
 sg13g2_buf_8 fanout2308 (.A(_03537_),
    .X(net2308));
 sg13g2_buf_8 fanout2309 (.A(_03537_),
    .X(net2309));
 sg13g2_buf_8 fanout2310 (.A(_03458_),
    .X(net2310));
 sg13g2_buf_8 fanout2311 (.A(net2312),
    .X(net2311));
 sg13g2_buf_8 fanout2312 (.A(_03187_),
    .X(net2312));
 sg13g2_buf_8 fanout2313 (.A(_03186_),
    .X(net2313));
 sg13g2_buf_1 fanout2314 (.A(_03186_),
    .X(net2314));
 sg13g2_buf_8 fanout2315 (.A(_02770_),
    .X(net2315));
 sg13g2_buf_8 fanout2316 (.A(_02770_),
    .X(net2316));
 sg13g2_buf_8 fanout2317 (.A(_02769_),
    .X(net2317));
 sg13g2_buf_8 fanout2318 (.A(net2319),
    .X(net2318));
 sg13g2_buf_8 fanout2319 (.A(_02740_),
    .X(net2319));
 sg13g2_buf_8 fanout2320 (.A(net2321),
    .X(net2320));
 sg13g2_buf_8 fanout2321 (.A(_02739_),
    .X(net2321));
 sg13g2_buf_8 fanout2322 (.A(_02708_),
    .X(net2322));
 sg13g2_buf_8 fanout2323 (.A(_02548_),
    .X(net2323));
 sg13g2_buf_2 fanout2324 (.A(_02548_),
    .X(net2324));
 sg13g2_buf_8 fanout2325 (.A(_02473_),
    .X(net2325));
 sg13g2_buf_8 fanout2326 (.A(_02472_),
    .X(net2326));
 sg13g2_buf_8 fanout2327 (.A(net2328),
    .X(net2327));
 sg13g2_buf_8 fanout2328 (.A(net2331),
    .X(net2328));
 sg13g2_buf_8 fanout2329 (.A(net2330),
    .X(net2329));
 sg13g2_buf_8 fanout2330 (.A(net2331),
    .X(net2330));
 sg13g2_buf_8 fanout2331 (.A(_02090_),
    .X(net2331));
 sg13g2_buf_8 fanout2332 (.A(_05364_),
    .X(net2332));
 sg13g2_buf_2 fanout2333 (.A(net2334),
    .X(net2333));
 sg13g2_buf_2 fanout2334 (.A(_04895_),
    .X(net2334));
 sg13g2_buf_8 fanout2335 (.A(net2336),
    .X(net2335));
 sg13g2_buf_8 fanout2336 (.A(_04894_),
    .X(net2336));
 sg13g2_buf_8 fanout2337 (.A(_04759_),
    .X(net2337));
 sg13g2_buf_8 fanout2338 (.A(net2339),
    .X(net2338));
 sg13g2_buf_2 fanout2339 (.A(net2340),
    .X(net2339));
 sg13g2_buf_1 fanout2340 (.A(net2341),
    .X(net2340));
 sg13g2_buf_8 fanout2341 (.A(_03464_),
    .X(net2341));
 sg13g2_buf_8 fanout2342 (.A(net2344),
    .X(net2342));
 sg13g2_buf_1 fanout2343 (.A(net2344),
    .X(net2343));
 sg13g2_buf_1 fanout2344 (.A(net2347),
    .X(net2344));
 sg13g2_buf_8 fanout2345 (.A(net2346),
    .X(net2345));
 sg13g2_buf_8 fanout2346 (.A(net2347),
    .X(net2346));
 sg13g2_buf_8 fanout2347 (.A(_03459_),
    .X(net2347));
 sg13g2_buf_8 fanout2348 (.A(net2349),
    .X(net2348));
 sg13g2_buf_2 fanout2349 (.A(_03457_),
    .X(net2349));
 sg13g2_buf_8 fanout2350 (.A(net2351),
    .X(net2350));
 sg13g2_buf_8 fanout2351 (.A(_03457_),
    .X(net2351));
 sg13g2_buf_8 fanout2352 (.A(net2354),
    .X(net2352));
 sg13g2_buf_1 fanout2353 (.A(net2354),
    .X(net2353));
 sg13g2_buf_8 fanout2354 (.A(net2356),
    .X(net2354));
 sg13g2_buf_8 fanout2355 (.A(net2356),
    .X(net2355));
 sg13g2_buf_8 fanout2356 (.A(_03388_),
    .X(net2356));
 sg13g2_buf_8 fanout2357 (.A(_02807_),
    .X(net2357));
 sg13g2_buf_8 fanout2358 (.A(net2359),
    .X(net2358));
 sg13g2_buf_8 fanout2359 (.A(net2360),
    .X(net2359));
 sg13g2_buf_8 fanout2360 (.A(_02563_),
    .X(net2360));
 sg13g2_buf_8 fanout2361 (.A(net2362),
    .X(net2361));
 sg13g2_buf_2 fanout2362 (.A(net2363),
    .X(net2362));
 sg13g2_buf_2 fanout2363 (.A(net2364),
    .X(net2363));
 sg13g2_buf_8 fanout2364 (.A(_02562_),
    .X(net2364));
 sg13g2_buf_8 fanout2365 (.A(_02555_),
    .X(net2365));
 sg13g2_buf_8 fanout2366 (.A(_02544_),
    .X(net2366));
 sg13g2_buf_8 fanout2367 (.A(net2368),
    .X(net2367));
 sg13g2_buf_8 fanout2368 (.A(net2369),
    .X(net2368));
 sg13g2_buf_8 fanout2369 (.A(_02543_),
    .X(net2369));
 sg13g2_buf_8 fanout2370 (.A(net2371),
    .X(net2370));
 sg13g2_buf_8 fanout2371 (.A(_02541_),
    .X(net2371));
 sg13g2_buf_8 fanout2372 (.A(net2375),
    .X(net2372));
 sg13g2_buf_1 fanout2373 (.A(net2375),
    .X(net2373));
 sg13g2_buf_8 fanout2374 (.A(net2375),
    .X(net2374));
 sg13g2_buf_8 fanout2375 (.A(_02540_),
    .X(net2375));
 sg13g2_buf_8 fanout2376 (.A(net2377),
    .X(net2376));
 sg13g2_buf_8 fanout2377 (.A(net2378),
    .X(net2377));
 sg13g2_buf_8 fanout2378 (.A(_02538_),
    .X(net2378));
 sg13g2_buf_8 fanout2379 (.A(_02523_),
    .X(net2379));
 sg13g2_buf_8 fanout2380 (.A(_02523_),
    .X(net2380));
 sg13g2_buf_8 fanout2381 (.A(net2383),
    .X(net2381));
 sg13g2_buf_8 fanout2382 (.A(net2383),
    .X(net2382));
 sg13g2_buf_8 fanout2383 (.A(net2384),
    .X(net2383));
 sg13g2_buf_8 fanout2384 (.A(_02522_),
    .X(net2384));
 sg13g2_buf_8 fanout2385 (.A(_02510_),
    .X(net2385));
 sg13g2_buf_8 fanout2386 (.A(_02505_),
    .X(net2386));
 sg13g2_buf_8 fanout2387 (.A(net2388),
    .X(net2387));
 sg13g2_buf_8 fanout2388 (.A(_02471_),
    .X(net2388));
 sg13g2_buf_8 fanout2389 (.A(net2390),
    .X(net2389));
 sg13g2_buf_8 fanout2390 (.A(_02470_),
    .X(net2390));
 sg13g2_buf_8 fanout2391 (.A(net2395),
    .X(net2391));
 sg13g2_buf_1 fanout2392 (.A(net2395),
    .X(net2392));
 sg13g2_buf_8 fanout2393 (.A(net2395),
    .X(net2393));
 sg13g2_buf_1 fanout2394 (.A(net2395),
    .X(net2394));
 sg13g2_buf_2 fanout2395 (.A(_02113_),
    .X(net2395));
 sg13g2_buf_8 fanout2396 (.A(net2397),
    .X(net2396));
 sg13g2_buf_8 fanout2397 (.A(net2398),
    .X(net2397));
 sg13g2_buf_8 fanout2398 (.A(_02112_),
    .X(net2398));
 sg13g2_buf_8 fanout2399 (.A(_02111_),
    .X(net2399));
 sg13g2_buf_8 fanout2400 (.A(_02110_),
    .X(net2400));
 sg13g2_buf_8 fanout2401 (.A(_02110_),
    .X(net2401));
 sg13g2_buf_8 fanout2402 (.A(net2405),
    .X(net2402));
 sg13g2_buf_8 fanout2403 (.A(net2405),
    .X(net2403));
 sg13g2_buf_1 fanout2404 (.A(net2405),
    .X(net2404));
 sg13g2_buf_2 fanout2405 (.A(_02109_),
    .X(net2405));
 sg13g2_buf_2 fanout2406 (.A(net2407),
    .X(net2406));
 sg13g2_buf_8 fanout2407 (.A(net2409),
    .X(net2407));
 sg13g2_buf_8 fanout2408 (.A(net2409),
    .X(net2408));
 sg13g2_buf_8 fanout2409 (.A(_02068_),
    .X(net2409));
 sg13g2_buf_8 fanout2410 (.A(_02038_),
    .X(net2410));
 sg13g2_buf_8 fanout2411 (.A(net2412),
    .X(net2411));
 sg13g2_buf_8 fanout2412 (.A(net2413),
    .X(net2412));
 sg13g2_buf_8 fanout2413 (.A(net2431),
    .X(net2413));
 sg13g2_buf_8 fanout2414 (.A(net2417),
    .X(net2414));
 sg13g2_buf_8 fanout2415 (.A(net2417),
    .X(net2415));
 sg13g2_buf_1 fanout2416 (.A(net2417),
    .X(net2416));
 sg13g2_buf_8 fanout2417 (.A(net2431),
    .X(net2417));
 sg13g2_buf_8 fanout2418 (.A(net2419),
    .X(net2418));
 sg13g2_buf_8 fanout2419 (.A(net2430),
    .X(net2419));
 sg13g2_buf_8 fanout2420 (.A(net2421),
    .X(net2420));
 sg13g2_buf_8 fanout2421 (.A(net2430),
    .X(net2421));
 sg13g2_buf_8 fanout2422 (.A(net2423),
    .X(net2422));
 sg13g2_buf_8 fanout2423 (.A(net2424),
    .X(net2423));
 sg13g2_buf_8 fanout2424 (.A(net2430),
    .X(net2424));
 sg13g2_buf_8 fanout2425 (.A(net2427),
    .X(net2425));
 sg13g2_buf_1 fanout2426 (.A(net2427),
    .X(net2426));
 sg13g2_buf_8 fanout2427 (.A(net2428),
    .X(net2427));
 sg13g2_buf_8 fanout2428 (.A(net2429),
    .X(net2428));
 sg13g2_buf_8 fanout2429 (.A(net2430),
    .X(net2429));
 sg13g2_buf_8 fanout2430 (.A(net2431),
    .X(net2430));
 sg13g2_buf_8 fanout2431 (.A(_02012_),
    .X(net2431));
 sg13g2_buf_8 fanout2432 (.A(net2434),
    .X(net2432));
 sg13g2_buf_2 fanout2433 (.A(net2434),
    .X(net2433));
 sg13g2_buf_8 fanout2434 (.A(_01992_),
    .X(net2434));
 sg13g2_buf_8 fanout2435 (.A(net2436),
    .X(net2435));
 sg13g2_buf_8 fanout2436 (.A(net2437),
    .X(net2436));
 sg13g2_buf_8 fanout2437 (.A(_01990_),
    .X(net2437));
 sg13g2_buf_8 fanout2438 (.A(_01989_),
    .X(net2438));
 sg13g2_buf_8 fanout2439 (.A(_01981_),
    .X(net2439));
 sg13g2_buf_8 fanout2440 (.A(net2441),
    .X(net2440));
 sg13g2_buf_8 fanout2441 (.A(_01967_),
    .X(net2441));
 sg13g2_buf_8 fanout2442 (.A(net2443),
    .X(net2442));
 sg13g2_buf_8 fanout2443 (.A(_01960_),
    .X(net2443));
 sg13g2_buf_8 fanout2444 (.A(net2451),
    .X(net2444));
 sg13g2_buf_1 fanout2445 (.A(net2451),
    .X(net2445));
 sg13g2_buf_8 fanout2446 (.A(net2451),
    .X(net2446));
 sg13g2_buf_8 fanout2447 (.A(net2448),
    .X(net2447));
 sg13g2_buf_8 fanout2448 (.A(net2449),
    .X(net2448));
 sg13g2_buf_8 fanout2449 (.A(net2450),
    .X(net2449));
 sg13g2_buf_8 fanout2450 (.A(net2451),
    .X(net2450));
 sg13g2_buf_8 fanout2451 (.A(_01960_),
    .X(net2451));
 sg13g2_buf_8 fanout2452 (.A(_01778_),
    .X(net2452));
 sg13g2_buf_8 fanout2453 (.A(_01776_),
    .X(net2453));
 sg13g2_buf_8 fanout2454 (.A(net2458),
    .X(net2454));
 sg13g2_buf_8 fanout2455 (.A(net2456),
    .X(net2455));
 sg13g2_buf_8 fanout2456 (.A(net2457),
    .X(net2456));
 sg13g2_buf_2 fanout2457 (.A(net2458),
    .X(net2457));
 sg13g2_buf_1 fanout2458 (.A(net5253),
    .X(net2458));
 sg13g2_buf_2 fanout2459 (.A(net5339),
    .X(net2459));
 sg13g2_buf_8 fanout2460 (.A(net5335),
    .X(net2460));
 sg13g2_buf_8 fanout2461 (.A(net5349),
    .X(net2461));
 sg13g2_buf_8 fanout2462 (.A(net2463),
    .X(net2462));
 sg13g2_buf_1 fanout2463 (.A(net5378),
    .X(net2463));
 sg13g2_buf_8 fanout2464 (.A(net4377),
    .X(net2464));
 sg13g2_buf_8 fanout2465 (.A(net5312),
    .X(net2465));
 sg13g2_buf_8 fanout2466 (.A(net5368),
    .X(net2466));
 sg13g2_buf_8 fanout2467 (.A(net2469),
    .X(net2467));
 sg13g2_buf_1 fanout2468 (.A(net2469),
    .X(net2468));
 sg13g2_buf_1 fanout2469 (.A(net2471),
    .X(net2469));
 sg13g2_buf_8 fanout2470 (.A(net2471),
    .X(net2470));
 sg13g2_buf_8 fanout2471 (.A(\addr[26] ),
    .X(net2471));
 sg13g2_buf_8 fanout2472 (.A(net5196),
    .X(net2472));
 sg13g2_buf_8 fanout2473 (.A(net2474),
    .X(net2473));
 sg13g2_buf_8 fanout2474 (.A(net2475),
    .X(net2474));
 sg13g2_buf_8 fanout2475 (.A(net2476),
    .X(net2475));
 sg13g2_buf_8 fanout2476 (.A(net5377),
    .X(net2476));
 sg13g2_buf_8 fanout2477 (.A(net2480),
    .X(net2477));
 sg13g2_buf_2 fanout2478 (.A(net2480),
    .X(net2478));
 sg13g2_buf_8 fanout2479 (.A(net2480),
    .X(net2479));
 sg13g2_buf_2 fanout2480 (.A(net2482),
    .X(net2480));
 sg13g2_buf_8 fanout2481 (.A(net2482),
    .X(net2481));
 sg13g2_buf_1 fanout2482 (.A(net2487),
    .X(net2482));
 sg13g2_buf_2 fanout2483 (.A(net2487),
    .X(net2483));
 sg13g2_buf_1 fanout2484 (.A(net2487),
    .X(net2484));
 sg13g2_buf_2 fanout2485 (.A(net2486),
    .X(net2485));
 sg13g2_buf_1 fanout2486 (.A(net2487),
    .X(net2486));
 sg13g2_buf_8 fanout2487 (.A(net5275),
    .X(net2487));
 sg13g2_buf_8 fanout2488 (.A(net2489),
    .X(net2488));
 sg13g2_buf_8 fanout2489 (.A(net2490),
    .X(net2489));
 sg13g2_buf_1 fanout2490 (.A(\i_seal.read_seq[1] ),
    .X(net2490));
 sg13g2_buf_8 fanout2491 (.A(net2492),
    .X(net2491));
 sg13g2_buf_2 fanout2492 (.A(\i_seal.read_seq[1] ),
    .X(net2492));
 sg13g2_buf_8 fanout2493 (.A(\i_seal.byte_idx[0] ),
    .X(net2493));
 sg13g2_buf_8 fanout2494 (.A(net2497),
    .X(net2494));
 sg13g2_buf_8 fanout2495 (.A(net2497),
    .X(net2495));
 sg13g2_buf_8 fanout2496 (.A(net2497),
    .X(net2496));
 sg13g2_buf_8 fanout2497 (.A(net2503),
    .X(net2497));
 sg13g2_buf_8 fanout2498 (.A(net2500),
    .X(net2498));
 sg13g2_buf_2 fanout2499 (.A(net2500),
    .X(net2499));
 sg13g2_buf_8 fanout2500 (.A(net2503),
    .X(net2500));
 sg13g2_buf_8 fanout2501 (.A(net2503),
    .X(net2501));
 sg13g2_buf_2 fanout2502 (.A(net2503),
    .X(net2502));
 sg13g2_buf_8 fanout2503 (.A(net5032),
    .X(net2503));
 sg13g2_buf_8 fanout2504 (.A(net5313),
    .X(net2504));
 sg13g2_buf_8 fanout2505 (.A(net5227),
    .X(net2505));
 sg13g2_buf_8 fanout2506 (.A(net5303),
    .X(net2506));
 sg13g2_buf_8 fanout2507 (.A(net5257),
    .X(net2507));
 sg13g2_buf_1 fanout2508 (.A(net5257),
    .X(net2508));
 sg13g2_buf_8 fanout2509 (.A(net2512),
    .X(net2509));
 sg13g2_buf_8 fanout2510 (.A(net2511),
    .X(net2510));
 sg13g2_buf_8 fanout2511 (.A(net2512),
    .X(net2511));
 sg13g2_buf_8 fanout2512 (.A(net5338),
    .X(net2512));
 sg13g2_buf_8 fanout2513 (.A(net5283),
    .X(net2513));
 sg13g2_buf_8 fanout2514 (.A(net5265),
    .X(net2514));
 sg13g2_buf_8 fanout2515 (.A(net5311),
    .X(net2515));
 sg13g2_buf_8 fanout2516 (.A(net2517),
    .X(net2516));
 sg13g2_buf_1 fanout2517 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .X(net2517));
 sg13g2_buf_8 fanout2518 (.A(net2519),
    .X(net2518));
 sg13g2_buf_8 fanout2519 (.A(net2520),
    .X(net2519));
 sg13g2_buf_8 fanout2520 (.A(net2526),
    .X(net2520));
 sg13g2_buf_2 fanout2521 (.A(net2522),
    .X(net2521));
 sg13g2_buf_2 fanout2522 (.A(net2523),
    .X(net2522));
 sg13g2_buf_8 fanout2523 (.A(net2525),
    .X(net2523));
 sg13g2_buf_8 fanout2524 (.A(net2525),
    .X(net2524));
 sg13g2_buf_8 fanout2525 (.A(net2526),
    .X(net2525));
 sg13g2_buf_8 fanout2526 (.A(net5274),
    .X(net2526));
 sg13g2_buf_8 fanout2527 (.A(net2528),
    .X(net2527));
 sg13g2_buf_8 fanout2528 (.A(\i_tinyqv.cpu.alu_op[1] ),
    .X(net2528));
 sg13g2_buf_8 fanout2529 (.A(net2530),
    .X(net2529));
 sg13g2_buf_8 fanout2530 (.A(net5379),
    .X(net2530));
 sg13g2_buf_8 fanout2531 (.A(net5371),
    .X(net2531));
 sg13g2_buf_8 fanout2532 (.A(\i_tinyqv.cpu.counter[4] ),
    .X(net2532));
 sg13g2_buf_8 fanout2533 (.A(\i_tinyqv.cpu.counter[4] ),
    .X(net2533));
 sg13g2_buf_8 fanout2534 (.A(net2536),
    .X(net2534));
 sg13g2_buf_2 fanout2535 (.A(net2536),
    .X(net2535));
 sg13g2_buf_8 fanout2536 (.A(\i_tinyqv.cpu.counter[4] ),
    .X(net2536));
 sg13g2_buf_8 fanout2537 (.A(net2538),
    .X(net2537));
 sg13g2_buf_1 fanout2538 (.A(\i_tinyqv.cpu.counter[3] ),
    .X(net2538));
 sg13g2_buf_8 fanout2539 (.A(net2540),
    .X(net2539));
 sg13g2_buf_8 fanout2540 (.A(net5360),
    .X(net2540));
 sg13g2_buf_8 fanout2541 (.A(net2542),
    .X(net2541));
 sg13g2_buf_8 fanout2542 (.A(\i_tinyqv.cpu.counter[2] ),
    .X(net2542));
 sg13g2_buf_8 fanout2543 (.A(net5184),
    .X(net2543));
 sg13g2_buf_8 fanout2544 (.A(net4976),
    .X(net2544));
 sg13g2_buf_8 fanout2545 (.A(\i_i2c_peri.i_i2c.state_reg[1] ),
    .X(net2545));
 sg13g2_buf_8 fanout2546 (.A(net5358),
    .X(net2546));
 sg13g2_buf_8 fanout2547 (.A(net5373),
    .X(net2547));
 sg13g2_buf_8 fanout2548 (.A(net4982),
    .X(net2548));
 sg13g2_buf_8 fanout2549 (.A(net2550),
    .X(net2549));
 sg13g2_buf_8 fanout2550 (.A(net4169),
    .X(net2550));
 sg13g2_buf_8 fanout2551 (.A(net4896),
    .X(net2551));
 sg13g2_buf_8 fanout2552 (.A(net4708),
    .X(net2552));
 sg13g2_buf_8 fanout2553 (.A(net4814),
    .X(net2553));
 sg13g2_buf_8 fanout2554 (.A(net4793),
    .X(net2554));
 sg13g2_buf_8 fanout2555 (.A(net4848),
    .X(net2555));
 sg13g2_buf_8 fanout2556 (.A(net5012),
    .X(net2556));
 sg13g2_buf_8 fanout2557 (.A(net5015),
    .X(net2557));
 sg13g2_buf_2 fanout2558 (.A(net5015),
    .X(net2558));
 sg13g2_buf_8 fanout2559 (.A(net4681),
    .X(net2559));
 sg13g2_buf_8 fanout2560 (.A(net2562),
    .X(net2560));
 sg13g2_buf_1 fanout2561 (.A(net2562),
    .X(net2561));
 sg13g2_buf_8 fanout2562 (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(net2562));
 sg13g2_buf_8 fanout2563 (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(net2563));
 sg13g2_buf_2 fanout2564 (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(net2564));
 sg13g2_buf_8 fanout2565 (.A(net5297),
    .X(net2565));
 sg13g2_buf_8 fanout2566 (.A(net5354),
    .X(net2566));
 sg13g2_buf_8 fanout2567 (.A(net5356),
    .X(net2567));
 sg13g2_buf_8 fanout2568 (.A(net5296),
    .X(net2568));
 sg13g2_buf_8 fanout2569 (.A(net5175),
    .X(net2569));
 sg13g2_buf_8 fanout2570 (.A(net5290),
    .X(net2570));
 sg13g2_buf_1 fanout2571 (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .X(net2571));
 sg13g2_buf_8 fanout2572 (.A(net5331),
    .X(net2572));
 sg13g2_buf_8 fanout2573 (.A(net5374),
    .X(net2573));
 sg13g2_buf_8 fanout2574 (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(net2574));
 sg13g2_buf_1 fanout2575 (.A(net5370),
    .X(net2575));
 sg13g2_buf_8 fanout2576 (.A(net4758),
    .X(net2576));
 sg13g2_buf_8 fanout2577 (.A(net5376),
    .X(net2577));
 sg13g2_buf_8 fanout2578 (.A(net4736),
    .X(net2578));
 sg13g2_buf_8 fanout2579 (.A(net5340),
    .X(net2579));
 sg13g2_buf_8 fanout2580 (.A(net5323),
    .X(net2580));
 sg13g2_buf_8 fanout2581 (.A(net5314),
    .X(net2581));
 sg13g2_buf_8 fanout2582 (.A(net5334),
    .X(net2582));
 sg13g2_buf_8 fanout2583 (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .X(net2583));
 sg13g2_buf_8 fanout2584 (.A(net4995),
    .X(net2584));
 sg13g2_buf_8 fanout2585 (.A(net4997),
    .X(net2585));
 sg13g2_buf_8 fanout2586 (.A(net4689),
    .X(net2586));
 sg13g2_buf_8 fanout2587 (.A(net4791),
    .X(net2587));
 sg13g2_buf_8 fanout2588 (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .X(net2588));
 sg13g2_buf_8 fanout2589 (.A(net5307),
    .X(net2589));
 sg13g2_buf_8 fanout2590 (.A(\i_tinyqv.cpu.instr_data_in[15] ),
    .X(net2590));
 sg13g2_buf_2 fanout2591 (.A(net5343),
    .X(net2591));
 sg13g2_buf_8 fanout2592 (.A(\i_tinyqv.cpu.instr_data_in[14] ),
    .X(net2592));
 sg13g2_buf_1 fanout2593 (.A(net5363),
    .X(net2593));
 sg13g2_buf_8 fanout2594 (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .X(net2594));
 sg13g2_buf_1 fanout2595 (.A(net5366),
    .X(net2595));
 sg13g2_buf_8 fanout2596 (.A(\i_tinyqv.cpu.instr_data_in[12] ),
    .X(net2596));
 sg13g2_buf_2 fanout2597 (.A(\i_tinyqv.cpu.instr_data_in[12] ),
    .X(net2597));
 sg13g2_buf_8 fanout2598 (.A(\i_tinyqv.cpu.instr_data_in[11] ),
    .X(net2598));
 sg13g2_buf_8 fanout2599 (.A(net5272),
    .X(net2599));
 sg13g2_buf_8 fanout2600 (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .X(net2600));
 sg13g2_buf_8 fanout2601 (.A(net5306),
    .X(net2601));
 sg13g2_buf_8 fanout2602 (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .X(net2602));
 sg13g2_buf_8 fanout2603 (.A(net5321),
    .X(net2603));
 sg13g2_buf_8 fanout2604 (.A(net5286),
    .X(net2604));
 sg13g2_buf_2 fanout2605 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(net2605));
 sg13g2_buf_8 fanout2606 (.A(net5327),
    .X(net2606));
 sg13g2_buf_8 fanout2607 (.A(net2608),
    .X(net2607));
 sg13g2_buf_8 fanout2608 (.A(net5361),
    .X(net2608));
 sg13g2_buf_8 fanout2609 (.A(net2610),
    .X(net2609));
 sg13g2_buf_8 fanout2610 (.A(net5282),
    .X(net2610));
 sg13g2_buf_8 fanout2611 (.A(net4859),
    .X(net2611));
 sg13g2_buf_8 fanout2612 (.A(net5333),
    .X(net2612));
 sg13g2_buf_8 fanout2613 (.A(net2614),
    .X(net2613));
 sg13g2_buf_8 fanout2614 (.A(net5310),
    .X(net2614));
 sg13g2_buf_8 fanout2615 (.A(net2617),
    .X(net2615));
 sg13g2_buf_8 fanout2616 (.A(net2617),
    .X(net2616));
 sg13g2_buf_8 fanout2617 (.A(net2618),
    .X(net2617));
 sg13g2_buf_8 fanout2618 (.A(net2619),
    .X(net2618));
 sg13g2_buf_8 fanout2619 (.A(net2620),
    .X(net2619));
 sg13g2_buf_2 fanout2620 (.A(net2674),
    .X(net2620));
 sg13g2_buf_8 fanout2621 (.A(net2625),
    .X(net2621));
 sg13g2_buf_1 fanout2622 (.A(net2623),
    .X(net2622));
 sg13g2_buf_8 fanout2623 (.A(net2625),
    .X(net2623));
 sg13g2_buf_8 fanout2624 (.A(net2625),
    .X(net2624));
 sg13g2_buf_8 fanout2625 (.A(net2674),
    .X(net2625));
 sg13g2_buf_8 fanout2626 (.A(net2629),
    .X(net2626));
 sg13g2_buf_8 fanout2627 (.A(net2628),
    .X(net2627));
 sg13g2_buf_8 fanout2628 (.A(net2629),
    .X(net2628));
 sg13g2_buf_8 fanout2629 (.A(net2630),
    .X(net2629));
 sg13g2_buf_8 fanout2630 (.A(net2634),
    .X(net2630));
 sg13g2_buf_8 fanout2631 (.A(net2633),
    .X(net2631));
 sg13g2_buf_2 fanout2632 (.A(net2633),
    .X(net2632));
 sg13g2_buf_8 fanout2633 (.A(net2634),
    .X(net2633));
 sg13g2_buf_8 fanout2634 (.A(net2674),
    .X(net2634));
 sg13g2_buf_8 fanout2635 (.A(net2650),
    .X(net2635));
 sg13g2_buf_8 fanout2636 (.A(net2650),
    .X(net2636));
 sg13g2_buf_8 fanout2637 (.A(net2639),
    .X(net2637));
 sg13g2_buf_8 fanout2638 (.A(net2639),
    .X(net2638));
 sg13g2_buf_8 fanout2639 (.A(net2650),
    .X(net2639));
 sg13g2_buf_8 fanout2640 (.A(net2641),
    .X(net2640));
 sg13g2_buf_8 fanout2641 (.A(net2642),
    .X(net2641));
 sg13g2_buf_8 fanout2642 (.A(net2650),
    .X(net2642));
 sg13g2_buf_8 fanout2643 (.A(net2645),
    .X(net2643));
 sg13g2_buf_8 fanout2644 (.A(net2645),
    .X(net2644));
 sg13g2_buf_8 fanout2645 (.A(net2649),
    .X(net2645));
 sg13g2_buf_8 fanout2646 (.A(net2648),
    .X(net2646));
 sg13g2_buf_1 fanout2647 (.A(net2648),
    .X(net2647));
 sg13g2_buf_8 fanout2648 (.A(net2649),
    .X(net2648));
 sg13g2_buf_2 fanout2649 (.A(net2650),
    .X(net2649));
 sg13g2_buf_8 fanout2650 (.A(net2674),
    .X(net2650));
 sg13g2_buf_8 fanout2651 (.A(net2654),
    .X(net2651));
 sg13g2_buf_1 fanout2652 (.A(net2654),
    .X(net2652));
 sg13g2_buf_8 fanout2653 (.A(net2654),
    .X(net2653));
 sg13g2_buf_2 fanout2654 (.A(net2659),
    .X(net2654));
 sg13g2_buf_8 fanout2655 (.A(net2656),
    .X(net2655));
 sg13g2_buf_8 fanout2656 (.A(net2659),
    .X(net2656));
 sg13g2_buf_8 fanout2657 (.A(net2658),
    .X(net2657));
 sg13g2_buf_8 fanout2658 (.A(net2659),
    .X(net2658));
 sg13g2_buf_8 fanout2659 (.A(net2669),
    .X(net2659));
 sg13g2_buf_8 fanout2660 (.A(net2664),
    .X(net2660));
 sg13g2_buf_8 fanout2661 (.A(net2664),
    .X(net2661));
 sg13g2_buf_8 fanout2662 (.A(net2664),
    .X(net2662));
 sg13g2_buf_8 fanout2663 (.A(net2664),
    .X(net2663));
 sg13g2_buf_8 fanout2664 (.A(net2669),
    .X(net2664));
 sg13g2_buf_8 fanout2665 (.A(net2666),
    .X(net2665));
 sg13g2_buf_8 fanout2666 (.A(net2669),
    .X(net2666));
 sg13g2_buf_8 fanout2667 (.A(net2668),
    .X(net2667));
 sg13g2_buf_8 fanout2668 (.A(net2669),
    .X(net2668));
 sg13g2_buf_8 fanout2669 (.A(net2674),
    .X(net2669));
 sg13g2_buf_8 fanout2670 (.A(net2671),
    .X(net2670));
 sg13g2_buf_8 fanout2671 (.A(net2672),
    .X(net2671));
 sg13g2_buf_8 fanout2672 (.A(net2673),
    .X(net2672));
 sg13g2_buf_8 fanout2673 (.A(net2674),
    .X(net2673));
 sg13g2_buf_8 fanout2674 (.A(net4215),
    .X(net2674));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_tiehi _16473__14 (.L_HI(net14));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_8 clkbuf_4_0__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sg13g2_buf_8 clkbuf_4_1__f_clk (.A(clknet_3_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sg13g2_buf_8 clkbuf_4_2__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_2__leaf_clk));
 sg13g2_buf_8 clkbuf_4_3__f_clk (.A(clknet_3_1_0_clk),
    .X(clknet_4_3__leaf_clk));
 sg13g2_buf_8 clkbuf_4_4__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_4__leaf_clk));
 sg13g2_buf_8 clkbuf_4_5__f_clk (.A(clknet_3_2_0_clk),
    .X(clknet_4_5__leaf_clk));
 sg13g2_buf_8 clkbuf_4_6__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_6__leaf_clk));
 sg13g2_buf_8 clkbuf_4_7__f_clk (.A(clknet_3_3_0_clk),
    .X(clknet_4_7__leaf_clk));
 sg13g2_buf_8 clkbuf_4_8__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_8__leaf_clk));
 sg13g2_buf_8 clkbuf_4_9__f_clk (.A(clknet_3_4_0_clk),
    .X(clknet_4_9__leaf_clk));
 sg13g2_buf_8 clkbuf_4_10__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_10__leaf_clk));
 sg13g2_buf_8 clkbuf_4_11__f_clk (.A(clknet_3_5_0_clk),
    .X(clknet_4_11__leaf_clk));
 sg13g2_buf_8 clkbuf_4_12__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_12__leaf_clk));
 sg13g2_buf_8 clkbuf_4_13__f_clk (.A(clknet_3_6_0_clk),
    .X(clknet_4_13__leaf_clk));
 sg13g2_buf_8 clkbuf_4_14__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_14__leaf_clk));
 sg13g2_buf_8 clkbuf_4_15__f_clk (.A(clknet_3_7_0_clk),
    .X(clknet_4_15__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_4_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_4_9__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_leaf_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_0_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_1_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_2_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_3_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_4_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_5_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_6_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_7_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_8_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_9_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_10_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_11_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_12_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_13_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_14_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_15_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_16_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_17_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_18_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_19_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_20_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_21_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_22_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_23_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_24_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_25_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_26_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_27_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_28_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_29_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_30_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_31_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_32_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_33_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_34_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_35_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_36_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_37_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_38_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_39_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_40_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_41_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_42_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_43_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_44_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_45_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_46_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_47_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_48_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_49_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_50_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_51_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_52_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_53_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_54_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_55_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_56_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_57_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_58_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_59_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_60_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_61_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_62_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_63_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_64_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_65_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_66_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_66_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_67_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_67_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_68_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_68_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_69_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_69_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_70_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_70_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_71_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_71_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_72_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_72_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_73_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_73_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_74_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_74_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_75_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_75_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_76_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_76_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_77_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_77_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_78_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_78_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_79_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_79_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_80_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_80_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_81_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_81_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_82_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_82_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_83_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_83_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_84_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_84_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_85_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_85_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_86_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_86_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_87_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_87_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_88_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_88_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_89_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_89_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_90_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_90_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_91_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_91_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_92_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_92_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_93_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_93_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_94_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_94_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_95_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_95_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_96_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_96_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_97_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_97_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_98_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_98_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_99_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_99_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_100_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_100_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_101_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_101_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_102_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_102_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_103_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_103_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_104_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_104_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_105_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_105_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_106_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_106_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_107_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_107_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_108_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_108_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_109_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_109_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_110_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_110_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_111_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_111_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_112_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_112_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_113_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_113_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_114_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_114_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_115_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_115_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_116_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_116_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_117_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_117_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_118_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_118_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_119_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_119_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_120_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_120_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_121_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_121_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_122_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_122_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_123_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_123_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_124_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_124_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_125_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_125_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_126_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_126_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_127_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_127_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_128_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_128_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_129_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_129_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_130_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_130_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_131_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_131_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_132_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_132_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_133_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_133_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_134_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_134_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_135_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_135_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_136_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_136_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_137_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_137_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_138_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_138_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_139_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_139_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_140_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_140_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_141_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_141_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_142_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_142_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_143_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_143_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_144_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_144_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_145_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_145_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_146_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_146_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_147_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_147_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_148_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_148_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_149_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_149_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_150_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_150_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_151_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_151_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_152_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_152_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_153_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_153_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_154_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_154_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_155_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_155_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_156_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_156_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_157_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_157_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_158_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_158_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_159_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_159_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_160_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_160_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_161_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_161_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_162_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_162_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_163_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_163_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_164_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_164_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_165_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_165_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_166_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_166_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_167_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_167_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_168_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_168_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_169_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_169_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_170_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_170_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_171_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_171_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_172_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_172_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_173_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_173_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_174_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_174_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_175_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_175_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_176_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_176_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_177_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_177_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_178_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_178_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_179_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_179_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_180_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_180_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_181_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_181_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_182_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_182_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_183_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_183_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_184_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_184_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_185_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_185_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_186_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_186_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_187_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_187_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_188_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_188_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_189_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_189_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_190_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_190_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_191_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_191_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_192_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_192_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_193_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_193_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_194_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_194_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_195_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_195_clk_regs));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_5_0__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_1__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_2__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_3__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_4__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_5__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_6__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_7__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_8__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_9__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_10__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_11__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_12__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_13__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_14__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_15__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_16__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_17__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_18__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_19__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_20__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_21__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_22__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_23__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_24__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_25__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_26__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_27__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_28__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_29__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_30__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_31__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_8 clkload4 (.A(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_8 clkload5 (.A(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_8 clkload6 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkload7 (.A(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkload8 (.A(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_8 clkload9 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkload10 (.A(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_8 clkload11 (.A(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_8 clkload12 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkload13 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkload14 (.A(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_8 clkload15 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_195_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold102 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold104 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold165 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold212 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold214 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold218 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold256 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold262 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold266 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold268 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold270 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold273 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold281 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold283 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold285 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold287 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold293 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold295 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold298 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold302 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold306 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold308 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold309 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold310 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold312 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold314 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold317 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold318 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold319 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold320 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold321 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold322 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold323 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold324 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold325 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold326 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold327 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold328 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold329 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold330 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold331 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold332 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold333 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold334 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold335 (.A(\i_i2c_peri.i_i2c.sda_i ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold336 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold337 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold338 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold339 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold340 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold341 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold342 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold343 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold344 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold345 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold346 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold347 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold348 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold349 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold350 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold351 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold352 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold353 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold354 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold355 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold356 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold357 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold358 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold359 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold360 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold361 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold362 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold363 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold364 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold365 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold366 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold367 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold368 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold369 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold370 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold371 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold372 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold373 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold374 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold375 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold376 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold377 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold378 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold379 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold380 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold381 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold382 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold383 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold384 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold385 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold386 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold387 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold388 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold389 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold390 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold391 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold392 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold393 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold394 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold395 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold396 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold397 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold398 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold399 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold400 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold401 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold402 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold403 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold404 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold405 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold406 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold407 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold408 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold409 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold410 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold411 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold412 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold414 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold415 (.A(\i_i2c_peri.i_i2c.sda_i_reg ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold416 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold417 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold418 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold419 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold420 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold421 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold423 (.A(\reset_hold_counter[5] ),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold424 (.A(combined_rst_n),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold425 (.A(\i_uart_rx.rxd_reg[1] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold426 (.A(\i_uart_rx.cycle_counter[0] ),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold427 (.A(\i_i2c_peri.i_i2c.delay_sda_reg ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold428 (.A(_01213_),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold429 (.A(\pps_sync[0] ),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold430 (.A(\us_divider[0] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold431 (.A(\pps_sync[1] ),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold432 (.A(\session_ms_div[9] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold433 (.A(_00388_),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold434 (.A(\session_ms_div[2] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold435 (.A(_00381_),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold436 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[6] ),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold437 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[3] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold438 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[0] ),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[5] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold440 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[0] ),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold441 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[0] ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold442 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[6] ),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold443 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[7] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold444 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[2] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold445 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[5] ),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold446 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[0] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[1] ),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold448 (.A(\reset_hold_counter[0] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold449 (.A(_00451_),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold450 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[2] ),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold451 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[1] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold452 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[0] ),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold453 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[7] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold454 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[1] ),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold455 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[2] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold456 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[1] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold457 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[5] ),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold458 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[7] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold459 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[5] ),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold460 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[0] ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold461 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[7] ),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold462 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[7] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold463 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[6] ),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold464 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[3] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold465 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[4] ),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold466 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[6] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold467 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[3] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold468 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[0] ),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold469 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[6] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold470 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[5] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold471 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[6] ),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold472 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[2] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold473 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[5] ),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold474 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[1] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold475 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[5] ),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold476 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[1] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold477 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[7] ),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold478 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[3] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold479 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[5] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold480 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[4] ),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold481 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[2] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold482 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[2] ),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold483 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[3] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold484 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[4] ),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold485 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[0] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold486 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[2] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold487 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[1] ),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold488 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[2] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold489 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[4] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold490 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[4] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold491 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[1] ),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold492 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[4] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold493 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[3] ),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold494 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[7] ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold495 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[2] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold496 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[2] ),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold497 (.A(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold498 (.A(_01252_),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold499 (.A(\i_crc16.bit_cnt[0] ),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold500 (.A(_00800_),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold501 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[4] ),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold502 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[0] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold503 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[3] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold504 (.A(\i_tinyqv.mem.qspi_data_buf[24] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold505 (.A(_00511_),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold506 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[7] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold507 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[6] ),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold508 (.A(\i_latch_mem.data_out[24] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold509 (.A(_00028_),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold510 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[2] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold511 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[0] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold512 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[2] ),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold513 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[2] ),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold514 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[1] ),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold515 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[3] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold516 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[6] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold517 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[5] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold518 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[4] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold519 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[5] ),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold520 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[6] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold521 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[6] ),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold522 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[7] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold523 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[3] ),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold524 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[6] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold525 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[1] ),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold526 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[4] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold527 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[7] ),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold528 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[1] ),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold529 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[6] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold530 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[5] ),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold531 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[5] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold532 (.A(\session_ms_div[7] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00386_),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold534 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[1] ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold535 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[5] ),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold536 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[3] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold537 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[3] ),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold538 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[0] ),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold539 (.A(\i_rtc.us_count[2] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold540 (.A(_00839_),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold541 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[0] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold542 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[7] ),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold543 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[6] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold544 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[7] ),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold545 (.A(\i_seal.sensor_id_reg[0] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold546 (.A(_01048_),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold547 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[4] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold548 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[1] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold549 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[4] ),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold550 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[5] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold551 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[7] ),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold552 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[5] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold553 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[2] ),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold554 (.A(\i_latch_mem.genblk1[0].l_ram.data_out[5] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold555 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[4] ),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold556 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[3] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold557 (.A(\i_seal.mono_count[29] ),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold558 (.A(_01013_),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold559 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[6] ),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold560 (.A(\i_spi.end_txn_reg ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold561 (.A(_01378_),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold562 (.A(\i_seal.sealed_crc[11] ),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold563 (.A(_00906_),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold564 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[3] ),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold565 (.A(\i_latch_mem.genblk1[27].l_ram.data_out[7] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[0] ),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold567 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[4] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold568 (.A(\i_seal.mono_count[26] ),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold569 (.A(_06550_),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold570 (.A(_01010_),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold571 (.A(\i_latch_mem.genblk1[9].l_ram.data_out[4] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold572 (.A(\i_seal.sealed_crc[8] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold573 (.A(_00903_),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold574 (.A(\i_tinyqv.cpu.i_core.mie[3] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold575 (.A(_01654_),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold576 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[2] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold577 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[6] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold578 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[2] ),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold579 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold580 (.A(_00553_),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold581 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[1] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold582 (.A(\i_seal.sealed_crc[10] ),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold583 (.A(_00905_),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold584 (.A(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold585 (.A(_00797_),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold586 (.A(\i_seal.sealed_crc[15] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold587 (.A(_00910_),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold588 (.A(\pps_count[12] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold589 (.A(_00409_),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold590 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[1] ),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold591 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[0] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold592 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[2] ),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold593 (.A(\us_divider[1] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold594 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[6] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_tinyqv.cpu.i_core.mie[4] ),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold596 (.A(_01653_),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[7] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold598 (.A(\i_latch_mem.genblk1[19].l_ram.data_out[3] ),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold599 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[1] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold600 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[3] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold601 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[6] ),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold602 (.A(\i_latch_mem.genblk1[8].l_ram.data_out[5] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold603 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[0] ),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold604 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[0] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold605 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[3] ),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold606 (.A(\i_seal.sealed_crc[14] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold607 (.A(_00909_),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold608 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[0] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold609 (.A(\i_uart_tx.data_to_send[7] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold610 (.A(_01337_),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold611 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[4] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold612 (.A(\i_i2c_peri.sda_sync[0] ),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold613 (.A(\i_latch_mem.genblk1[7].l_ram.data_out[0] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold614 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[1] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold615 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[0] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold616 (.A(\i_latch_mem.genblk1[2].l_ram.data_out[5] ),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold617 (.A(\i_latch_mem.genblk1[16].l_ram.data_out[3] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold618 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[2] ),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold619 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[4] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold620 (.A(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold621 (.A(_06013_),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold622 (.A(_00781_),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold623 (.A(\i_rtc.us_count[3] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold624 (.A(_06233_),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold625 (.A(\i_rtc.us_count[17] ),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold626 (.A(_00854_),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold627 (.A(\i_i2c_peri.i_i2c.data_reg[7] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold628 (.A(_01643_),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold629 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[2] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold630 (.A(\i_seal.sensor_id_reg[2] ),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold631 (.A(_01050_),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold632 (.A(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold633 (.A(_00758_),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold634 (.A(\i_seal.sensor_id_reg[5] ),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold635 (.A(_01053_),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold636 (.A(\i_latch_mem.genblk1[1].l_ram.data_out[7] ),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold637 (.A(\i_spi.clock_count[1] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold638 (.A(_01669_),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold639 (.A(_01380_),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold640 (.A(\i_latch_mem.genblk1[24].l_ram.data_out[0] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold641 (.A(\i_latch_mem.data_out[29] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold642 (.A(_00033_),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold643 (.A(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold644 (.A(_00786_),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold645 (.A(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold646 (.A(_00783_),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold647 (.A(\i_spi.data[1] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold648 (.A(_01177_),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold649 (.A(\i_i2c_peri.i_i2c.last_sda_i_reg ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold650 (.A(_06891_),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold651 (.A(_01215_),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold652 (.A(\i_tinyqv.mem.qspi_data_buf[31] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold653 (.A(_00518_),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold654 (.A(\i_tinyqv.cpu.instr_data[2][3] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold655 (.A(_01187_),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold656 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[6] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold657 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[1] ),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold658 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[4] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold659 (.A(\i_latch_mem.data_out[28] ),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold660 (.A(_00032_),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold661 (.A(\i_spi.data[4] ),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold662 (.A(_01180_),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold663 (.A(\i_seal.sensor_id_reg[3] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold664 (.A(_01051_),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold665 (.A(\i_seal.sensor_id_reg[4] ),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold666 (.A(_01052_),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold667 (.A(\i_spi.data[2] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold668 (.A(\i_i2c_peri.i_i2c.mode_write_multiple_reg ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold669 (.A(_01242_),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold670 (.A(debug_data_continue),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold671 (.A(_00480_),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold672 (.A(\i_seal.mono_count[9] ),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold673 (.A(_01025_),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold674 (.A(\i_latch_mem.genblk1[25].l_ram.data_out[4] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold675 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[6] ),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold676 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[2] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold677 (.A(\i_spi.data[5] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold678 (.A(_01181_),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold679 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[1] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold680 (.A(\i_latch_mem.data_out[30] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold681 (.A(_00035_),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold682 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[4] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold683 (.A(\i_seal.mono_count[20] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold684 (.A(_01036_),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold685 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[0] ),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold686 (.A(\i_seal.sealed_crc[12] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold687 (.A(_00907_),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold688 (.A(\i_spi.data[3] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold689 (.A(_01179_),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold690 (.A(\i_latch_mem.genblk1[3].l_ram.data_out[7] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold691 (.A(\i_seal.mono_count[24] ),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold692 (.A(_01040_),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold693 (.A(\i_seal.sensor_id_reg[1] ),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold694 (.A(_01049_),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold695 (.A(\i_seal.sealed_crc[9] ),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold696 (.A(_00904_),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold697 (.A(\i_tinyqv.cpu.instr_data[1][0] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold698 (.A(_00556_),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold699 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[7] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold700 (.A(\i_tinyqv.cpu.i_core.mepc[4] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold701 (.A(_01113_),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold702 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[1] ),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold703 (.A(\i_seal.mono_count[30] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold704 (.A(_06557_),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold705 (.A(_01014_),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold706 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[6] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold707 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[4] ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold708 (.A(\i_latch_mem.data_out[19] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold709 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[4] ),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold710 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[2] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold711 (.A(\i_tinyqv.cpu.instr_data[2][8] ),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold712 (.A(_01192_),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold713 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[1] ),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold714 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[3] ),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold715 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[3] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold716 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[7] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold717 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[0] ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold718 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[3] ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold719 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[5] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold720 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[5] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold721 (.A(\i_latch_mem.data_out[15] ),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold722 (.A(\us_divider[2] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold723 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[7] ),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold724 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[7] ),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold725 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[3] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold726 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[5] ),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold727 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[0] ),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold728 (.A(\session_ms_div[4] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold729 (.A(_04346_),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold730 (.A(_00383_),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold731 (.A(\i_seal.mono_count[6] ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold732 (.A(_01022_),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold733 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[6] ),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold734 (.A(\i_spi.data[7] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold735 (.A(_01183_),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold736 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[5] ),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold737 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold738 (.A(_04892_),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold739 (.A(_00541_),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold740 (.A(\i_i2c_peri.i_i2c.delay_reg[13] ),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold741 (.A(_06971_),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold742 (.A(\i_tinyqv.mem.qspi_data_buf[8] ),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold743 (.A(_00495_),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold744 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[5] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold745 (.A(\i_seal.mono_count[10] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold746 (.A(_01026_),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold747 (.A(\i_tinyqv.cpu.instr_data[3][3] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold748 (.A(_01254_),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold749 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[2] ),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold750 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[7] ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold751 (.A(\i_latch_mem.genblk1[26].l_ram.data_out[4] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold752 (.A(\i_latch_mem.data_out[1] ),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold753 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[5] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold754 (.A(\i_latch_mem.data_out[18] ),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold755 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[3] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold756 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[3] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold757 (.A(\i_latch_mem.genblk1[10].l_ram.data_out[1] ),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold758 (.A(\i_tinyqv.mem.qspi_data_buf[10] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold759 (.A(_00497_),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold760 (.A(\i_tinyqv.cpu.instr_data[1][1] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold761 (.A(_00557_),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold762 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold763 (.A(_00554_),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold764 (.A(\session_ms_div[1] ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold765 (.A(_04333_),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold766 (.A(_00380_),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold767 (.A(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold768 (.A(_00784_),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold769 (.A(\i_i2c_peri.cmd_addr_reg[0] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold770 (.A(_01294_),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold771 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[6] ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold772 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[6] ),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold773 (.A(\session_ms_div[8] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold774 (.A(_04357_),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold775 (.A(\i_latch_mem.data_out[17] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold776 (.A(\i_seal.mono_count[19] ),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold777 (.A(_06539_),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold778 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[6] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold779 (.A(\i_latch_mem.data_out[9] ),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold780 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[6] ),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold781 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[2] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold782 (.A(\i_latch_mem.data_out[31] ),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold783 (.A(\i_seal.sealed_mono[12] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold784 (.A(_00923_),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold785 (.A(\i_rtc.us_count[1] ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold786 (.A(_06228_),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold787 (.A(_00838_),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold788 (.A(\i_i2c_peri.i_i2c.addr_reg[0] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold789 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[2] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold790 (.A(\i_tinyqv.cpu.instr_data[0][0] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold791 (.A(_01376_),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold792 (.A(\i_tinyqv.cpu.i_core.mcause[3] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold793 (.A(_00458_),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold794 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[4] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold795 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[3] ),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold796 (.A(\i_latch_mem.genblk1[17].l_ram.data_out[5] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold797 (.A(\i_seal.session_ctr_in[4] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold798 (.A(_04367_),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold799 (.A(_00393_),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold800 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[0] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold801 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[1] ),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold802 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[6] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold803 (.A(\i_seal.value_reg[8] ),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold804 (.A(_00951_),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold805 (.A(\i_latch_mem.data_out[7] ),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold806 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[4] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold807 (.A(\i_seal.session_ctr_in[1] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold808 (.A(_00977_),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold809 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[1] ),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold810 (.A(\i_latch_mem.genblk1[6].l_ram.data_out[5] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold811 (.A(\i_tinyqv.mem.data_from_read[16] ),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold812 (.A(_04758_),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold813 (.A(_00503_),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold814 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[7] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold815 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[0] ),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold816 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[2] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold817 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[3] ),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold818 (.A(\i_i2c_peri.cmd_addr_reg[6] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold819 (.A(_01300_),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold820 (.A(\i_tinyqv.cpu.instr_data[3][8] ),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold821 (.A(_01259_),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold822 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[5] ),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold823 (.A(\i_i2c_peri.i_i2c.addr_reg[6] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold824 (.A(\i_latch_mem.data_out[2] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold825 (.A(\i_tinyqv.cpu.instr_data[0][1] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold826 (.A(_01377_),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold827 (.A(\i_latch_mem.data_out[25] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold828 (.A(\i_latch_mem.data_out[27] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold829 (.A(\i_uart_rx.cycle_counter[3] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold830 (.A(_07205_),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold831 (.A(_01362_),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold832 (.A(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold833 (.A(_00792_),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold834 (.A(\i_latch_mem.data_out[23] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold835 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[5] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold836 (.A(\i_uart_rx.cycle_counter[6] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold837 (.A(_07210_),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold838 (.A(_01365_),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold839 (.A(\i_latch_mem.genblk1[11].l_ram.data_out[7] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold840 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[4] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold841 (.A(\i_tinyqv.mem.qspi_data_buf[11] ),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold842 (.A(_00498_),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold843 (.A(\i_seal.cur_mono[25] ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold844 (.A(_00936_),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold845 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[3] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold846 (.A(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold847 (.A(_00779_),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold848 (.A(\session_ms_div[5] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold849 (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[7] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold850 (.A(_01212_),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold851 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[5] ),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold852 (.A(\i_latch_mem.data_out[26] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold853 (.A(\i_seal.mono_count[21] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold854 (.A(_01037_),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold855 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[4] ),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold856 (.A(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold857 (.A(_00777_),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold858 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[4] ),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold859 (.A(\i_tinyqv.cpu.instr_data[3][0] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold860 (.A(_01200_),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold861 (.A(\i_tinyqv.cpu.imm[27] ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold862 (.A(\i_seal.cur_mono[28] ),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold863 (.A(_00939_),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold864 (.A(\i_seal.cur_mono[30] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold865 (.A(_06591_),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold866 (.A(\i_tinyqv.mem.qspi_data_buf[12] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold867 (.A(_00499_),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold868 (.A(\i_spi.data[6] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold869 (.A(_01182_),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold870 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[2] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold871 (.A(\i_latch_mem.data_out[10] ),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold872 (.A(_00013_),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold873 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[0] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold874 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[2] ),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold875 (.A(\pps_count[13] ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold876 (.A(_04399_),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold877 (.A(\i_latch_mem.genblk1[28].l_ram.data_out[7] ),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold878 (.A(\i_tinyqv.cpu.load_started ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold879 (.A(_00656_),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold880 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[2] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold881 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[0] ),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold882 (.A(\i_seal.mono_count[14] ),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold883 (.A(_01030_),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold884 (.A(\i_tinyqv.cpu.i_core.load_done ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold885 (.A(_00751_),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold886 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[7] ),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold887 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[1] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold888 (.A(\i_seal.mono_count[15] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold889 (.A(_01031_),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold890 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[5] ),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold891 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[1] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold892 (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold893 (.A(\i_latch_mem.data_out[8] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold894 (.A(\i_i2c_peri.i_i2c.delay_reg[14] ),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold895 (.A(_06976_),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold896 (.A(\i_tinyqv.mem.qspi_data_buf[13] ),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold897 (.A(_00500_),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold898 (.A(\i_tinyqv.mem.qspi_data_buf[15] ),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold899 (.A(_00502_),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold900 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[0] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold901 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[1] ),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold902 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[3] ),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold903 (.A(\i_seal.session_ctr_in[5] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold904 (.A(_00981_),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold905 (.A(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold906 (.A(_00790_),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold907 (.A(\i_seal.mono_count[5] ),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold908 (.A(_06516_),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold909 (.A(_00990_),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold910 (.A(\i_seal.mono_count[16] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold911 (.A(_01032_),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold912 (.A(\i_latch_mem.data_out[3] ),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold913 (.A(\i_seal.mono_count[12] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold914 (.A(_06526_),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold915 (.A(_00996_),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold916 (.A(\i_latch_mem.genblk1[18].l_ram.data_out[2] ),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold917 (.A(\i_seal.session_ctr_in[0] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold918 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[0] ),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold919 (.A(\i_seal.mono_count[13] ),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold920 (.A(_06529_),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold921 (.A(\i_latch_mem.genblk1[4].l_ram.data_out[3] ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold922 (.A(\gpio_out[1] ),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold923 (.A(_00371_),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold924 (.A(\i_uart_tx.cycle_counter[2] ),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold925 (.A(_07167_),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold926 (.A(_01340_),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold927 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[7] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold928 (.A(\i_tinyqv.cpu.instr_data[2][1] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold929 (.A(_00799_),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold930 (.A(\i_seal.sensor_id_reg[6] ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold931 (.A(_01054_),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold932 (.A(\i_latch_mem.data_out[16] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold933 (.A(_00019_),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold934 (.A(\i_spi.read_latency ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold935 (.A(\i_seal.mono_count[27] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold936 (.A(_01043_),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold937 (.A(\i_seal.mono_count[28] ),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold938 (.A(\i_latch_mem.data_out[0] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold939 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[7] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold940 (.A(\i_seal.sealed_mono[11] ),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold941 (.A(_00922_),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold942 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[1] ),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold943 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[5] ),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold944 (.A(\i_seal.value_reg[7] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold945 (.A(_00950_),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold946 (.A(\i_seal.session_ctr_in[6] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold947 (.A(_00982_),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold948 (.A(\i_latch_mem.data_out[11] ),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold949 (.A(\i_seal.mono_count[8] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold950 (.A(_06519_),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold951 (.A(_00992_),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold952 (.A(\i_latch_mem.genblk1[5].l_ram.data_out[7] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold953 (.A(\pps_count[15] ),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold954 (.A(_00412_),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold955 (.A(\i_seal.mono_count[31] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold956 (.A(_01015_),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold957 (.A(\i_spi.clock_divider[2] ),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold958 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[5] ),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold959 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[1] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold960 (.A(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold961 (.A(_00795_),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold962 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold963 (.A(_00721_),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold964 (.A(\i_seal.sealed_mono[15] ),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold965 (.A(_00926_),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold966 (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[2] ),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold967 (.A(_01207_),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold968 (.A(\i_seal.value_reg[6] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold969 (.A(_00949_),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold970 (.A(\i_tinyqv.cpu.i_core.mepc[22] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold971 (.A(_01131_),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold972 (.A(\i_seal.mono_count[3] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold973 (.A(_01019_),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold974 (.A(\i_seal.value_reg[4] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold975 (.A(_00947_),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold976 (.A(\i_seal.crc_byte[0] ),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold977 (.A(_01091_),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold978 (.A(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold979 (.A(_00761_),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold980 (.A(\i_seal.value_reg[17] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold981 (.A(_00960_),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold982 (.A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold983 (.A(_00770_),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold984 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[4] ),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold985 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[2] ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold986 (.A(\i_seal.crc_byte[7] ),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold987 (.A(_01098_),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold988 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[1] ),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold989 (.A(\i_seal.mono_count[18] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold990 (.A(_06536_),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold991 (.A(_01002_),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold992 (.A(\i2c_data_out[5] ),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold993 (.A(_01318_),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold994 (.A(\i_tinyqv.cpu.instr_data[2][0] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold995 (.A(_00798_),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold996 (.A(\i_latch_mem.data_out[5] ),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold997 (.A(\i_seal.mono_count[25] ),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold998 (.A(\i_tinyqv.mem.qspi_data_buf[14] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold999 (.A(_00501_),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\i_seal.cur_mono[26] ),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1001 (.A(_00937_),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\i_tinyqv.cpu.instr_data[0][3] ),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1003 (.A(_01134_),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\i_seal.cur_mono[8] ),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1005 (.A(\i_latch_mem.genblk1[15].l_ram.data_out[6] ),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\i_i2c_peri.cmd_stop_reg ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1007 (.A(_01216_),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\i_seal.session_ctr_in[7] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1009 (.A(_00396_),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1010 (.A(\i_seal.sealed_sid[7] ),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1011 (.A(_06505_),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1012 (.A(_00983_),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1013 (.A(\i_uart_tx.cycle_counter[7] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_07177_),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1015 (.A(_01345_),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1016 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[4] ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\i_seal.mono_count[23] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1018 (.A(_01039_),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[4] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1020 (.A(\i_latch_mem.genblk1[12].l_ram.data_out[2] ),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\i_tinyqv.cpu.i_core.mepc[21] ),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1022 (.A(_01130_),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1023 (.A(\i_seal.value_reg[16] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1024 (.A(_00959_),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1025 (.A(\i_seal.value_reg[20] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1026 (.A(_00963_),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1027 (.A(\pps_count[6] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1028 (.A(_04387_),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_00403_),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1030 (.A(\i_rtc.us_count[8] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1031 (.A(_06258_),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_00845_),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1033 (.A(\i_seal.cur_mono[18] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\i_seal.value_reg[18] ),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1035 (.A(_00961_),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1036 (.A(\i_spi.clock_divider[0] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1038 (.A(\i_seal.sealed_sid[4] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\i_uart_tx.fsm_state[1] ),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1040 (.A(_01348_),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\pps_count[10] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_04394_),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1043 (.A(_00407_),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1044 (.A(\i2c_data_out[1] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1045 (.A(_01314_),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1046 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[3] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\i_seal.value_reg[14] ),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_00957_),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\i_seal.mono_count[22] ),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1050 (.A(_01038_),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\i_tinyqv.mem.qspi_write_done ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1052 (.A(_04731_),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1053 (.A(_06111_),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1054 (.A(\i_latch_mem.genblk1[23].l_ram.data_out[3] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\i_seal.sensor_id_reg[7] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1056 (.A(_01055_),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\i_seal.mono_count[17] ),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1058 (.A(_01033_),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1059 (.A(\pps_count[1] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1060 (.A(_04378_),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1061 (.A(_00398_),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1062 (.A(\i_uart_rx.bit_sample ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1063 (.A(_07219_),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1064 (.A(_01368_),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\i_seal.cur_mono[31] ),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1066 (.A(_06592_),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\i_tinyqv.cpu.instr_data[3][1] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1068 (.A(_01201_),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\i_latch_mem.genblk1[20].l_ram.data_out[3] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1070 (.A(\i_seal.mono_count[2] ),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1071 (.A(_00986_),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1072 (.A(\i_latch_mem.genblk1[31].l_ram.data_out[2] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\i_i2c_peri.cmd_pending ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1074 (.A(_01290_),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[6] ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1076 (.A(_01211_),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\i_seal.cur_mono[19] ),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\i_latch_mem.data_out[21] ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\i_tinyqv.cpu.i_core.mepc[20] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_00764_),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\i_latch_mem.data_out[14] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\i2c_data_out[3] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1083 (.A(_01316_),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[6] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1085 (.A(\i_seal.cur_mono[5] ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\i_i2c_peri.cmd_addr_reg[4] ),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_01247_),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[7] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1089 (.A(\i_seal.value_reg[28] ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1090 (.A(_00971_),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1091 (.A(\i_i2c_peri.i_i2c.delay_reg[12] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1092 (.A(_01233_),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1093 (.A(\i_latch_mem.genblk1[13].l_ram.data_out[6] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\i_rtc.us_count[4] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\i_seal.value_reg[30] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1096 (.A(_00973_),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\i_seal.cur_mono[2] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1098 (.A(_00913_),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\dio1_sync[0] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1100 (.A(\i_spi.clock_divider[1] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[0] ),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1102 (.A(\i_seal.sealed_sid[0] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1103 (.A(_06498_),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1104 (.A(_00976_),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[4] ),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1106 (.A(\i_tinyqv.mem.qspi_data_buf[28] ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1107 (.A(_00515_),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1109 (.A(_00543_),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\i_rtc.us_count[18] ),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1111 (.A(_06276_),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\i_seal.cur_mono[29] ),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\i_latch_mem.data_out[13] ),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1114 (.A(\i_tinyqv.mem.data_from_read[20] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1115 (.A(_00507_),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\i_seal.value_reg[22] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1117 (.A(_00965_),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\i_tinyqv.mem.qspi_data_buf[27] ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1119 (.A(_00514_),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\i_latch_mem.genblk1[30].l_ram.data_out[1] ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\i_tinyqv.mem.qspi_data_buf[9] ),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1122 (.A(_00496_),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1124 (.A(_00772_),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\i_latch_mem.genblk1[22].l_ram.data_out[6] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[5] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1127 (.A(_01210_),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1128 (.A(\i_seal.cur_mono[1] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1129 (.A(_00912_),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1130 (.A(\i2c_data_out[4] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1131 (.A(_01317_),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1132 (.A(\i_seal.cur_mono[4] ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1133 (.A(_00915_),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1134 (.A(\addr[10] ),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1135 (.A(_01163_),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\i_seal.value_reg[15] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1137 (.A(_00958_),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\i_seal.mono_count[1] ),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1139 (.A(\i_latch_mem.data_out[22] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\i_tinyqv.cpu.i_core.mie[1] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1141 (.A(_01656_),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\i_seal.commit_dropped ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1144 (.A(_00544_),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1145 (.A(\i_i2c_peri.i_i2c.addr_reg[3] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1146 (.A(_01246_),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\us_divider[3] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1148 (.A(\i_tinyqv.mem.qspi_data_buf[30] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1149 (.A(_00517_),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\i_wdt.wdt_reset ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1151 (.A(_00460_),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\i_seal.value_reg[23] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1153 (.A(_00966_),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold1155 (.A(_05874_),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\i_seal.session_ctr_in[3] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold1157 (.A(_00979_),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold1158 (.A(\i_seal.crc_byte[3] ),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold1159 (.A(_01094_),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold1160 (.A(\i_seal.cur_mono[27] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold1161 (.A(_00938_),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold1162 (.A(\i_latch_mem.data_out[20] ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\i_tinyqv.mem.qspi_data_buf[26] ),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold1164 (.A(_00513_),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\i_seal.cur_mono[17] ),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold1166 (.A(_00928_),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold1167 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[1] ),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[7] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold1169 (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold1170 (.A(_00762_),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\i_tinyqv.mem.qspi_data_buf[29] ),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_00516_),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\i_seal.value_reg[21] ),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold1174 (.A(_00964_),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[6] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold1176 (.A(\i_tinyqv.mem.qspi_data_buf[25] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold1177 (.A(_00512_),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\i_seal.sealed_mono[5] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold1179 (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[0] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold1180 (.A(_01205_),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold1181 (.A(\i_tinyqv.cpu.instr_data[1][8] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold1182 (.A(_00467_),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold1183 (.A(\i_i2c_peri.i_i2c.last_reg ),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold1184 (.A(_01219_),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold1185 (.A(\i_tinyqv.mem.data_from_read[21] ),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold1186 (.A(_00508_),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold1187 (.A(\data_to_write[8] ),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\i_crc16.bit_cnt[3] ),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold1189 (.A(_06123_),
    .X(net4171));
 sg13g2_dlygate4sd3_1 hold1190 (.A(_00802_),
    .X(net4172));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\i_seal.cur_mono[24] ),
    .X(net4173));
 sg13g2_dlygate4sd3_1 hold1192 (.A(_00935_),
    .X(net4174));
 sg13g2_dlygate4sd3_1 hold1193 (.A(\i_tinyqv.mem.data_from_read[17] ),
    .X(net4175));
 sg13g2_dlygate4sd3_1 hold1194 (.A(_00504_),
    .X(net4176));
 sg13g2_dlygate4sd3_1 hold1195 (.A(\i_tinyqv.cpu.i_core.mie[2] ),
    .X(net4177));
 sg13g2_dlygate4sd3_1 hold1196 (.A(_01655_),
    .X(net4178));
 sg13g2_dlygate4sd3_1 hold1197 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .X(net4179));
 sg13g2_dlygate4sd3_1 hold1198 (.A(_00542_),
    .X(net4180));
 sg13g2_dlygate4sd3_1 hold1199 (.A(\i_seal.cur_mono[13] ),
    .X(net4181));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\i_i2c_peri.i_i2c.delay_reg[16] ),
    .X(net4182));
 sg13g2_dlygate4sd3_1 hold1201 (.A(_06980_),
    .X(net4183));
 sg13g2_dlygate4sd3_1 hold1202 (.A(_01237_),
    .X(net4184));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\addr[13] ),
    .X(net4185));
 sg13g2_dlygate4sd3_1 hold1204 (.A(_01166_),
    .X(net4186));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\i_seal.cur_mono[0] ),
    .X(net4187));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_00911_),
    .X(net4188));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\i_seal.value_reg[24] ),
    .X(net4189));
 sg13g2_dlygate4sd3_1 hold1208 (.A(_00967_),
    .X(net4190));
 sg13g2_dlygate4sd3_1 hold1209 (.A(\i_seal.crc_byte[1] ),
    .X(net4191));
 sg13g2_dlygate4sd3_1 hold1210 (.A(_01092_),
    .X(net4192));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\i_uart_rx.recieved_data[0] ),
    .X(net4193));
 sg13g2_dlygate4sd3_1 hold1212 (.A(_01351_),
    .X(net4194));
 sg13g2_dlygate4sd3_1 hold1213 (.A(\i_tinyqv.mem.data_from_read[22] ),
    .X(net4195));
 sg13g2_dlygate4sd3_1 hold1214 (.A(_00509_),
    .X(net4196));
 sg13g2_dlygate4sd3_1 hold1215 (.A(\i_seal.value_reg[9] ),
    .X(net4197));
 sg13g2_dlygate4sd3_1 hold1216 (.A(_00952_),
    .X(net4198));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\i_spi.bits_remaining[3] ),
    .X(net4199));
 sg13g2_dlygate4sd3_1 hold1218 (.A(_01686_),
    .X(net4200));
 sg13g2_dlygate4sd3_1 hold1219 (.A(_01387_),
    .X(net4201));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\i_seal.mono_count[0] ),
    .X(net4202));
 sg13g2_dlygate4sd3_1 hold1221 (.A(\i2c_data_out[7] ),
    .X(net4203));
 sg13g2_dlygate4sd3_1 hold1222 (.A(_01320_),
    .X(net4204));
 sg13g2_dlygate4sd3_1 hold1223 (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .X(net4205));
 sg13g2_dlygate4sd3_1 hold1224 (.A(_00763_),
    .X(net4206));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[4] ),
    .X(net4207));
 sg13g2_dlygate4sd3_1 hold1226 (.A(_01209_),
    .X(net4208));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\i_tinyqv.cpu.instr_data[0][8] ),
    .X(net4209));
 sg13g2_dlygate4sd3_1 hold1228 (.A(_01139_),
    .X(net4210));
 sg13g2_dlygate4sd3_1 hold1229 (.A(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .X(net4211));
 sg13g2_dlygate4sd3_1 hold1230 (.A(_00776_),
    .X(net4212));
 sg13g2_dlygate4sd3_1 hold1231 (.A(\i_seal.crc_byte[4] ),
    .X(net4213));
 sg13g2_dlygate4sd3_1 hold1232 (.A(_01095_),
    .X(net4214));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\i_crc16.rst_n ),
    .X(net4215));
 sg13g2_dlygate4sd3_1 hold1234 (.A(\i_rtc.us_count[12] ),
    .X(net4216));
 sg13g2_dlygate4sd3_1 hold1235 (.A(_06265_),
    .X(net4217));
 sg13g2_dlygate4sd3_1 hold1236 (.A(_00849_),
    .X(net4218));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[0] ),
    .X(net4219));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\i_latch_mem.genblk1[14].l_ram.data_out[6] ),
    .X(net4220));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\i_seal.value_reg[13] ),
    .X(net4221));
 sg13g2_dlygate4sd3_1 hold1240 (.A(_00956_),
    .X(net4222));
 sg13g2_dlygate4sd3_1 hold1241 (.A(\i_i2c_peri.cmd_addr_reg[1] ),
    .X(net4223));
 sg13g2_dlygate4sd3_1 hold1242 (.A(_01295_),
    .X(net4224));
 sg13g2_dlygate4sd3_1 hold1243 (.A(\addr[11] ),
    .X(net4225));
 sg13g2_dlygate4sd3_1 hold1244 (.A(_01164_),
    .X(net4226));
 sg13g2_dlygate4sd3_1 hold1245 (.A(\i_seal.value_reg[31] ),
    .X(net4227));
 sg13g2_dlygate4sd3_1 hold1246 (.A(_00974_),
    .X(net4228));
 sg13g2_dlygate4sd3_1 hold1247 (.A(\i_spi.bits_remaining[0] ),
    .X(net4229));
 sg13g2_dlygate4sd3_1 hold1248 (.A(_01681_),
    .X(net4230));
 sg13g2_dlygate4sd3_1 hold1249 (.A(_01384_),
    .X(net4231));
 sg13g2_dlygate4sd3_1 hold1250 (.A(\addr[7] ),
    .X(net4232));
 sg13g2_dlygate4sd3_1 hold1251 (.A(_01160_),
    .X(net4233));
 sg13g2_dlygate4sd3_1 hold1252 (.A(\addr[8] ),
    .X(net4234));
 sg13g2_dlygate4sd3_1 hold1253 (.A(_01161_),
    .X(net4235));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\i_wdt.counter[24] ),
    .X(net4236));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_06201_),
    .X(net4237));
 sg13g2_dlygate4sd3_1 hold1256 (.A(_00828_),
    .X(net4238));
 sg13g2_dlygate4sd3_1 hold1257 (.A(\i_tinyqv.mem.data_from_read[19] ),
    .X(net4239));
 sg13g2_dlygate4sd3_1 hold1258 (.A(_00506_),
    .X(net4240));
 sg13g2_dlygate4sd3_1 hold1259 (.A(\i_i2c_peri.i_i2c.addr_reg[2] ),
    .X(net4241));
 sg13g2_dlygate4sd3_1 hold1260 (.A(_01245_),
    .X(net4242));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\i_seal.crc_byte[5] ),
    .X(net4243));
 sg13g2_dlygate4sd3_1 hold1262 (.A(_01096_),
    .X(net4244));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\i_i2c_peri.i_i2c.delay_reg[7] ),
    .X(net4245));
 sg13g2_dlygate4sd3_1 hold1264 (.A(_06942_),
    .X(net4246));
 sg13g2_dlygate4sd3_1 hold1265 (.A(_01228_),
    .X(net4247));
 sg13g2_dlygate4sd3_1 hold1266 (.A(\i_i2c_peri.i_i2c.addr_reg[5] ),
    .X(net4248));
 sg13g2_dlygate4sd3_1 hold1267 (.A(_01248_),
    .X(net4249));
 sg13g2_dlygate4sd3_1 hold1268 (.A(\i_spi.spi_select ),
    .X(net4250));
 sg13g2_dlygate4sd3_1 hold1269 (.A(_01688_),
    .X(net4251));
 sg13g2_dlygate4sd3_1 hold1270 (.A(_01389_),
    .X(net4252));
 sg13g2_dlygate4sd3_1 hold1271 (.A(\i_seal.cur_mono[7] ),
    .X(net4253));
 sg13g2_dlygate4sd3_1 hold1272 (.A(_00918_),
    .X(net4254));
 sg13g2_dlygate4sd3_1 hold1273 (.A(\i_i2c_peri.i_i2c.addr_reg[1] ),
    .X(net4255));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[3] ),
    .X(net4256));
 sg13g2_dlygate4sd3_1 hold1275 (.A(\i_tinyqv.cpu.imm[29] ),
    .X(net4257));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\i_i2c_peri.cmd_addr_reg[5] ),
    .X(net4258));
 sg13g2_dlygate4sd3_1 hold1277 (.A(_01299_),
    .X(net4259));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\i_spi.clock_divider[3] ),
    .X(net4260));
 sg13g2_dlygate4sd3_1 hold1279 (.A(\i_i2c_peri.i_i2c.m_axis_data_tdata_reg[3] ),
    .X(net4261));
 sg13g2_dlygate4sd3_1 hold1280 (.A(_01208_),
    .X(net4262));
 sg13g2_dlygate4sd3_1 hold1281 (.A(\i_tinyqv.mem.data_from_read[18] ),
    .X(net4263));
 sg13g2_dlygate4sd3_1 hold1282 (.A(_00505_),
    .X(net4264));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\i_wdt.counter[25] ),
    .X(net4265));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_00829_),
    .X(net4266));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\i_seal.value_reg[10] ),
    .X(net4267));
 sg13g2_dlygate4sd3_1 hold1286 (.A(_00953_),
    .X(net4268));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\i_tinyqv.cpu.instr_data[1][3] ),
    .X(net4269));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_00462_),
    .X(net4270));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\i_i2c_peri.i_i2c.m_axis_data_tvalid_reg ),
    .X(net4271));
 sg13g2_dlygate4sd3_1 hold1290 (.A(_01312_),
    .X(net4272));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\i_seal.mono_count[11] ),
    .X(net4273));
 sg13g2_dlygate4sd3_1 hold1292 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[4] ),
    .X(net4274));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\i_tinyqv.cpu.i_core.mepc[2] ),
    .X(net4275));
 sg13g2_dlygate4sd3_1 hold1294 (.A(_00766_),
    .X(net4276));
 sg13g2_dlygate4sd3_1 hold1295 (.A(\i_latch_mem.data_out[6] ),
    .X(net4277));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\i_seal.crc_init ),
    .X(net4278));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_01185_),
    .X(net4279));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\i_crc16.bit_cnt[1] ),
    .X(net4280));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .X(net4281));
 sg13g2_dlygate4sd3_1 hold1300 (.A(_00529_),
    .X(net4282));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .X(net4283));
 sg13g2_dlygate4sd3_1 hold1302 (.A(_00082_),
    .X(net4284));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .X(net4285));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_00787_),
    .X(net4286));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\i_tinyqv.cpu.imm[24] ),
    .X(net4287));
 sg13g2_dlygate4sd3_1 hold1306 (.A(\i_latch_mem.genblk1[21].l_ram.data_out[7] ),
    .X(net4288));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\i_i2c_peri.i_i2c.missed_ack_reg ),
    .X(net4289));
 sg13g2_dlygate4sd3_1 hold1308 (.A(_07088_),
    .X(net4290));
 sg13g2_dlygate4sd3_1 hold1309 (.A(\i_tinyqv.cpu.imm[28] ),
    .X(net4291));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\i_i2c_peri.addr_latch[4] ),
    .X(net4292));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\i_rtc.us_count[5] ),
    .X(net4293));
 sg13g2_dlygate4sd3_1 hold1312 (.A(\i_latch_mem.data_out[4] ),
    .X(net4294));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\i_uart_rx.recieved_data[7] ),
    .X(net4295));
 sg13g2_dlygate4sd3_1 hold1314 (.A(\i_tinyqv.cpu.i_core.mepc[19] ),
    .X(net4296));
 sg13g2_dlygate4sd3_1 hold1315 (.A(_01132_),
    .X(net4297));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\reset_hold_counter[1] ),
    .X(net4298));
 sg13g2_dlygate4sd3_1 hold1317 (.A(\addr[22] ),
    .X(net4299));
 sg13g2_dlygate4sd3_1 hold1318 (.A(_01175_),
    .X(net4300));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\addr[18] ),
    .X(net4301));
 sg13g2_dlygate4sd3_1 hold1320 (.A(_01171_),
    .X(net4302));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\i_seal.crc_byte[2] ),
    .X(net4303));
 sg13g2_dlygate4sd3_1 hold1322 (.A(_01093_),
    .X(net4304));
 sg13g2_dlygate4sd3_1 hold1323 (.A(\i_rtc.us_count[15] ),
    .X(net4305));
 sg13g2_dlygate4sd3_1 hold1324 (.A(_06271_),
    .X(net4306));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_00852_),
    .X(net4307));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\i_seal.mono_count[7] ),
    .X(net4308));
 sg13g2_dlygate4sd3_1 hold1327 (.A(\i_tinyqv.cpu.data_ready_sync ),
    .X(net4309));
 sg13g2_dlygate4sd3_1 hold1328 (.A(_00664_),
    .X(net4310));
 sg13g2_dlygate4sd3_1 hold1329 (.A(\i_seal.session_ctr_in[2] ),
    .X(net4311));
 sg13g2_dlygate4sd3_1 hold1330 (.A(_00978_),
    .X(net4312));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\i2c_data_out[6] ),
    .X(net4313));
 sg13g2_dlygate4sd3_1 hold1332 (.A(\i_seal.sealed_mono[31] ),
    .X(net4314));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .X(net4315));
 sg13g2_dlygate4sd3_1 hold1334 (.A(_05823_),
    .X(net4316));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\i_seal.value_reg[19] ),
    .X(net4317));
 sg13g2_dlygate4sd3_1 hold1336 (.A(_00962_),
    .X(net4318));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\i_seal.mono_count[4] ),
    .X(net4319));
 sg13g2_dlygate4sd3_1 hold1338 (.A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .X(net4320));
 sg13g2_dlygate4sd3_1 hold1339 (.A(_04563_),
    .X(net4321));
 sg13g2_dlygate4sd3_1 hold1340 (.A(\reset_hold_counter[4] ),
    .X(net4322));
 sg13g2_dlygate4sd3_1 hold1341 (.A(_04543_),
    .X(net4323));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\i_seal.value_reg[26] ),
    .X(net4324));
 sg13g2_dlygate4sd3_1 hold1343 (.A(_00969_),
    .X(net4325));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\i_seal.sealed_mono[18] ),
    .X(net4326));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\i_seal.value_reg[27] ),
    .X(net4327));
 sg13g2_dlygate4sd3_1 hold1346 (.A(_00970_),
    .X(net4328));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\i_i2c_peri.i_i2c.phy_rx_data_reg ),
    .X(net4329));
 sg13g2_dlygate4sd3_1 hold1348 (.A(_01694_),
    .X(net4330));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\i_i2c_peri.cmd_addr_reg[3] ),
    .X(net4331));
 sg13g2_dlygate4sd3_1 hold1350 (.A(_01297_),
    .X(net4332));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\timer_count[11] ),
    .X(net4333));
 sg13g2_dlygate4sd3_1 hold1352 (.A(_04458_),
    .X(net4334));
 sg13g2_dlygate4sd3_1 hold1353 (.A(_00428_),
    .X(net4335));
 sg13g2_dlygate4sd3_1 hold1354 (.A(\i_seal.cur_mono[21] ),
    .X(net4336));
 sg13g2_dlygate4sd3_1 hold1355 (.A(_00932_),
    .X(net4337));
 sg13g2_dlygate4sd3_1 hold1356 (.A(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .X(net4338));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\i_i2c_peri.i_i2c.data_reg[0] ),
    .X(net4339));
 sg13g2_dlygate4sd3_1 hold1358 (.A(_01206_),
    .X(net4340));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .X(net4341));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\addr[9] ),
    .X(net4342));
 sg13g2_dlygate4sd3_1 hold1361 (.A(_01162_),
    .X(net4343));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .X(net4344));
 sg13g2_dlygate4sd3_1 hold1363 (.A(_05996_),
    .X(net4345));
 sg13g2_dlygate4sd3_1 hold1364 (.A(\i_wdt.counter[30] ),
    .X(net4346));
 sg13g2_dlygate4sd3_1 hold1365 (.A(_06218_),
    .X(net4347));
 sg13g2_dlygate4sd3_1 hold1366 (.A(_00834_),
    .X(net4348));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\i_seal.cur_mono[12] ),
    .X(net4349));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\i_tinyqv.cpu.i_core.mepc[23] ),
    .X(net4350));
 sg13g2_dlygate4sd3_1 hold1369 (.A(_00767_),
    .X(net4351));
 sg13g2_dlygate4sd3_1 hold1370 (.A(\i_tinyqv.cpu.alu_op[1] ),
    .X(net4352));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\i_seal.read_seq[0] ),
    .X(net4353));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\i_uart_tx.cycle_counter[0] ),
    .X(net4354));
 sg13g2_dlygate4sd3_1 hold1373 (.A(_07163_),
    .X(net4355));
 sg13g2_dlygate4sd3_1 hold1374 (.A(_01338_),
    .X(net4356));
 sg13g2_dlygate4sd3_1 hold1375 (.A(\i_tinyqv.cpu.i_core.mip[0] ),
    .X(net4357));
 sg13g2_dlygate4sd3_1 hold1376 (.A(_01659_),
    .X(net4358));
 sg13g2_dlygate4sd3_1 hold1377 (.A(\i_i2c_peri.cmd_addr_reg[2] ),
    .X(net4359));
 sg13g2_dlygate4sd3_1 hold1378 (.A(_01296_),
    .X(net4360));
 sg13g2_dlygate4sd3_1 hold1379 (.A(\i_tinyqv.cpu.imm[25] ),
    .X(net4361));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\i_latch_mem.genblk1[29].l_ram.data_out[0] ),
    .X(net4362));
 sg13g2_dlygate4sd3_1 hold1381 (.A(\i_seal.byte_sent ),
    .X(net4363));
 sg13g2_dlygate4sd3_1 hold1382 (.A(_06394_),
    .X(net4364));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\i_seal.cur_mono[23] ),
    .X(net4365));
 sg13g2_dlygate4sd3_1 hold1384 (.A(_00934_),
    .X(net4366));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\i_i2c_peri.i_i2c.data_reg[4] ),
    .X(net4367));
 sg13g2_dlygate4sd3_1 hold1386 (.A(_01646_),
    .X(net4368));
 sg13g2_dlygate4sd3_1 hold1387 (.A(\i2c_config_out[1] ),
    .X(net4369));
 sg13g2_dlygate4sd3_1 hold1388 (.A(_01268_),
    .X(net4370));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\i_seal.cur_mono[11] ),
    .X(net4371));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\i_tinyqv.mem.data_from_read[23] ),
    .X(net4372));
 sg13g2_dlygate4sd3_1 hold1391 (.A(_00510_),
    .X(net4373));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\i_i2c_peri.i_i2c.data_reg[3] ),
    .X(net4374));
 sg13g2_dlygate4sd3_1 hold1393 (.A(_01647_),
    .X(net4375));
 sg13g2_dlygate4sd3_1 hold1394 (.A(\i_tinyqv.cpu.imm[26] ),
    .X(net4376));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\i_i2c_peri.i_i2c.phy_state_reg[1] ),
    .X(net4377));
 sg13g2_dlygate4sd3_1 hold1396 (.A(_06888_),
    .X(net4378));
 sg13g2_dlygate4sd3_1 hold1397 (.A(\i_wdt.enabled ),
    .X(net4379));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .X(net4380));
 sg13g2_dlygate4sd3_1 hold1399 (.A(_00528_),
    .X(net4381));
 sg13g2_dlygate4sd3_1 hold1400 (.A(\i_seal.value_reg[29] ),
    .X(net4382));
 sg13g2_dlygate4sd3_1 hold1401 (.A(_00972_),
    .X(net4383));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\i_seal.sealed_mono[29] ),
    .X(net4384));
 sg13g2_dlygate4sd3_1 hold1403 (.A(\timer_count[15] ),
    .X(net4385));
 sg13g2_dlygate4sd3_1 hold1404 (.A(_04469_),
    .X(net4386));
 sg13g2_dlygate4sd3_1 hold1405 (.A(_00432_),
    .X(net4387));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .X(net4388));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_06104_),
    .X(net4389));
 sg13g2_dlygate4sd3_1 hold1408 (.A(_00794_),
    .X(net4390));
 sg13g2_dlygate4sd3_1 hold1409 (.A(\i_wdt.counter[31] ),
    .X(net4391));
 sg13g2_dlygate4sd3_1 hold1410 (.A(_00835_),
    .X(net4392));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\i_seal.value_reg[25] ),
    .X(net4393));
 sg13g2_dlygate4sd3_1 hold1412 (.A(_00968_),
    .X(net4394));
 sg13g2_dlygate4sd3_1 hold1413 (.A(\i_wdt.counter[7] ),
    .X(net4395));
 sg13g2_dlygate4sd3_1 hold1414 (.A(_00811_),
    .X(net4396));
 sg13g2_dlygate4sd3_1 hold1415 (.A(\i_tinyqv.cpu.mem_op_increment_reg ),
    .X(net4397));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .X(net4398));
 sg13g2_dlygate4sd3_1 hold1417 (.A(_00735_),
    .X(net4399));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\addr[14] ),
    .X(net4400));
 sg13g2_dlygate4sd3_1 hold1419 (.A(_01167_),
    .X(net4401));
 sg13g2_dlygate4sd3_1 hold1420 (.A(\addr[4] ),
    .X(net4402));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\i_seal.sealed_mono[30] ),
    .X(net4403));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\i_tinyqv.cpu.i_core.mepc[11] ),
    .X(net4404));
 sg13g2_dlygate4sd3_1 hold1423 (.A(_01124_),
    .X(net4405));
 sg13g2_dlygate4sd3_1 hold1424 (.A(\i_tinyqv.cpu.imm[18] ),
    .X(net4406));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\i_tinyqv.cpu.instr_data[3][9] ),
    .X(net4407));
 sg13g2_dlygate4sd3_1 hold1426 (.A(_01260_),
    .X(net4408));
 sg13g2_dlygate4sd3_1 hold1427 (.A(\i_tinyqv.cpu.is_branch ),
    .X(net4409));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\i_tinyqv.cpu.i_core.mepc[8] ),
    .X(net4410));
 sg13g2_dlygate4sd3_1 hold1429 (.A(_01121_),
    .X(net4411));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\i_tinyqv.cpu.i_core.mepc[7] ),
    .X(net4412));
 sg13g2_dlygate4sd3_1 hold1431 (.A(\i_tinyqv.cpu.i_core.mepc[18] ),
    .X(net4413));
 sg13g2_dlygate4sd3_1 hold1432 (.A(_01127_),
    .X(net4414));
 sg13g2_dlygate4sd3_1 hold1433 (.A(\i_rtc.us_count[6] ),
    .X(net4415));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .X(net4416));
 sg13g2_dlygate4sd3_1 hold1435 (.A(_01112_),
    .X(net4417));
 sg13g2_dlygate4sd3_1 hold1436 (.A(\i_tinyqv.cpu.instr_data[1][7] ),
    .X(net4418));
 sg13g2_dlygate4sd3_1 hold1437 (.A(_00466_),
    .X(net4419));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\i_seal.value_reg[2] ),
    .X(net4420));
 sg13g2_dlygate4sd3_1 hold1439 (.A(_00945_),
    .X(net4421));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\i_latch_mem.data_out[12] ),
    .X(net4422));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\i2c_data_out[2] ),
    .X(net4423));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\i_tinyqv.cpu.instr_data[3][11] ),
    .X(net4424));
 sg13g2_dlygate4sd3_1 hold1443 (.A(_01262_),
    .X(net4425));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .X(net4426));
 sg13g2_dlygate4sd3_1 hold1445 (.A(\i_tinyqv.cpu.instr_data[3][7] ),
    .X(net4427));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_01258_),
    .X(net4428));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\i_seal.sealed_mono[13] ),
    .X(net4429));
 sg13g2_dlygate4sd3_1 hold1448 (.A(\i_seal.value_reg[11] ),
    .X(net4430));
 sg13g2_dlygate4sd3_1 hold1449 (.A(_00954_),
    .X(net4431));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\i_wdt.counter[26] ),
    .X(net4432));
 sg13g2_dlygate4sd3_1 hold1451 (.A(_00830_),
    .X(net4433));
 sg13g2_dlygate4sd3_1 hold1452 (.A(\i_tinyqv.cpu.instr_data[1][4] ),
    .X(net4434));
 sg13g2_dlygate4sd3_1 hold1453 (.A(_00463_),
    .X(net4435));
 sg13g2_dlygate4sd3_1 hold1454 (.A(timer_irq),
    .X(net4436));
 sg13g2_dlygate4sd3_1 hold1455 (.A(_04531_),
    .X(net4437));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\i_tinyqv.cpu.i_core.mepc[5] ),
    .X(net4438));
 sg13g2_dlygate4sd3_1 hold1457 (.A(_01114_),
    .X(net4439));
 sg13g2_dlygate4sd3_1 hold1458 (.A(\i_tinyqv.cpu.counter[3] ),
    .X(net4440));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\i_i2c_peri.i_i2c.data_reg[6] ),
    .X(net4441));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_01644_),
    .X(net4442));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\i_seal.sealed_value[5] ),
    .X(net4443));
 sg13g2_dlygate4sd3_1 hold1462 (.A(_00948_),
    .X(net4444));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\i_i2c_peri.i_i2c.scl_o_reg ),
    .X(net4445));
 sg13g2_dlygate4sd3_1 hold1464 (.A(_01204_),
    .X(net4446));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\i_tinyqv.cpu.imm[13] ),
    .X(net4447));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\i_tinyqv.cpu.instr_data[3][5] ),
    .X(net4448));
 sg13g2_dlygate4sd3_1 hold1467 (.A(_01256_),
    .X(net4449));
 sg13g2_dlygate4sd3_1 hold1468 (.A(\gpio_out[2] ),
    .X(net4450));
 sg13g2_dlygate4sd3_1 hold1469 (.A(_00372_),
    .X(net4451));
 sg13g2_dlygate4sd3_1 hold1470 (.A(\i_tinyqv.cpu.instr_data[0][9] ),
    .X(net4452));
 sg13g2_dlygate4sd3_1 hold1471 (.A(_01140_),
    .X(net4453));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\i_tinyqv.cpu.instr_data[0][12] ),
    .X(net4454));
 sg13g2_dlygate4sd3_1 hold1473 (.A(_01143_),
    .X(net4455));
 sg13g2_dlygate4sd3_1 hold1474 (.A(\gpio_out[5] ),
    .X(net4456));
 sg13g2_dlygate4sd3_1 hold1475 (.A(_00375_),
    .X(net4457));
 sg13g2_dlygate4sd3_1 hold1476 (.A(\i_tinyqv.cpu.instr_data[2][14] ),
    .X(net4458));
 sg13g2_dlygate4sd3_1 hold1477 (.A(_01198_),
    .X(net4459));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[7] ),
    .X(net4460));
 sg13g2_dlygate4sd3_1 hold1479 (.A(_01310_),
    .X(net4461));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\timer_count[22] ),
    .X(net4462));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_00439_),
    .X(net4463));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\i_tinyqv.cpu.instr_data[1][5] ),
    .X(net4464));
 sg13g2_dlygate4sd3_1 hold1483 (.A(_00464_),
    .X(net4465));
 sg13g2_dlygate4sd3_1 hold1484 (.A(\i_uart_tx.cycle_counter[6] ),
    .X(net4466));
 sg13g2_dlygate4sd3_1 hold1485 (.A(_07175_),
    .X(net4467));
 sg13g2_dlygate4sd3_1 hold1486 (.A(_01344_),
    .X(net4468));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\i_tinyqv.cpu.i_core.mepc[9] ),
    .X(net4469));
 sg13g2_dlygate4sd3_1 hold1488 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[0] ),
    .X(net4470));
 sg13g2_dlygate4sd3_1 hold1489 (.A(_01706_),
    .X(net4471));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\i_tinyqv.cpu.imm[17] ),
    .X(net4472));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\i_tinyqv.cpu.instr_data[2][9] ),
    .X(net4473));
 sg13g2_dlygate4sd3_1 hold1492 (.A(_01193_),
    .X(net4474));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\i_tinyqv.cpu.instr_data[1][13] ),
    .X(net4475));
 sg13g2_dlygate4sd3_1 hold1494 (.A(_00472_),
    .X(net4476));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\i_i2c_peri.i_i2c.data_reg[5] ),
    .X(net4477));
 sg13g2_dlygate4sd3_1 hold1496 (.A(_01645_),
    .X(net4478));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\i_seal.value_reg[3] ),
    .X(net4479));
 sg13g2_dlygate4sd3_1 hold1498 (.A(_00946_),
    .X(net4480));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\i_tinyqv.cpu.i_core.mepc[1] ),
    .X(net4481));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\i_tinyqv.cpu.instr_data[1][15] ),
    .X(net4482));
 sg13g2_dlygate4sd3_1 hold1501 (.A(_00474_),
    .X(net4483));
 sg13g2_dlygate4sd3_1 hold1502 (.A(\i_tinyqv.cpu.instr_data[1][10] ),
    .X(net4484));
 sg13g2_dlygate4sd3_1 hold1503 (.A(_00469_),
    .X(net4485));
 sg13g2_dlygate4sd3_1 hold1504 (.A(\i2c_data_out[0] ),
    .X(net4486));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\i_tinyqv.cpu.instr_data[3][12] ),
    .X(net4487));
 sg13g2_dlygate4sd3_1 hold1506 (.A(_01263_),
    .X(net4488));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\i_seal.sealed_mono[8] ),
    .X(net4489));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\i_i2c_peri.i_i2c.delay_reg[10] ),
    .X(net4490));
 sg13g2_dlygate4sd3_1 hold1509 (.A(_06957_),
    .X(net4491));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\i_tinyqv.cpu.instr_data[0][15] ),
    .X(net4492));
 sg13g2_dlygate4sd3_1 hold1511 (.A(_01146_),
    .X(net4493));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\i_tinyqv.cpu.instr_data[3][6] ),
    .X(net4494));
 sg13g2_dlygate4sd3_1 hold1513 (.A(_01257_),
    .X(net4495));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\i_tinyqv.cpu.instr_data[0][11] ),
    .X(net4496));
 sg13g2_dlygate4sd3_1 hold1515 (.A(_01142_),
    .X(net4497));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\i_tinyqv.cpu.instr_data[0][7] ),
    .X(net4498));
 sg13g2_dlygate4sd3_1 hold1517 (.A(_01138_),
    .X(net4499));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\i_rtc.us_count[9] ),
    .X(net4500));
 sg13g2_dlygate4sd3_1 hold1519 (.A(_06260_),
    .X(net4501));
 sg13g2_dlygate4sd3_1 hold1520 (.A(_00846_),
    .X(net4502));
 sg13g2_dlygate4sd3_1 hold1521 (.A(\i_tinyqv.cpu.instr_data[0][5] ),
    .X(net4503));
 sg13g2_dlygate4sd3_1 hold1522 (.A(_01136_),
    .X(net4504));
 sg13g2_dlygate4sd3_1 hold1523 (.A(\i_tinyqv.cpu.instr_data[0][13] ),
    .X(net4505));
 sg13g2_dlygate4sd3_1 hold1524 (.A(_01144_),
    .X(net4506));
 sg13g2_dlygate4sd3_1 hold1525 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[6] ),
    .X(net4507));
 sg13g2_dlygate4sd3_1 hold1526 (.A(_01309_),
    .X(net4508));
 sg13g2_dlygate4sd3_1 hold1527 (.A(\i_tinyqv.cpu.i_core.mepc[13] ),
    .X(net4509));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\i_tinyqv.cpu.i_core.mepc[6] ),
    .X(net4510));
 sg13g2_dlygate4sd3_1 hold1529 (.A(_01119_),
    .X(net4511));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\i_tinyqv.cpu.i_core.mepc[3] ),
    .X(net4512));
 sg13g2_dlygate4sd3_1 hold1531 (.A(\gpio_out[6] ),
    .X(net4513));
 sg13g2_dlygate4sd3_1 hold1532 (.A(_00376_),
    .X(net4514));
 sg13g2_dlygate4sd3_1 hold1533 (.A(\i_tinyqv.cpu.imm[30] ),
    .X(net4515));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\i_tinyqv.cpu.instr_data[1][14] ),
    .X(net4516));
 sg13g2_dlygate4sd3_1 hold1535 (.A(_00473_),
    .X(net4517));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\i_tinyqv.cpu.instr_data[2][5] ),
    .X(net4518));
 sg13g2_dlygate4sd3_1 hold1537 (.A(_01189_),
    .X(net4519));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\session_ms_div[6] ),
    .X(net4520));
 sg13g2_dlygate4sd3_1 hold1539 (.A(\i_tinyqv.cpu.instr_data[1][12] ),
    .X(net4521));
 sg13g2_dlygate4sd3_1 hold1540 (.A(_00471_),
    .X(net4522));
 sg13g2_dlygate4sd3_1 hold1541 (.A(\i_tinyqv.cpu.instr_data[2][11] ),
    .X(net4523));
 sg13g2_dlygate4sd3_1 hold1542 (.A(_01195_),
    .X(net4524));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\i_tinyqv.cpu.instr_data[2][15] ),
    .X(net4525));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_01199_),
    .X(net4526));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\i_seal.sealed_crc[5] ),
    .X(net4527));
 sg13g2_dlygate4sd3_1 hold1546 (.A(_00900_),
    .X(net4528));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\i_seal.sealed_crc[7] ),
    .X(net4529));
 sg13g2_dlygate4sd3_1 hold1548 (.A(_00902_),
    .X(net4530));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\addr[15] ),
    .X(net4531));
 sg13g2_dlygate4sd3_1 hold1550 (.A(_01168_),
    .X(net4532));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\i_tinyqv.cpu.imm[19] ),
    .X(net4533));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\i_rtc.us_count[0] ),
    .X(net4534));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\i_i2c_peri.i_i2c.data_reg[2] ),
    .X(net4535));
 sg13g2_dlygate4sd3_1 hold1554 (.A(_01648_),
    .X(net4536));
 sg13g2_dlygate4sd3_1 hold1555 (.A(\addr[17] ),
    .X(net4537));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\i_seal.session_locked ),
    .X(net4538));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\i_uart_rx.cycle_counter[4] ),
    .X(net4539));
 sg13g2_dlygate4sd3_1 hold1558 (.A(_07207_),
    .X(net4540));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\i_seal.sealed_value[0] ),
    .X(net4541));
 sg13g2_dlygate4sd3_1 hold1560 (.A(_00943_),
    .X(net4542));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\i_seal.cur_mono[20] ),
    .X(net4543));
 sg13g2_dlygate4sd3_1 hold1562 (.A(_00931_),
    .X(net4544));
 sg13g2_dlygate4sd3_1 hold1563 (.A(\i_tinyqv.cpu.instr_data[2][2] ),
    .X(net4545));
 sg13g2_dlygate4sd3_1 hold1564 (.A(_01186_),
    .X(net4546));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\i_tinyqv.cpu.instr_data[3][14] ),
    .X(net4547));
 sg13g2_dlygate4sd3_1 hold1566 (.A(_01265_),
    .X(net4548));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\i_tinyqv.cpu.instr_data[3][2] ),
    .X(net4549));
 sg13g2_dlygate4sd3_1 hold1568 (.A(_01253_),
    .X(net4550));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\i_tinyqv.cpu.i_core.mepc[17] ),
    .X(net4551));
 sg13g2_dlygate4sd3_1 hold1570 (.A(_05191_),
    .X(net4552));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\i_tinyqv.cpu.imm[15] ),
    .X(net4553));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\i_tinyqv.cpu.imm[12] ),
    .X(net4554));
 sg13g2_dlygate4sd3_1 hold1573 (.A(\i_seal.cur_mono[10] ),
    .X(net4555));
 sg13g2_dlygate4sd3_1 hold1574 (.A(_00921_),
    .X(net4556));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\i_tinyqv.cpu.instr_data[0][4] ),
    .X(net4557));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_01135_),
    .X(net4558));
 sg13g2_dlygate4sd3_1 hold1577 (.A(\i_seal.cur_mono[22] ),
    .X(net4559));
 sg13g2_dlygate4sd3_1 hold1578 (.A(_00933_),
    .X(net4560));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\i_seal.sealed_mono[19] ),
    .X(net4561));
 sg13g2_dlygate4sd3_1 hold1580 (.A(\i_tinyqv.cpu.instr_data[1][2] ),
    .X(net4562));
 sg13g2_dlygate4sd3_1 hold1581 (.A(_00461_),
    .X(net4563));
 sg13g2_dlygate4sd3_1 hold1582 (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .X(net4564));
 sg13g2_dlygate4sd3_1 hold1583 (.A(_00488_),
    .X(net4565));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\i_i2c_peri.i_i2c.mode_read_reg ),
    .X(net4566));
 sg13g2_dlygate4sd3_1 hold1585 (.A(_01250_),
    .X(net4567));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .X(net4568));
 sg13g2_dlygate4sd3_1 hold1587 (.A(_01111_),
    .X(net4569));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\i_tinyqv.cpu.instr_data[0][14] ),
    .X(net4570));
 sg13g2_dlygate4sd3_1 hold1589 (.A(_01145_),
    .X(net4571));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\i_seal.value_reg[1] ),
    .X(net4572));
 sg13g2_dlygate4sd3_1 hold1591 (.A(_00944_),
    .X(net4573));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\i_tinyqv.cpu.instr_data[2][7] ),
    .X(net4574));
 sg13g2_dlygate4sd3_1 hold1593 (.A(_01191_),
    .X(net4575));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\i_seal.cur_mono[6] ),
    .X(net4576));
 sg13g2_dlygate4sd3_1 hold1595 (.A(_00917_),
    .X(net4577));
 sg13g2_dlygate4sd3_1 hold1596 (.A(\addr[19] ),
    .X(net4578));
 sg13g2_dlygate4sd3_1 hold1597 (.A(_01172_),
    .X(net4579));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\i_rtc.us_count[10] ),
    .X(net4580));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_06262_),
    .X(net4581));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\i_tinyqv.cpu.instr_data[0][10] ),
    .X(net4582));
 sg13g2_dlygate4sd3_1 hold1601 (.A(_01141_),
    .X(net4583));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\i_tinyqv.cpu.instr_data[0][2] ),
    .X(net4584));
 sg13g2_dlygate4sd3_1 hold1603 (.A(_01133_),
    .X(net4585));
 sg13g2_dlygate4sd3_1 hold1604 (.A(\i_seal.sealed_crc[6] ),
    .X(net4586));
 sg13g2_dlygate4sd3_1 hold1605 (.A(_00901_),
    .X(net4587));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\i_tinyqv.cpu.i_core.mepc[14] ),
    .X(net4588));
 sg13g2_dlygate4sd3_1 hold1607 (.A(_01123_),
    .X(net4589));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\i_tinyqv.cpu.instr_data[2][4] ),
    .X(net4590));
 sg13g2_dlygate4sd3_1 hold1609 (.A(_01188_),
    .X(net4591));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\i_tinyqv.cpu.instr_data[1][11] ),
    .X(net4592));
 sg13g2_dlygate4sd3_1 hold1611 (.A(_00470_),
    .X(net4593));
 sg13g2_dlygate4sd3_1 hold1612 (.A(\i_tinyqv.cpu.instr_data[1][9] ),
    .X(net4594));
 sg13g2_dlygate4sd3_1 hold1613 (.A(_00468_),
    .X(net4595));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\i_seal.sealed_value[12] ),
    .X(net4596));
 sg13g2_dlygate4sd3_1 hold1615 (.A(_00955_),
    .X(net4597));
 sg13g2_dlygate4sd3_1 hold1616 (.A(\i_tinyqv.cpu.i_core.mepc[15] ),
    .X(net4598));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\addr[23] ),
    .X(net4599));
 sg13g2_dlygate4sd3_1 hold1618 (.A(_04822_),
    .X(net4600));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\i_tinyqv.cpu.instr_data[2][13] ),
    .X(net4601));
 sg13g2_dlygate4sd3_1 hold1620 (.A(_01197_),
    .X(net4602));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\i_spi.bits_remaining[2] ),
    .X(net4603));
 sg13g2_dlygate4sd3_1 hold1622 (.A(_01684_),
    .X(net4604));
 sg13g2_dlygate4sd3_1 hold1623 (.A(_01386_),
    .X(net4605));
 sg13g2_dlygate4sd3_1 hold1624 (.A(\i_uart_tx.cycle_counter[8] ),
    .X(net4606));
 sg13g2_dlygate4sd3_1 hold1625 (.A(_07179_),
    .X(net4607));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\gpio_out[0] ),
    .X(net4608));
 sg13g2_dlygate4sd3_1 hold1627 (.A(_00370_),
    .X(net4609));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\gpio_out[7] ),
    .X(net4610));
 sg13g2_dlygate4sd3_1 hold1629 (.A(_00377_),
    .X(net4611));
 sg13g2_dlygate4sd3_1 hold1630 (.A(\i_i2c_peri.i_i2c.s_axis_data_tlast ),
    .X(net4612));
 sg13g2_dlygate4sd3_1 hold1631 (.A(_01302_),
    .X(net4613));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\i_tinyqv.cpu.instr_data[1][6] ),
    .X(net4614));
 sg13g2_dlygate4sd3_1 hold1633 (.A(_00465_),
    .X(net4615));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\i_tinyqv.cpu.instr_data[3][13] ),
    .X(net4616));
 sg13g2_dlygate4sd3_1 hold1635 (.A(_01264_),
    .X(net4617));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\i_i2c_peri.i_i2c.delay_reg[9] ),
    .X(net4618));
 sg13g2_dlygate4sd3_1 hold1637 (.A(_06951_),
    .X(net4619));
 sg13g2_dlygate4sd3_1 hold1638 (.A(_01230_),
    .X(net4620));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\i_tinyqv.cpu.instr_data[2][6] ),
    .X(net4621));
 sg13g2_dlygate4sd3_1 hold1640 (.A(_01190_),
    .X(net4622));
 sg13g2_dlygate4sd3_1 hold1641 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .X(net4623));
 sg13g2_dlygate4sd3_1 hold1642 (.A(_00736_),
    .X(net4624));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .X(net4625));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\i_seal.cur_mono[3] ),
    .X(net4626));
 sg13g2_dlygate4sd3_1 hold1645 (.A(_00914_),
    .X(net4627));
 sg13g2_dlygate4sd3_1 hold1646 (.A(\i_wdt.counter[3] ),
    .X(net4628));
 sg13g2_dlygate4sd3_1 hold1647 (.A(_00807_),
    .X(net4629));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\addr[12] ),
    .X(net4630));
 sg13g2_dlygate4sd3_1 hold1649 (.A(_01165_),
    .X(net4631));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .X(net4632));
 sg13g2_dlygate4sd3_1 hold1651 (.A(_06099_),
    .X(net4633));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\i_tinyqv.cpu.instr_data[3][15] ),
    .X(net4634));
 sg13g2_dlygate4sd3_1 hold1653 (.A(_01266_),
    .X(net4635));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\gpio_out[3] ),
    .X(net4636));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\i_tinyqv.cpu.i_core.mip[1] ),
    .X(net4637));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\i_seal.sealed_mono[9] ),
    .X(net4638));
 sg13g2_dlygate4sd3_1 hold1657 (.A(_00920_),
    .X(net4639));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\i_i2c_peri.i_i2c.data_reg[1] ),
    .X(net4640));
 sg13g2_dlygate4sd3_1 hold1659 (.A(_01649_),
    .X(net4641));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\i_tinyqv.cpu.i_core.mepc[12] ),
    .X(net4642));
 sg13g2_dlygate4sd3_1 hold1661 (.A(_01125_),
    .X(net4643));
 sg13g2_dlygate4sd3_1 hold1662 (.A(\i_tinyqv.cpu.instr_data[2][12] ),
    .X(net4644));
 sg13g2_dlygate4sd3_1 hold1663 (.A(_01196_),
    .X(net4645));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\i_uart_tx.cycle_counter[4] ),
    .X(net4646));
 sg13g2_dlygate4sd3_1 hold1665 (.A(_07171_),
    .X(net4647));
 sg13g2_dlygate4sd3_1 hold1666 (.A(_01342_),
    .X(net4648));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\i_tinyqv.cpu.instr_data_in[3] ),
    .X(net4649));
 sg13g2_dlygate4sd3_1 hold1668 (.A(_00490_),
    .X(net4650));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\i2c_config_out[0] ),
    .X(net4651));
 sg13g2_dlygate4sd3_1 hold1670 (.A(_01267_),
    .X(net4652));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\i_seal.sealed_crc[13] ),
    .X(net4653));
 sg13g2_dlygate4sd3_1 hold1672 (.A(_00908_),
    .X(net4654));
 sg13g2_dlygate4sd3_1 hold1673 (.A(\i_seal.sealed_mono[16] ),
    .X(net4655));
 sg13g2_dlygate4sd3_1 hold1674 (.A(_00927_),
    .X(net4656));
 sg13g2_dlygate4sd3_1 hold1675 (.A(\i_tinyqv.cpu.instr_data[0][6] ),
    .X(net4657));
 sg13g2_dlygate4sd3_1 hold1676 (.A(_01137_),
    .X(net4658));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\addr[16] ),
    .X(net4659));
 sg13g2_dlygate4sd3_1 hold1678 (.A(_01169_),
    .X(net4660));
 sg13g2_dlygate4sd3_1 hold1679 (.A(\i_tinyqv.cpu.instr_data[3][10] ),
    .X(net4661));
 sg13g2_dlygate4sd3_1 hold1680 (.A(_01261_),
    .X(net4662));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\i_wdt.counter[21] ),
    .X(net4663));
 sg13g2_dlygate4sd3_1 hold1682 (.A(_06191_),
    .X(net4664));
 sg13g2_dlygate4sd3_1 hold1683 (.A(_00825_),
    .X(net4665));
 sg13g2_dlygate4sd3_1 hold1684 (.A(\i_tinyqv.cpu.instr_data[3][4] ),
    .X(net4666));
 sg13g2_dlygate4sd3_1 hold1685 (.A(_01255_),
    .X(net4667));
 sg13g2_dlygate4sd3_1 hold1686 (.A(\i_tinyqv.cpu.instr_data[2][10] ),
    .X(net4668));
 sg13g2_dlygate4sd3_1 hold1687 (.A(_01194_),
    .X(net4669));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\i_tinyqv.cpu.i_core.mcause[1] ),
    .X(net4670));
 sg13g2_dlygate4sd3_1 hold1689 (.A(_00457_),
    .X(net4671));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .X(net4672));
 sg13g2_dlygate4sd3_1 hold1691 (.A(_00737_),
    .X(net4673));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\session_ms_div[0] ),
    .X(net4674));
 sg13g2_dlygate4sd3_1 hold1693 (.A(\i_uart_tx.cycle_counter[3] ),
    .X(net4675));
 sg13g2_dlygate4sd3_1 hold1694 (.A(_07169_),
    .X(net4676));
 sg13g2_dlygate4sd3_1 hold1695 (.A(_01341_),
    .X(net4677));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .X(net4678));
 sg13g2_dlygate4sd3_1 hold1697 (.A(_00093_),
    .X(net4679));
 sg13g2_dlygate4sd3_1 hold1698 (.A(\i_rtc.us_count[19] ),
    .X(net4680));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\crc_peri_data[0] ),
    .X(net4681));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\i_seal.sealed_crc[0] ),
    .X(net4682));
 sg13g2_dlygate4sd3_1 hold1701 (.A(_00895_),
    .X(net4683));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\addr[24] ),
    .X(net4684));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\reset_hold_counter[2] ),
    .X(net4685));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .X(net4686));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\i_seal.sealed_crc[1] ),
    .X(net4687));
 sg13g2_dlygate4sd3_1 hold1706 (.A(_00896_),
    .X(net4688));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .X(net4689));
 sg13g2_dlygate4sd3_1 hold1708 (.A(_00560_),
    .X(net4690));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\i_uart_tx.cycle_counter[5] ),
    .X(net4691));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\pps_count[0] ),
    .X(net4692));
 sg13g2_dlygate4sd3_1 hold1711 (.A(_04376_),
    .X(net4693));
 sg13g2_dlygate4sd3_1 hold1712 (.A(_00397_),
    .X(net4694));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\i_i2c_peri.i_i2c.delay_reg[4] ),
    .X(net4695));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_01225_),
    .X(net4696));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\i_uart_rx.recieved_data[2] ),
    .X(net4697));
 sg13g2_dlygate4sd3_1 hold1716 (.A(_01352_),
    .X(net4698));
 sg13g2_dlygate4sd3_1 hold1717 (.A(\i_uart_rx.recieved_data[3] ),
    .X(net4699));
 sg13g2_dlygate4sd3_1 hold1718 (.A(\i_i2c_peri.i_i2c.delay_reg[8] ),
    .X(net4700));
 sg13g2_dlygate4sd3_1 hold1719 (.A(_01229_),
    .X(net4701));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\i_wdt.counter[19] ),
    .X(net4702));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_00823_),
    .X(net4703));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\i_rtc.us_count[13] ),
    .X(net4704));
 sg13g2_dlygate4sd3_1 hold1723 (.A(_06267_),
    .X(net4705));
 sg13g2_dlygate4sd3_1 hold1724 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .X(net4706));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ),
    .X(net4707));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\crc_peri_data[6] ),
    .X(net4708));
 sg13g2_dlygate4sd3_1 hold1727 (.A(_01336_),
    .X(net4709));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\i_i2c_peri.i_i2c.state_reg[1] ),
    .X(net4710));
 sg13g2_dlygate4sd3_1 hold1729 (.A(_06879_),
    .X(net4711));
 sg13g2_dlygate4sd3_1 hold1730 (.A(_06898_),
    .X(net4712));
 sg13g2_dlygate4sd3_1 hold1731 (.A(\i_uart_rx.cycle_counter[8] ),
    .X(net4713));
 sg13g2_dlygate4sd3_1 hold1732 (.A(_07215_),
    .X(net4714));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\i_uart_tx.fsm_state[3] ),
    .X(net4715));
 sg13g2_dlygate4sd3_1 hold1734 (.A(_01350_),
    .X(net4716));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\i_wdt.counter[5] ),
    .X(net4717));
 sg13g2_dlygate4sd3_1 hold1736 (.A(_00809_),
    .X(net4718));
 sg13g2_dlygate4sd3_1 hold1737 (.A(\crc16_read[4] ),
    .X(net4719));
 sg13g2_dlygate4sd3_1 hold1738 (.A(_00899_),
    .X(net4720));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\gpio_out[4] ),
    .X(net4721));
 sg13g2_dlygate4sd3_1 hold1740 (.A(_00374_),
    .X(net4722));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\i_i2c_peri.cmd_read_reg ),
    .X(net4723));
 sg13g2_dlygate4sd3_1 hold1742 (.A(_01292_),
    .X(net4724));
 sg13g2_dlygate4sd3_1 hold1743 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[2] ),
    .X(net4725));
 sg13g2_dlygate4sd3_1 hold1744 (.A(_01305_),
    .X(net4726));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\pps_count[9] ),
    .X(net4727));
 sg13g2_dlygate4sd3_1 hold1746 (.A(_04393_),
    .X(net4728));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[1] ),
    .X(net4729));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\i_tinyqv.cpu.i_core.mepc[16] ),
    .X(net4730));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\i_uart_rx.recieved_data[5] ),
    .X(net4731));
 sg13g2_dlygate4sd3_1 hold1750 (.A(_01356_),
    .X(net4732));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\i_rtc.seconds_out[24] ),
    .X(net4733));
 sg13g2_dlygate4sd3_1 hold1752 (.A(_06358_),
    .X(net4734));
 sg13g2_dlygate4sd3_1 hold1753 (.A(_00881_),
    .X(net4735));
 sg13g2_dlygate4sd3_1 hold1754 (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .X(net4736));
 sg13g2_dlygate4sd3_1 hold1755 (.A(_00572_),
    .X(net4737));
 sg13g2_dlygate4sd3_1 hold1756 (.A(\i_uart_rx.recieved_data[4] ),
    .X(net4738));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\reset_hold_counter[3] ),
    .X(net4739));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\i_spi.clock_count[0] ),
    .X(net4740));
 sg13g2_dlygate4sd3_1 hold1759 (.A(_01379_),
    .X(net4741));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\i_tinyqv.cpu.is_jal ),
    .X(net4742));
 sg13g2_dlygate4sd3_1 hold1761 (.A(_00674_),
    .X(net4743));
 sg13g2_dlygate4sd3_1 hold1762 (.A(\i_spi.clock_count[3] ),
    .X(net4744));
 sg13g2_dlygate4sd3_1 hold1763 (.A(_01672_),
    .X(net4745));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\i_tinyqv.cpu.imm[20] ),
    .X(net4746));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\i_seal.sealed_crc[2] ),
    .X(net4747));
 sg13g2_dlygate4sd3_1 hold1766 (.A(_00897_),
    .X(net4748));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[4] ),
    .X(net4749));
 sg13g2_dlygate4sd3_1 hold1768 (.A(_01307_),
    .X(net4750));
 sg13g2_dlygate4sd3_1 hold1769 (.A(\crc16_read[13] ),
    .X(net4751));
 sg13g2_dlygate4sd3_1 hold1770 (.A(_05862_),
    .X(net4752));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_00747_),
    .X(net4753));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\i_rtc.us_count[11] ),
    .X(net4754));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\timer_count[18] ),
    .X(net4755));
 sg13g2_dlygate4sd3_1 hold1774 (.A(_04478_),
    .X(net4756));
 sg13g2_dlygate4sd3_1 hold1775 (.A(_00435_),
    .X(net4757));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .X(net4758));
 sg13g2_dlygate4sd3_1 hold1777 (.A(_00574_),
    .X(net4759));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\i_i2c_peri.i_i2c.delay_reg[3] ),
    .X(net4760));
 sg13g2_dlygate4sd3_1 hold1779 (.A(_01224_),
    .X(net4761));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\i_uart_tx.fsm_state[2] ),
    .X(net4762));
 sg13g2_dlygate4sd3_1 hold1781 (.A(_01349_),
    .X(net4763));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\i_uart_rx.cycle_counter[7] ),
    .X(net4764));
 sg13g2_dlygate4sd3_1 hold1783 (.A(_07212_),
    .X(net4765));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\addr[21] ),
    .X(net4766));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[3] ),
    .X(net4767));
 sg13g2_dlygate4sd3_1 hold1786 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .X(net4768));
 sg13g2_dlygate4sd3_1 hold1787 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .X(net4769));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\i_tinyqv.cpu.instr_len[1] ),
    .X(net4770));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\i_spi.clock_count[2] ),
    .X(net4771));
 sg13g2_dlygate4sd3_1 hold1790 (.A(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .X(net4772));
 sg13g2_dlygate4sd3_1 hold1791 (.A(_00780_),
    .X(net4773));
 sg13g2_dlygate4sd3_1 hold1792 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .X(net4774));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\i_uart_rx.recieved_data[6] ),
    .X(net4775));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .X(net4776));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\i_seal.cur_mono[14] ),
    .X(net4777));
 sg13g2_dlygate4sd3_1 hold1796 (.A(_00925_),
    .X(net4778));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\addr[20] ),
    .X(net4779));
 sg13g2_dlygate4sd3_1 hold1798 (.A(_01173_),
    .X(net4780));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .X(net4781));
 sg13g2_dlygate4sd3_1 hold1800 (.A(_06044_),
    .X(net4782));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\i_i2c_peri.i_i2c.s_axis_cmd_ready_reg ),
    .X(net4783));
 sg13g2_dlygate4sd3_1 hold1802 (.A(\i_spi.data[0] ),
    .X(net4784));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\crc16_read[14] ),
    .X(net4785));
 sg13g2_dlygate4sd3_1 hold1804 (.A(_00749_),
    .X(net4786));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\i_uart_rx.fsm_state[2] ),
    .X(net4787));
 sg13g2_dlygate4sd3_1 hold1806 (.A(_01373_),
    .X(net4788));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\pps_count[5] ),
    .X(net4789));
 sg13g2_dlygate4sd3_1 hold1808 (.A(_04386_),
    .X(net4790));
 sg13g2_dlygate4sd3_1 hold1809 (.A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .X(net4791));
 sg13g2_dlygate4sd3_1 hold1810 (.A(_00563_),
    .X(net4792));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\crc_peri_data[4] ),
    .X(net4793));
 sg13g2_dlygate4sd3_1 hold1812 (.A(_01334_),
    .X(net4794));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .X(net4795));
 sg13g2_dlygate4sd3_1 hold1814 (.A(_00575_),
    .X(net4796));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\i_tinyqv.cpu.imm[31] ),
    .X(net4797));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .X(net4798));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\timer_count[20] ),
    .X(net4799));
 sg13g2_dlygate4sd3_1 hold1818 (.A(_04485_),
    .X(net4800));
 sg13g2_dlygate4sd3_1 hold1819 (.A(_00437_),
    .X(net4801));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .X(net4802));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\i_rtc.us_count[16] ),
    .X(net4803));
 sg13g2_dlygate4sd3_1 hold1822 (.A(_06273_),
    .X(net4804));
 sg13g2_dlygate4sd3_1 hold1823 (.A(\i2c_config_out[3] ),
    .X(net4805));
 sg13g2_dlygate4sd3_1 hold1824 (.A(_01270_),
    .X(net4806));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .X(net4807));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .X(net4808));
 sg13g2_dlygate4sd3_1 hold1827 (.A(_00571_),
    .X(net4809));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .X(net4810));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .X(net4811));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\i_i2c_peri.i_i2c.s_axis_data_tdata[5] ),
    .X(net4812));
 sg13g2_dlygate4sd3_1 hold1831 (.A(_01308_),
    .X(net4813));
 sg13g2_dlygate4sd3_1 hold1832 (.A(\crc_peri_data[5] ),
    .X(net4814));
 sg13g2_dlygate4sd3_1 hold1833 (.A(_01335_),
    .X(net4815));
 sg13g2_dlygate4sd3_1 hold1834 (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .X(net4816));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\i_wdt.counter[17] ),
    .X(net4817));
 sg13g2_dlygate4sd3_1 hold1836 (.A(_06180_),
    .X(net4818));
 sg13g2_dlygate4sd3_1 hold1837 (.A(_00821_),
    .X(net4819));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\i_uart_rx.cycle_counter[5] ),
    .X(net4820));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\i_uart_rx.cycle_counter[2] ),
    .X(net4821));
 sg13g2_dlygate4sd3_1 hold1840 (.A(_07204_),
    .X(net4822));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\i_i2c_peri.i_i2c.sda_o_reg ),
    .X(net4823));
 sg13g2_dlygate4sd3_1 hold1842 (.A(_01203_),
    .X(net4824));
 sg13g2_dlygate4sd3_1 hold1843 (.A(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .X(net4825));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\gpio_out_sel[7] ),
    .X(net4826));
 sg13g2_dlygate4sd3_1 hold1845 (.A(_00369_),
    .X(net4827));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\i_tinyqv.cpu.i_core.mie[0] ),
    .X(net4828));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\session_ms_div[3] ),
    .X(net4829));
 sg13g2_dlygate4sd3_1 hold1848 (.A(_00382_),
    .X(net4830));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\i_tinyqv.cpu.imm[21] ),
    .X(net4831));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\crc16_read[0] ),
    .X(net4832));
 sg13g2_dlygate4sd3_1 hold1851 (.A(_01322_),
    .X(net4833));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\gpio_out_sel[1] ),
    .X(net4834));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\i_tinyqv.cpu.imm[23] ),
    .X(net4835));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .X(net4836));
 sg13g2_dlygate4sd3_1 hold1855 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .X(net4837));
 sg13g2_dlygate4sd3_1 hold1856 (.A(\i_tinyqv.cpu.instr_len[2] ),
    .X(net4838));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .X(net4839));
 sg13g2_dlygate4sd3_1 hold1858 (.A(_06071_),
    .X(net4840));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .X(net4841));
 sg13g2_dlygate4sd3_1 hold1860 (.A(_05835_),
    .X(net4842));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\i_seal.sealed_crc[3] ),
    .X(net4843));
 sg13g2_dlygate4sd3_1 hold1862 (.A(_00898_),
    .X(net4844));
 sg13g2_dlygate4sd3_1 hold1863 (.A(\us_divider[4] ),
    .X(net4845));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\i_tinyqv.cpu.imm[14] ),
    .X(net4846));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .X(net4847));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\crc_peri_data[3] ),
    .X(net4848));
 sg13g2_dlygate4sd3_1 hold1867 (.A(_01333_),
    .X(net4849));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\crc16_read[15] ),
    .X(net4850));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .X(net4851));
 sg13g2_dlygate4sd3_1 hold1870 (.A(_00573_),
    .X(net4852));
 sg13g2_dlygate4sd3_1 hold1871 (.A(\pps_count[3] ),
    .X(net4853));
 sg13g2_dlygate4sd3_1 hold1872 (.A(_04383_),
    .X(net4854));
 sg13g2_dlygate4sd3_1 hold1873 (.A(_00400_),
    .X(net4855));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\pps_count[4] ),
    .X(net4856));
 sg13g2_dlygate4sd3_1 hold1875 (.A(_04385_),
    .X(net4857));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\i_tinyqv.cpu.imm[16] ),
    .X(net4858));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\i_tinyqv.mem.instr_active ),
    .X(net4859));
 sg13g2_dlygate4sd3_1 hold1878 (.A(_04780_),
    .X(net4860));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\i_rtc.us_count[7] ),
    .X(net4861));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\i2c_config_out[4] ),
    .X(net4862));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\i_rtc.us_count[14] ),
    .X(net4863));
 sg13g2_dlygate4sd3_1 hold1882 (.A(_06270_),
    .X(net4864));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\i_i2c_peri.i_i2c.bit_count_reg[3] ),
    .X(net4865));
 sg13g2_dlygate4sd3_1 hold1884 (.A(_00757_),
    .X(net4866));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .X(net4867));
 sg13g2_dlygate4sd3_1 hold1886 (.A(_05834_),
    .X(net4868));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\i_wdt.counter[27] ),
    .X(net4869));
 sg13g2_dlygate4sd3_1 hold1888 (.A(_06211_),
    .X(net4870));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\i_i2c_peri.i_i2c.delay_reg[5] ),
    .X(net4871));
 sg13g2_dlygate4sd3_1 hold1890 (.A(_01226_),
    .X(net4872));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\i_tinyqv.mem.q_ctrl.data_req ),
    .X(net4873));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\crc16_read[2] ),
    .X(net4874));
 sg13g2_dlygate4sd3_1 hold1893 (.A(_01323_),
    .X(net4875));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .X(net4876));
 sg13g2_dlygate4sd3_1 hold1895 (.A(\data_to_write[18] ),
    .X(net4877));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .X(net4878));
 sg13g2_dlygate4sd3_1 hold1897 (.A(_00487_),
    .X(net4879));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .X(net4880));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\i_i2c_peri.i_i2c.bit_count_reg[2] ),
    .X(net4881));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\pps_count[2] ),
    .X(net4882));
 sg13g2_dlygate4sd3_1 hold1901 (.A(_04381_),
    .X(net4883));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .X(net4884));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\i_i2c_peri.i_i2c.delay_reg[2] ),
    .X(net4885));
 sg13g2_dlygate4sd3_1 hold1904 (.A(_01223_),
    .X(net4886));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .X(net4887));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\pps_count[8] ),
    .X(net4888));
 sg13g2_dlygate4sd3_1 hold1907 (.A(_04392_),
    .X(net4889));
 sg13g2_dlygate4sd3_1 hold1908 (.A(_00405_),
    .X(net4890));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\i_uart_tx.cycle_counter[1] ),
    .X(net4891));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\data_to_write[16] ),
    .X(net4892));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\i_wdt.counter[28] ),
    .X(net4893));
 sg13g2_dlygate4sd3_1 hold1912 (.A(_00832_),
    .X(net4894));
 sg13g2_dlygate4sd3_1 hold1913 (.A(\gpio_out_sel[4] ),
    .X(net4895));
 sg13g2_dlygate4sd3_1 hold1914 (.A(\crc_peri_data[7] ),
    .X(net4896));
 sg13g2_dlygate4sd3_1 hold1915 (.A(\i2c_config_out[5] ),
    .X(net4897));
 sg13g2_dlygate4sd3_1 hold1916 (.A(\i2c_config_out[6] ),
    .X(net4898));
 sg13g2_dlygate4sd3_1 hold1917 (.A(\i_i2c_peri.i_i2c.delay_reg[11] ),
    .X(net4899));
 sg13g2_dlygate4sd3_1 hold1918 (.A(_01232_),
    .X(net4900));
 sg13g2_dlygate4sd3_1 hold1919 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .X(net4901));
 sg13g2_dlygate4sd3_1 hold1920 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .X(net4902));
 sg13g2_dlygate4sd3_1 hold1921 (.A(\i_i2c_peri.cmd_write_m_reg ),
    .X(net4903));
 sg13g2_dlygate4sd3_1 hold1922 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .X(net4904));
 sg13g2_dlygate4sd3_1 hold1923 (.A(\data_to_write[22] ),
    .X(net4905));
 sg13g2_dlygate4sd3_1 hold1924 (.A(\i_i2c_peri.i_i2c.delay_reg[6] ),
    .X(net4906));
 sg13g2_dlygate4sd3_1 hold1925 (.A(\i_seal.crc_byte[6] ),
    .X(net4907));
 sg13g2_dlygate4sd3_1 hold1926 (.A(_06691_),
    .X(net4908));
 sg13g2_dlygate4sd3_1 hold1927 (.A(_01097_),
    .X(net4909));
 sg13g2_dlygate4sd3_1 hold1928 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .X(net4910));
 sg13g2_dlygate4sd3_1 hold1929 (.A(_00524_),
    .X(net4911));
 sg13g2_dlygate4sd3_1 hold1930 (.A(\data_to_write[19] ),
    .X(net4912));
 sg13g2_dlygate4sd3_1 hold1931 (.A(_00436_),
    .X(net4913));
 sg13g2_dlygate4sd3_1 hold1932 (.A(\data_to_write[17] ),
    .X(net4914));
 sg13g2_dlygate4sd3_1 hold1933 (.A(_00434_),
    .X(net4915));
 sg13g2_dlygate4sd3_1 hold1934 (.A(\i_spi.bits_remaining[1] ),
    .X(net4916));
 sg13g2_dlygate4sd3_1 hold1935 (.A(\pps_count[14] ),
    .X(net4917));
 sg13g2_dlygate4sd3_1 hold1936 (.A(\gpio_out_sel[5] ),
    .X(net4918));
 sg13g2_dlygate4sd3_1 hold1937 (.A(\pps_count[11] ),
    .X(net4919));
 sg13g2_dlygate4sd3_1 hold1938 (.A(\i_tinyqv.cpu.data_read_n[0] ),
    .X(net4920));
 sg13g2_dlygate4sd3_1 hold1939 (.A(_05346_),
    .X(net4921));
 sg13g2_dlygate4sd3_1 hold1940 (.A(_00653_),
    .X(net4922));
 sg13g2_dlygate4sd3_1 hold1941 (.A(\i2c_config_out[15] ),
    .X(net4923));
 sg13g2_dlygate4sd3_1 hold1942 (.A(_06979_),
    .X(net4924));
 sg13g2_dlygate4sd3_1 hold1943 (.A(_01236_),
    .X(net4925));
 sg13g2_dlygate4sd3_1 hold1944 (.A(\pps_count[7] ),
    .X(net4926));
 sg13g2_dlygate4sd3_1 hold1945 (.A(\data_to_write[28] ),
    .X(net4927));
 sg13g2_dlygate4sd3_1 hold1946 (.A(\data_to_write[23] ),
    .X(net4928));
 sg13g2_dlygate4sd3_1 hold1947 (.A(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .X(net4929));
 sg13g2_dlygate4sd3_1 hold1948 (.A(_00578_),
    .X(net4930));
 sg13g2_dlygate4sd3_1 hold1949 (.A(\i2c_config_out[7] ),
    .X(net4931));
 sg13g2_dlygate4sd3_1 hold1950 (.A(\i_tinyqv.cpu.imm[22] ),
    .X(net4932));
 sg13g2_dlygate4sd3_1 hold1951 (.A(\data_to_write[21] ),
    .X(net4933));
 sg13g2_dlygate4sd3_1 hold1952 (.A(\gpio_out_sel[0] ),
    .X(net4934));
 sg13g2_dlygate4sd3_1 hold1953 (.A(\i_i2c_peri.i_i2c.delay_reg[1] ),
    .X(net4935));
 sg13g2_dlygate4sd3_1 hold1954 (.A(_01222_),
    .X(net4936));
 sg13g2_dlygate4sd3_1 hold1955 (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .X(net4937));
 sg13g2_dlygate4sd3_1 hold1956 (.A(\crc16_read[11] ),
    .X(net4938));
 sg13g2_dlygate4sd3_1 hold1957 (.A(_00746_),
    .X(net4939));
 sg13g2_dlygate4sd3_1 hold1958 (.A(\i_uart_tx.data_to_send[0] ),
    .X(net4940));
 sg13g2_dlygate4sd3_1 hold1959 (.A(_00836_),
    .X(net4941));
 sg13g2_dlygate4sd3_1 hold1960 (.A(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .X(net4942));
 sg13g2_dlygate4sd3_1 hold1961 (.A(\crc16_read[8] ),
    .X(net4943));
 sg13g2_dlygate4sd3_1 hold1962 (.A(_00743_),
    .X(net4944));
 sg13g2_dlygate4sd3_1 hold1963 (.A(\i_tinyqv.cpu.i_core.mstatus_mte ),
    .X(net4945));
 sg13g2_dlygate4sd3_1 hold1964 (.A(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .X(net4946));
 sg13g2_dlygate4sd3_1 hold1965 (.A(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .X(net4947));
 sg13g2_dlygate4sd3_1 hold1966 (.A(_00576_),
    .X(net4948));
 sg13g2_dlygate4sd3_1 hold1967 (.A(\i_tinyqv.cpu.data_read_n[1] ),
    .X(net4949));
 sg13g2_dlygate4sd3_1 hold1968 (.A(_00654_),
    .X(net4950));
 sg13g2_dlygate4sd3_1 hold1969 (.A(\i_tinyqv.cpu.data_ready_latch ),
    .X(net4951));
 sg13g2_dlygate4sd3_1 hold1970 (.A(_05449_),
    .X(net4952));
 sg13g2_dlygate4sd3_1 hold1971 (.A(\i_uart_rx.cycle_counter[1] ),
    .X(net4953));
 sg13g2_dlygate4sd3_1 hold1972 (.A(\i2c_config_out[2] ),
    .X(net4954));
 sg13g2_dlygate4sd3_1 hold1973 (.A(_01269_),
    .X(net4955));
 sg13g2_dlygate4sd3_1 hold1974 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .X(net4956));
 sg13g2_dlygate4sd3_1 hold1975 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .X(net4957));
 sg13g2_dlygate4sd3_1 hold1976 (.A(\data_to_write[10] ),
    .X(net4958));
 sg13g2_dlygate4sd3_1 hold1977 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .X(net4959));
 sg13g2_dlygate4sd3_1 hold1978 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .X(net4960));
 sg13g2_dlygate4sd3_1 hold1979 (.A(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .X(net4961));
 sg13g2_dlygate4sd3_1 hold1980 (.A(\data_to_write[14] ),
    .X(net4962));
 sg13g2_dlygate4sd3_1 hold1981 (.A(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .X(net4963));
 sg13g2_dlygate4sd3_1 hold1982 (.A(\crc16_read[3] ),
    .X(net4964));
 sg13g2_dlygate4sd3_1 hold1983 (.A(\gpio_out_sel[3] ),
    .X(net4965));
 sg13g2_dlygate4sd3_1 hold1984 (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .X(net4966));
 sg13g2_dlygate4sd3_1 hold1985 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .X(net4967));
 sg13g2_dlygate4sd3_1 hold1986 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .X(net4968));
 sg13g2_dlygate4sd3_1 hold1987 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .X(net4969));
 sg13g2_dlygate4sd3_1 hold1988 (.A(\timer_count[26] ),
    .X(net4970));
 sg13g2_dlygate4sd3_1 hold1989 (.A(_04506_),
    .X(net4971));
 sg13g2_dlygate4sd3_1 hold1990 (.A(_00443_),
    .X(net4972));
 sg13g2_dlygate4sd3_1 hold1991 (.A(\gpio_out_sel[2] ),
    .X(net4973));
 sg13g2_dlygate4sd3_1 hold1992 (.A(_00364_),
    .X(net4974));
 sg13g2_dlygate4sd3_1 hold1993 (.A(\i_i2c_peri.cmd_start_reg ),
    .X(net4975));
 sg13g2_dlygate4sd3_1 hold1994 (.A(\i_i2c_peri.i_i2c.state_reg[2] ),
    .X(net4976));
 sg13g2_dlygate4sd3_1 hold1995 (.A(_05394_),
    .X(net4977));
 sg13g2_dlygate4sd3_1 hold1996 (.A(_00658_),
    .X(net4978));
 sg13g2_dlygate4sd3_1 hold1997 (.A(\data_to_write[15] ),
    .X(net4979));
 sg13g2_dlygate4sd3_1 hold1998 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .X(net4980));
 sg13g2_dlygate4sd3_1 hold1999 (.A(\crc16_read[10] ),
    .X(net4981));
 sg13g2_dlygate4sd3_1 hold2000 (.A(\data_to_write[9] ),
    .X(net4982));
 sg13g2_dlygate4sd3_1 hold2001 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .X(net4983));
 sg13g2_dlygate4sd3_1 hold2002 (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .X(net4984));
 sg13g2_dlygate4sd3_1 hold2003 (.A(\i_tinyqv.cpu.is_lui ),
    .X(net4985));
 sg13g2_dlygate4sd3_1 hold2004 (.A(\data_to_write[24] ),
    .X(net4986));
 sg13g2_dlygate4sd3_1 hold2005 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .X(net4987));
 sg13g2_dlygate4sd3_1 hold2006 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .X(net4988));
 sg13g2_dlygate4sd3_1 hold2007 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .X(net4989));
 sg13g2_dlygate4sd3_1 hold2008 (.A(\crc16_read[7] ),
    .X(net4990));
 sg13g2_dlygate4sd3_1 hold2009 (.A(_01328_),
    .X(net4991));
 sg13g2_dlygate4sd3_1 hold2010 (.A(\crc16_read[6] ),
    .X(net4992));
 sg13g2_dlygate4sd3_1 hold2011 (.A(_01327_),
    .X(net4993));
 sg13g2_dlygate4sd3_1 hold2012 (.A(\data_to_write[20] ),
    .X(net4994));
 sg13g2_dlygate4sd3_1 hold2013 (.A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .X(net4995));
 sg13g2_dlygate4sd3_1 hold2014 (.A(_00562_),
    .X(net4996));
 sg13g2_dlygate4sd3_1 hold2015 (.A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .X(net4997));
 sg13g2_dlygate4sd3_1 hold2016 (.A(_00561_),
    .X(net4998));
 sg13g2_dlygate4sd3_1 hold2017 (.A(\i_i2c_peri.i_i2c.delay_reg[0] ),
    .X(net4999));
 sg13g2_dlygate4sd3_1 hold2018 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .X(net5000));
 sg13g2_dlygate4sd3_1 hold2019 (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .X(net5001));
 sg13g2_dlygate4sd3_1 hold2020 (.A(\i2c_config_out[11] ),
    .X(net5002));
 sg13g2_dlygate4sd3_1 hold2021 (.A(_01278_),
    .X(net5003));
 sg13g2_dlygate4sd3_1 hold2022 (.A(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .X(net5004));
 sg13g2_dlygate4sd3_1 hold2023 (.A(\data_to_write[30] ),
    .X(net5005));
 sg13g2_dlygate4sd3_1 hold2024 (.A(\i_wdt.counter[20] ),
    .X(net5006));
 sg13g2_dlygate4sd3_1 hold2025 (.A(\i_spi.spi_clk_out ),
    .X(net5007));
 sg13g2_dlygate4sd3_1 hold2026 (.A(\i_tinyqv.cpu.instr_data_in[4] ),
    .X(net5008));
 sg13g2_dlygate4sd3_1 hold2027 (.A(_00491_),
    .X(net5009));
 sg13g2_dlygate4sd3_1 hold2028 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .X(net5010));
 sg13g2_dlygate4sd3_1 hold2029 (.A(\i_wdt.counter[8] ),
    .X(net5011));
 sg13g2_dlygate4sd3_1 hold2030 (.A(\crc_peri_data[2] ),
    .X(net5012));
 sg13g2_dlygate4sd3_1 hold2031 (.A(\crc16_read[5] ),
    .X(net5013));
 sg13g2_dlygate4sd3_1 hold2032 (.A(_01326_),
    .X(net5014));
 sg13g2_dlygate4sd3_1 hold2033 (.A(\crc_peri_data[1] ),
    .X(net5015));
 sg13g2_dlygate4sd3_1 hold2034 (.A(\i_tinyqv.cpu.instr_data_in[6] ),
    .X(net5016));
 sg13g2_dlygate4sd3_1 hold2035 (.A(_00493_),
    .X(net5017));
 sg13g2_dlygate4sd3_1 hold2036 (.A(\timer_count[2] ),
    .X(net5018));
 sg13g2_dlygate4sd3_1 hold2037 (.A(_04431_),
    .X(net5019));
 sg13g2_dlygate4sd3_1 hold2038 (.A(\data_to_write[31] ),
    .X(net5020));
 sg13g2_dlygate4sd3_1 hold2039 (.A(_00888_),
    .X(net5021));
 sg13g2_dlygate4sd3_1 hold2040 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .X(net5022));
 sg13g2_dlygate4sd3_1 hold2041 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .X(net5023));
 sg13g2_dlygate4sd3_1 hold2042 (.A(\i_latch_mem.cycle[1] ),
    .X(net5024));
 sg13g2_dlygate4sd3_1 hold2043 (.A(_01695_),
    .X(net5025));
 sg13g2_dlygate4sd3_1 hold2044 (.A(_01642_),
    .X(net5026));
 sg13g2_dlygate4sd3_1 hold2045 (.A(\i_wdt.counter[18] ),
    .X(net5027));
 sg13g2_dlygate4sd3_1 hold2046 (.A(_00822_),
    .X(net5028));
 sg13g2_dlygate4sd3_1 hold2047 (.A(\i_tinyqv.cpu.is_alu_imm ),
    .X(net5029));
 sg13g2_dlygate4sd3_1 hold2048 (.A(\i_rtc.seconds_out[17] ),
    .X(net5030));
 sg13g2_dlygate4sd3_1 hold2049 (.A(_06338_),
    .X(net5031));
 sg13g2_dlygate4sd3_1 hold2050 (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .X(net5032));
 sg13g2_dlygate4sd3_1 hold2051 (.A(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .X(net5033));
 sg13g2_dlygate4sd3_1 hold2052 (.A(_00526_),
    .X(net5034));
 sg13g2_dlygate4sd3_1 hold2053 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .X(net5035));
 sg13g2_dlygate4sd3_1 hold2054 (.A(\timer_count[13] ),
    .X(net5036));
 sg13g2_dlygate4sd3_1 hold2055 (.A(_04466_),
    .X(net5037));
 sg13g2_dlygate4sd3_1 hold2056 (.A(_00430_),
    .X(net5038));
 sg13g2_dlygate4sd3_1 hold2057 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .X(net5039));
 sg13g2_dlygate4sd3_1 hold2058 (.A(\i_uart_tx.fsm_state[0] ),
    .X(net5040));
 sg13g2_dlygate4sd3_1 hold2059 (.A(_07183_),
    .X(net5041));
 sg13g2_dlygate4sd3_1 hold2060 (.A(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .X(net5042));
 sg13g2_dlygate4sd3_1 hold2061 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .X(net5043));
 sg13g2_dlygate4sd3_1 hold2062 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .X(net5044));
 sg13g2_dlygate4sd3_1 hold2063 (.A(\i_seal.value_reg[0] ),
    .X(net5045));
 sg13g2_dlygate4sd3_1 hold2064 (.A(\i_rtc.seconds_out[30] ),
    .X(net5046));
 sg13g2_dlygate4sd3_1 hold2065 (.A(_06379_),
    .X(net5047));
 sg13g2_dlygate4sd3_1 hold2066 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .X(net5048));
 sg13g2_dlygate4sd3_1 hold2067 (.A(\gpio_out_sel[6] ),
    .X(net5049));
 sg13g2_dlygate4sd3_1 hold2068 (.A(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .X(net5050));
 sg13g2_dlygate4sd3_1 hold2069 (.A(_00726_),
    .X(net5051));
 sg13g2_dlygate4sd3_1 hold2070 (.A(\addr[6] ),
    .X(net5052));
 sg13g2_dlygate4sd3_1 hold2071 (.A(\data_to_write[13] ),
    .X(net5053));
 sg13g2_dlygate4sd3_1 hold2072 (.A(\data_to_write[26] ),
    .X(net5054));
 sg13g2_dlygate4sd3_1 hold2073 (.A(\data_to_write[29] ),
    .X(net5055));
 sg13g2_dlygate4sd3_1 hold2074 (.A(\i_rtc.seconds_out[19] ),
    .X(net5056));
 sg13g2_dlygate4sd3_1 hold2075 (.A(_06343_),
    .X(net5057));
 sg13g2_dlygate4sd3_1 hold2076 (.A(_06345_),
    .X(net5058));
 sg13g2_dlygate4sd3_1 hold2077 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .X(net5059));
 sg13g2_dlygate4sd3_1 hold2078 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .X(net5060));
 sg13g2_dlygate4sd3_1 hold2079 (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .X(net5061));
 sg13g2_dlygate4sd3_1 hold2080 (.A(\i_tinyqv.cpu.is_system ),
    .X(net5062));
 sg13g2_dlygate4sd3_1 hold2081 (.A(\timer_count[5] ),
    .X(net5063));
 sg13g2_dlygate4sd3_1 hold2082 (.A(_04440_),
    .X(net5064));
 sg13g2_dlygate4sd3_1 hold2083 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .X(net5065));
 sg13g2_dlygate4sd3_1 hold2084 (.A(_05845_),
    .X(net5066));
 sg13g2_dlygate4sd3_1 hold2085 (.A(_00740_),
    .X(net5067));
 sg13g2_dlygate4sd3_1 hold2086 (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .X(net5068));
 sg13g2_dlygate4sd3_1 hold2087 (.A(_05830_),
    .X(net5069));
 sg13g2_dlygate4sd3_1 hold2088 (.A(_00732_),
    .X(net5070));
 sg13g2_dlygate4sd3_1 hold2089 (.A(\data_to_write[25] ),
    .X(net5071));
 sg13g2_dlygate4sd3_1 hold2090 (.A(\timer_count[16] ),
    .X(net5072));
 sg13g2_dlygate4sd3_1 hold2091 (.A(\i_tinyqv.cpu.no_write_in_progress ),
    .X(net5073));
 sg13g2_dlygate4sd3_1 hold2092 (.A(\i_tinyqv.cpu.instr_data_in[2] ),
    .X(net5074));
 sg13g2_dlygate4sd3_1 hold2093 (.A(_00489_),
    .X(net5075));
 sg13g2_dlygate4sd3_1 hold2094 (.A(\i_rtc.seconds_out[2] ),
    .X(net5076));
 sg13g2_dlygate4sd3_1 hold2095 (.A(_06289_),
    .X(net5077));
 sg13g2_dlygate4sd3_1 hold2096 (.A(\i2c_config_out[9] ),
    .X(net5078));
 sg13g2_dlygate4sd3_1 hold2097 (.A(\data_to_write[27] ),
    .X(net5079));
 sg13g2_dlygate4sd3_1 hold2098 (.A(_00884_),
    .X(net5080));
 sg13g2_dlygate4sd3_1 hold2099 (.A(\i2c_config_out[10] ),
    .X(net5081));
 sg13g2_dlygate4sd3_1 hold2100 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .X(net5082));
 sg13g2_dlygate4sd3_1 hold2101 (.A(\i_seal.value_reg[5] ),
    .X(net5083));
 sg13g2_dlygate4sd3_1 hold2102 (.A(\i_wdt.counter[4] ),
    .X(net5084));
 sg13g2_dlygate4sd3_1 hold2103 (.A(_06140_),
    .X(net5085));
 sg13g2_dlygate4sd3_1 hold2104 (.A(\i2c_config_out[14] ),
    .X(net5086));
 sg13g2_dlygate4sd3_1 hold2105 (.A(\i_rtc.seconds_out[26] ),
    .X(net5087));
 sg13g2_dlygate4sd3_1 hold2106 (.A(_06366_),
    .X(net5088));
 sg13g2_dlygate4sd3_1 hold2107 (.A(_00883_),
    .X(net5089));
 sg13g2_dlygate4sd3_1 hold2108 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .X(net5090));
 sg13g2_dlygate4sd3_1 hold2109 (.A(_05844_),
    .X(net5091));
 sg13g2_dlygate4sd3_1 hold2110 (.A(_00739_),
    .X(net5092));
 sg13g2_dlygate4sd3_1 hold2111 (.A(\i_i2c_peri.tx_pending ),
    .X(net5093));
 sg13g2_dlygate4sd3_1 hold2112 (.A(_07077_),
    .X(net5094));
 sg13g2_dlygate4sd3_1 hold2113 (.A(\i_seal.value_reg[12] ),
    .X(net5095));
 sg13g2_dlygate4sd3_1 hold2114 (.A(_01068_),
    .X(net5096));
 sg13g2_dlygate4sd3_1 hold2115 (.A(\i_tinyqv.cpu.instr_data_in[5] ),
    .X(net5097));
 sg13g2_dlygate4sd3_1 hold2116 (.A(_00492_),
    .X(net5098));
 sg13g2_dlygate4sd3_1 hold2117 (.A(\crc16_read[9] ),
    .X(net5099));
 sg13g2_dlygate4sd3_1 hold2118 (.A(\i_rtc.seconds_out[21] ),
    .X(net5100));
 sg13g2_dlygate4sd3_1 hold2119 (.A(_06350_),
    .X(net5101));
 sg13g2_dlygate4sd3_1 hold2120 (.A(\i_wdt.counter[13] ),
    .X(net5102));
 sg13g2_dlygate4sd3_1 hold2121 (.A(_06169_),
    .X(net5103));
 sg13g2_dlygate4sd3_1 hold2122 (.A(\data_to_write[11] ),
    .X(net5104));
 sg13g2_dlygate4sd3_1 hold2123 (.A(\i_wdt.counter[10] ),
    .X(net5105));
 sg13g2_dlygate4sd3_1 hold2124 (.A(_06159_),
    .X(net5106));
 sg13g2_dlygate4sd3_1 hold2125 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .X(net5107));
 sg13g2_dlygate4sd3_1 hold2126 (.A(\timer_count[6] ),
    .X(net5108));
 sg13g2_dlygate4sd3_1 hold2127 (.A(_04443_),
    .X(net5109));
 sg13g2_dlygate4sd3_1 hold2128 (.A(\i2c_config_out[8] ),
    .X(net5110));
 sg13g2_dlygate4sd3_1 hold2129 (.A(\i_tinyqv.cpu.instr_fetch_running ),
    .X(net5111));
 sg13g2_dlygate4sd3_1 hold2130 (.A(\i_tinyqv.cpu.is_store ),
    .X(net5112));
 sg13g2_dlygate4sd3_1 hold2131 (.A(\addr[25] ),
    .X(net5113));
 sg13g2_dlygate4sd3_1 hold2132 (.A(\i_rtc.seconds_out[16] ),
    .X(net5114));
 sg13g2_dlygate4sd3_1 hold2133 (.A(_06333_),
    .X(net5115));
 sg13g2_dlygate4sd3_1 hold2134 (.A(_06336_),
    .X(net5116));
 sg13g2_dlygate4sd3_1 hold2135 (.A(\i_wdt.counter[16] ),
    .X(net5117));
 sg13g2_dlygate4sd3_1 hold2136 (.A(\i2c_config_out[13] ),
    .X(net5118));
 sg13g2_dlygate4sd3_1 hold2137 (.A(\i_tinyqv.cpu.is_auipc ),
    .X(net5119));
 sg13g2_dlygate4sd3_1 hold2138 (.A(\i_seal.byte_idx[3] ),
    .X(net5120));
 sg13g2_dlygate4sd3_1 hold2139 (.A(_00894_),
    .X(net5121));
 sg13g2_dlygate4sd3_1 hold2140 (.A(\i_tinyqv.cpu.data_write_n[1] ),
    .X(net5122));
 sg13g2_dlygate4sd3_1 hold2141 (.A(\i_wdt.counter[22] ),
    .X(net5123));
 sg13g2_dlygate4sd3_1 hold2142 (.A(\i_tinyqv.cpu.no_write_in_progress ),
    .X(net5124));
 sg13g2_dlygate4sd3_1 hold2143 (.A(\i_wdt.counter[23] ),
    .X(net5125));
 sg13g2_dlygate4sd3_1 hold2144 (.A(\i2c_config_out[12] ),
    .X(net5126));
 sg13g2_dlygate4sd3_1 hold2145 (.A(_01279_),
    .X(net5127));
 sg13g2_dlygate4sd3_1 hold2146 (.A(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .X(net5128));
 sg13g2_dlygate4sd3_1 hold2147 (.A(\timer_count[10] ),
    .X(net5129));
 sg13g2_dlygate4sd3_1 hold2148 (.A(_04456_),
    .X(net5130));
 sg13g2_dlygate4sd3_1 hold2149 (.A(\timer_count[1] ),
    .X(net5131));
 sg13g2_dlygate4sd3_1 hold2150 (.A(_04427_),
    .X(net5132));
 sg13g2_dlygate4sd3_1 hold2151 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .X(net5133));
 sg13g2_dlygate4sd3_1 hold2152 (.A(\timer_count[23] ),
    .X(net5134));
 sg13g2_dlygate4sd3_1 hold2153 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .X(net5135));
 sg13g2_dlygate4sd3_1 hold2154 (.A(\i_wdt.counter[11] ),
    .X(net5136));
 sg13g2_dlygate4sd3_1 hold2155 (.A(\i_tinyqv.cpu.i_core.mcause[0] ),
    .X(net5137));
 sg13g2_dlygate4sd3_1 hold2156 (.A(_04555_),
    .X(net5138));
 sg13g2_dlygate4sd3_1 hold2157 (.A(\i_i2c_peri.addr_latch[6] ),
    .X(net5139));
 sg13g2_dlygate4sd3_1 hold2158 (.A(\i_rtc.seconds_out[15] ),
    .X(net5140));
 sg13g2_dlygate4sd3_1 hold2159 (.A(_06331_),
    .X(net5141));
 sg13g2_dlygate4sd3_1 hold2160 (.A(\i_tinyqv.cpu.data_write_n[0] ),
    .X(net5142));
 sg13g2_dlygate4sd3_1 hold2161 (.A(\i_wdt.counter[1] ),
    .X(net5143));
 sg13g2_dlygate4sd3_1 hold2162 (.A(_00805_),
    .X(net5144));
 sg13g2_dlygate4sd3_1 hold2163 (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .X(net5145));
 sg13g2_dlygate4sd3_1 hold2164 (.A(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .X(net5146));
 sg13g2_dlygate4sd3_1 hold2165 (.A(\i_i2c_peri.addr_latch[5] ),
    .X(net5147));
 sg13g2_dlygate4sd3_1 hold2166 (.A(\addr[1] ),
    .X(net5148));
 sg13g2_dlygate4sd3_1 hold2167 (.A(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .X(net5149));
 sg13g2_dlygate4sd3_1 hold2168 (.A(\i_rtc.seconds_out[23] ),
    .X(net5150));
 sg13g2_dlygate4sd3_1 hold2169 (.A(_06357_),
    .X(net5151));
 sg13g2_dlygate4sd3_1 hold2170 (.A(\i_wdt.counter[2] ),
    .X(net5152));
 sg13g2_dlygate4sd3_1 hold2171 (.A(_06134_),
    .X(net5153));
 sg13g2_dlygate4sd3_1 hold2172 (.A(\timer_count[12] ),
    .X(net5154));
 sg13g2_dlygate4sd3_1 hold2173 (.A(_00429_),
    .X(net5155));
 sg13g2_dlygate4sd3_1 hold2174 (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .X(net5156));
 sg13g2_dlygate4sd3_1 hold2175 (.A(\i_wdt.counter[15] ),
    .X(net5157));
 sg13g2_dlygate4sd3_1 hold2176 (.A(_06175_),
    .X(net5158));
 sg13g2_dlygate4sd3_1 hold2177 (.A(\i_i2c_peri.i_i2c.phy_state_reg[0] ),
    .X(net5159));
 sg13g2_dlygate4sd3_1 hold2178 (.A(_06985_),
    .X(net5160));
 sg13g2_dlygate4sd3_1 hold2179 (.A(_01238_),
    .X(net5161));
 sg13g2_dlygate4sd3_1 hold2180 (.A(\i_rtc.seconds_out[3] ),
    .X(net5162));
 sg13g2_dlygate4sd3_1 hold2181 (.A(_06292_),
    .X(net5163));
 sg13g2_dlygate4sd3_1 hold2182 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .X(net5164));
 sg13g2_dlygate4sd3_1 hold2183 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .X(net5165));
 sg13g2_dlygate4sd3_1 hold2184 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .X(net5166));
 sg13g2_dlygate4sd3_1 hold2185 (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .X(net5167));
 sg13g2_dlygate4sd3_1 hold2186 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .X(net5168));
 sg13g2_dlygate4sd3_1 hold2187 (.A(\i_i2c_peri.addr_latch[1] ),
    .X(net5169));
 sg13g2_dlygate4sd3_1 hold2188 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .X(net5170));
 sg13g2_dlygate4sd3_1 hold2189 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .X(net5171));
 sg13g2_dlygate4sd3_1 hold2190 (.A(\addr[27] ),
    .X(net5172));
 sg13g2_dlygate4sd3_1 hold2191 (.A(\i_wdt.counter[9] ),
    .X(net5173));
 sg13g2_dlygate4sd3_1 hold2192 (.A(\timer_count[27] ),
    .X(net5174));
 sg13g2_dlygate4sd3_1 hold2193 (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .X(net5175));
 sg13g2_dlygate4sd3_1 hold2194 (.A(\i_rtc.seconds_out[25] ),
    .X(net5176));
 sg13g2_dlygate4sd3_1 hold2195 (.A(_06364_),
    .X(net5177));
 sg13g2_dlygate4sd3_1 hold2196 (.A(\timer_count[14] ),
    .X(net5178));
 sg13g2_dlygate4sd3_1 hold2197 (.A(\i_rtc.seconds_out[4] ),
    .X(net5179));
 sg13g2_dlygate4sd3_1 hold2198 (.A(\i_rtc.seconds_out[18] ),
    .X(net5180));
 sg13g2_dlygate4sd3_1 hold2199 (.A(\i_rtc.seconds_out[11] ),
    .X(net5181));
 sg13g2_dlygate4sd3_1 hold2200 (.A(_06317_),
    .X(net5182));
 sg13g2_dlygate4sd3_1 hold2201 (.A(_00868_),
    .X(net5183));
 sg13g2_dlygate4sd3_1 hold2202 (.A(\i_i2c_peri.i_i2c.state_reg[3] ),
    .X(net5184));
 sg13g2_dlygate4sd3_1 hold2203 (.A(\i_tinyqv.cpu.is_alu_reg ),
    .X(net5185));
 sg13g2_dlygate4sd3_1 hold2204 (.A(\timer_count[25] ),
    .X(net5186));
 sg13g2_dlygate4sd3_1 hold2205 (.A(_04504_),
    .X(net5187));
 sg13g2_dlygate4sd3_1 hold2206 (.A(\i_i2c_peri.addr_latch[0] ),
    .X(net5188));
 sg13g2_dlygate4sd3_1 hold2207 (.A(\i_tinyqv.cpu.alu_op[3] ),
    .X(net5189));
 sg13g2_dlygate4sd3_1 hold2208 (.A(\i_seal.byte_idx[2] ),
    .X(net5190));
 sg13g2_dlygate4sd3_1 hold2209 (.A(_06406_),
    .X(net5191));
 sg13g2_dlygate4sd3_1 hold2210 (.A(\i_tinyqv.cpu.instr_data_start[23] ),
    .X(net5192));
 sg13g2_dlygate4sd3_1 hold2211 (.A(\i_rtc.seconds_out[22] ),
    .X(net5193));
 sg13g2_dlygate4sd3_1 hold2212 (.A(_06352_),
    .X(net5194));
 sg13g2_dlygate4sd3_1 hold2213 (.A(_06355_),
    .X(net5195));
 sg13g2_dlygate4sd3_1 hold2214 (.A(\addr[26] ),
    .X(net5196));
 sg13g2_dlygate4sd3_1 hold2215 (.A(\i_rtc.seconds_out[8] ),
    .X(net5197));
 sg13g2_dlygate4sd3_1 hold2216 (.A(_06306_),
    .X(net5198));
 sg13g2_dlygate4sd3_1 hold2217 (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(net5199));
 sg13g2_dlygate4sd3_1 hold2218 (.A(\i_i2c_peri.addr_latch[3] ),
    .X(net5200));
 sg13g2_dlygate4sd3_1 hold2219 (.A(\i_seal.state[1] ),
    .X(net5201));
 sg13g2_dlygate4sd3_1 hold2220 (.A(_06413_),
    .X(net5202));
 sg13g2_dlygate4sd3_1 hold2221 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .X(net5203));
 sg13g2_dlygate4sd3_1 hold2222 (.A(\i_tinyqv.cpu.i_core.load_top_bit ),
    .X(net5204));
 sg13g2_dlygate4sd3_1 hold2223 (.A(_04260_),
    .X(net5205));
 sg13g2_dlygate4sd3_1 hold2224 (.A(\i_i2c_peri.addr_latch[2] ),
    .X(net5206));
 sg13g2_dlygate4sd3_1 hold2225 (.A(\timer_count[28] ),
    .X(net5207));
 sg13g2_dlygate4sd3_1 hold2226 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .X(net5208));
 sg13g2_dlygate4sd3_1 hold2227 (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .X(net5209));
 sg13g2_dlygate4sd3_1 hold2228 (.A(\i_wdt.counter[14] ),
    .X(net5210));
 sg13g2_dlygate4sd3_1 hold2229 (.A(_04289_),
    .X(net5211));
 sg13g2_dlygate4sd3_1 hold2230 (.A(_00818_),
    .X(net5212));
 sg13g2_dlygate4sd3_1 hold2231 (.A(\i_rtc.seconds_out[20] ),
    .X(net5213));
 sg13g2_dlygate4sd3_1 hold2232 (.A(\i_tinyqv.cpu.is_jalr ),
    .X(net5214));
 sg13g2_dlygate4sd3_1 hold2233 (.A(\i_wdt.counter[29] ),
    .X(net5215));
 sg13g2_dlygate4sd3_1 hold2234 (.A(_04326_),
    .X(net5216));
 sg13g2_dlygate4sd3_1 hold2235 (.A(_00378_),
    .X(net5217));
 sg13g2_dlygate4sd3_1 hold2236 (.A(\timer_count[8] ),
    .X(net5218));
 sg13g2_dlygate4sd3_1 hold2237 (.A(_04447_),
    .X(net5219));
 sg13g2_dlygate4sd3_1 hold2238 (.A(_04449_),
    .X(net5220));
 sg13g2_dlygate4sd3_1 hold2239 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .X(net5221));
 sg13g2_dlygate4sd3_1 hold2240 (.A(\i_rtc.seconds_out[29] ),
    .X(net5222));
 sg13g2_dlygate4sd3_1 hold2241 (.A(_06376_),
    .X(net5223));
 sg13g2_dlygate4sd3_1 hold2242 (.A(_06377_),
    .X(net5224));
 sg13g2_dlygate4sd3_1 hold2243 (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .X(net5225));
 sg13g2_dlygate4sd3_1 hold2244 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .X(net5226));
 sg13g2_dlygate4sd3_1 hold2245 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .X(net5227));
 sg13g2_dlygate4sd3_1 hold2246 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .X(net5228));
 sg13g2_dlygate4sd3_1 hold2247 (.A(\timer_count[7] ),
    .X(net5229));
 sg13g2_dlygate4sd3_1 hold2248 (.A(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .X(net5230));
 sg13g2_dlygate4sd3_1 hold2249 (.A(\i_rtc.seconds_out[10] ),
    .X(net5231));
 sg13g2_dlygate4sd3_1 hold2250 (.A(_06312_),
    .X(net5232));
 sg13g2_dlygate4sd3_1 hold2251 (.A(_00867_),
    .X(net5233));
 sg13g2_dlygate4sd3_1 hold2252 (.A(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .X(net5234));
 sg13g2_dlygate4sd3_1 hold2253 (.A(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .X(net5235));
 sg13g2_dlygate4sd3_1 hold2254 (.A(\i_uart_rx.fsm_state[3] ),
    .X(net5236));
 sg13g2_dlygate4sd3_1 hold2255 (.A(_01662_),
    .X(net5237));
 sg13g2_dlygate4sd3_1 hold2256 (.A(_01374_),
    .X(net5238));
 sg13g2_dlygate4sd3_1 hold2257 (.A(\i_rtc.seconds_out[13] ),
    .X(net5239));
 sg13g2_dlygate4sd3_1 hold2258 (.A(_06323_),
    .X(net5240));
 sg13g2_dlygate4sd3_1 hold2259 (.A(_06326_),
    .X(net5241));
 sg13g2_dlygate4sd3_1 hold2260 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .X(net5242));
 sg13g2_dlygate4sd3_1 hold2261 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .X(net5243));
 sg13g2_dlygate4sd3_1 hold2262 (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(net5244));
 sg13g2_dlygate4sd3_1 hold2263 (.A(\i_rtc.seconds_out[14] ),
    .X(net5245));
 sg13g2_dlygate4sd3_1 hold2264 (.A(_06327_),
    .X(net5246));
 sg13g2_dlygate4sd3_1 hold2265 (.A(\addr[0] ),
    .X(net5247));
 sg13g2_dlygate4sd3_1 hold2266 (.A(_01153_),
    .X(net5248));
 sg13g2_dlygate4sd3_1 hold2267 (.A(\i_tinyqv.cpu.instr_data_start[15] ),
    .X(net5249));
 sg13g2_dlygate4sd3_1 hold2268 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .X(net5250));
 sg13g2_dlygate4sd3_1 hold2269 (.A(\timer_count[3] ),
    .X(net5251));
 sg13g2_dlygate4sd3_1 hold2270 (.A(_04432_),
    .X(net5252));
 sg13g2_dlygate4sd3_1 hold2271 (.A(\i_spi.busy ),
    .X(net5253));
 sg13g2_dlygate4sd3_1 hold2272 (.A(\i_tinyqv.cpu.instr_data_in[7] ),
    .X(net5254));
 sg13g2_dlygate4sd3_1 hold2273 (.A(_00494_),
    .X(net5255));
 sg13g2_dlygate4sd3_1 hold2274 (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .X(net5256));
 sg13g2_dlygate4sd3_1 hold2275 (.A(\i_i2c_peri.i_i2c.bit_count_reg[0] ),
    .X(net5257));
 sg13g2_dlygate4sd3_1 hold2276 (.A(\i_rtc.seconds_out[5] ),
    .X(net5258));
 sg13g2_dlygate4sd3_1 hold2277 (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .X(net5259));
 sg13g2_dlygate4sd3_1 hold2278 (.A(\i_tinyqv.cpu.pc[2] ),
    .X(net5260));
 sg13g2_dlygate4sd3_1 hold2279 (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .X(net5261));
 sg13g2_dlygate4sd3_1 hold2280 (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(net5262));
 sg13g2_dlygate4sd3_1 hold2281 (.A(\addr[5] ),
    .X(net5263));
 sg13g2_dlygate4sd3_1 hold2282 (.A(_01158_),
    .X(net5264));
 sg13g2_dlygate4sd3_1 hold2283 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .X(net5265));
 sg13g2_dlygate4sd3_1 hold2284 (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .X(net5266));
 sg13g2_dlygate4sd3_1 hold2285 (.A(_04948_),
    .X(net5267));
 sg13g2_dlygate4sd3_1 hold2286 (.A(_00549_),
    .X(net5268));
 sg13g2_dlygate4sd3_1 hold2287 (.A(\i_tinyqv.cpu.instr_fetch_started ),
    .X(net5269));
 sg13g2_dlygate4sd3_1 hold2288 (.A(_05274_),
    .X(net5270));
 sg13g2_dlygate4sd3_1 hold2289 (.A(_05275_),
    .X(net5271));
 sg13g2_dlygate4sd3_1 hold2290 (.A(\i_tinyqv.cpu.instr_data_in[11] ),
    .X(net5272));
 sg13g2_dlygate4sd3_1 hold2291 (.A(_00548_),
    .X(net5273));
 sg13g2_dlygate4sd3_1 hold2292 (.A(\i_tinyqv.cpu.alu_op[2] ),
    .X(net5274));
 sg13g2_dlygate4sd3_1 hold2293 (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(net5275));
 sg13g2_dlygate4sd3_1 hold2294 (.A(\i_rtc.seconds_out[28] ),
    .X(net5276));
 sg13g2_dlygate4sd3_1 hold2295 (.A(_06371_),
    .X(net5277));
 sg13g2_dlygate4sd3_1 hold2296 (.A(_06373_),
    .X(net5278));
 sg13g2_dlygate4sd3_1 hold2297 (.A(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .X(net5279));
 sg13g2_dlygate4sd3_1 hold2298 (.A(\timer_count[21] ),
    .X(net5280));
 sg13g2_dlygate4sd3_1 hold2299 (.A(\i_wdt.counter[28] ),
    .X(net5281));
 sg13g2_dlygate4sd3_1 hold2300 (.A(\i_tinyqv.mem.q_ctrl.is_writing ),
    .X(net5282));
 sg13g2_dlygate4sd3_1 hold2301 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .X(net5283));
 sg13g2_dlygate4sd3_1 hold2302 (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .X(net5284));
 sg13g2_dlygate4sd3_1 hold2303 (.A(\i_tinyqv.cpu.pc[1] ),
    .X(net5285));
 sg13g2_dlygate4sd3_1 hold2304 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(net5286));
 sg13g2_dlygate4sd3_1 hold2305 (.A(\timer_count[24] ),
    .X(net5287));
 sg13g2_dlygate4sd3_1 hold2306 (.A(\i_rtc.seconds_out[9] ),
    .X(net5288));
 sg13g2_dlygate4sd3_1 hold2307 (.A(_06309_),
    .X(net5289));
 sg13g2_dlygate4sd3_1 hold2308 (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .X(net5290));
 sg13g2_dlygate4sd3_1 hold2309 (.A(\i_wdt.counter[0] ),
    .X(net5291));
 sg13g2_dlygate4sd3_1 hold2310 (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .X(net5292));
 sg13g2_dlygate4sd3_1 hold2311 (.A(\i_rtc.seconds_out[12] ),
    .X(net5293));
 sg13g2_dlygate4sd3_1 hold2312 (.A(_00869_),
    .X(net5294));
 sg13g2_dlygate4sd3_1 hold2313 (.A(\i_uart_tx.data_to_send[1] ),
    .X(net5295));
 sg13g2_dlygate4sd3_1 hold2314 (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .X(net5296));
 sg13g2_dlygate4sd3_1 hold2315 (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .X(net5297));
 sg13g2_dlygate4sd3_1 hold2316 (.A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .X(net5298));
 sg13g2_dlygate4sd3_1 hold2317 (.A(\i_seal.byte_idx[1] ),
    .X(net5299));
 sg13g2_dlygate4sd3_1 hold2318 (.A(_06404_),
    .X(net5300));
 sg13g2_dlygate4sd3_1 hold2319 (.A(\i_uart_tx.data_to_send[3] ),
    .X(net5301));
 sg13g2_dlygate4sd3_1 hold2320 (.A(_07147_),
    .X(net5302));
 sg13g2_dlygate4sd3_1 hold2321 (.A(\i_i2c_peri.i_i2c.bit_count_reg[1] ),
    .X(net5303));
 sg13g2_dlygate4sd3_1 hold2322 (.A(\i_wdt.counter[12] ),
    .X(net5304));
 sg13g2_dlygate4sd3_1 hold2323 (.A(\i_uart_tx.data_to_send[2] ),
    .X(net5305));
 sg13g2_dlygate4sd3_1 hold2324 (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .X(net5306));
 sg13g2_dlygate4sd3_1 hold2325 (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .X(net5307));
 sg13g2_dlygate4sd3_1 hold2326 (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(net5308));
 sg13g2_dlygate4sd3_1 hold2327 (.A(\i_rtc.seconds_out[6] ),
    .X(net5309));
 sg13g2_dlygate4sd3_1 hold2328 (.A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .X(net5310));
 sg13g2_dlygate4sd3_1 hold2329 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .X(net5311));
 sg13g2_dlygate4sd3_1 hold2330 (.A(\i_latch_mem.cycle[0] ),
    .X(net5312));
 sg13g2_dlygate4sd3_1 hold2331 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .X(net5313));
 sg13g2_dlygate4sd3_1 hold2332 (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .X(net5314));
 sg13g2_dlygate4sd3_1 hold2333 (.A(_00569_),
    .X(net5315));
 sg13g2_dlygate4sd3_1 hold2334 (.A(\addr[2] ),
    .X(net5316));
 sg13g2_dlygate4sd3_1 hold2335 (.A(\i_wdt.counter[6] ),
    .X(net5317));
 sg13g2_dlygate4sd3_1 hold2336 (.A(\timer_count[31] ),
    .X(net5318));
 sg13g2_dlygate4sd3_1 hold2337 (.A(_04528_),
    .X(net5319));
 sg13g2_dlygate4sd3_1 hold2338 (.A(\i_rtc.seconds_out[1] ),
    .X(net5320));
 sg13g2_dlygate4sd3_1 hold2339 (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .X(net5321));
 sg13g2_dlygate4sd3_1 hold2340 (.A(\timer_count[29] ),
    .X(net5322));
 sg13g2_dlygate4sd3_1 hold2341 (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .X(net5323));
 sg13g2_dlygate4sd3_1 hold2342 (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .X(net5324));
 sg13g2_dlygate4sd3_1 hold2343 (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .X(net5325));
 sg13g2_dlygate4sd3_1 hold2344 (.A(\i_tinyqv.cpu.is_load ),
    .X(net5326));
 sg13g2_dlygate4sd3_1 hold2345 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .X(net5327));
 sg13g2_dlygate4sd3_1 hold2346 (.A(_04849_),
    .X(net5328));
 sg13g2_dlygate4sd3_1 hold2347 (.A(\timer_count[30] ),
    .X(net5329));
 sg13g2_dlygate4sd3_1 hold2348 (.A(\timer_count[4] ),
    .X(net5330));
 sg13g2_dlygate4sd3_1 hold2349 (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .X(net5331));
 sg13g2_dlygate4sd3_1 hold2350 (.A(\i_rtc.seconds_out[7] ),
    .X(net5332));
 sg13g2_dlygate4sd3_1 hold2351 (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .X(net5333));
 sg13g2_dlygate4sd3_1 hold2352 (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .X(net5334));
 sg13g2_dlygate4sd3_1 hold2353 (.A(\i_uart_rx.fsm_state[0] ),
    .X(net5335));
 sg13g2_dlygate4sd3_1 hold2354 (.A(_07228_),
    .X(net5336));
 sg13g2_dlygate4sd3_1 hold2355 (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .X(net5337));
 sg13g2_dlygate4sd3_1 hold2356 (.A(debug_instr_valid),
    .X(net5338));
 sg13g2_dlygate4sd3_1 hold2357 (.A(\i_uart_rx.fsm_state[1] ),
    .X(net5339));
 sg13g2_dlygate4sd3_1 hold2358 (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .X(net5340));
 sg13g2_dlygate4sd3_1 hold2359 (.A(_00567_),
    .X(net5341));
 sg13g2_dlygate4sd3_1 hold2360 (.A(\timer_count[0] ),
    .X(net5342));
 sg13g2_dlygate4sd3_1 hold2361 (.A(\i_tinyqv.cpu.instr_data_in[15] ),
    .X(net5343));
 sg13g2_dlygate4sd3_1 hold2362 (.A(_00552_),
    .X(net5344));
 sg13g2_dlygate4sd3_1 hold2363 (.A(\i_seal.state[0] ),
    .X(net5345));
 sg13g2_dlygate4sd3_1 hold2364 (.A(_06399_),
    .X(net5346));
 sg13g2_dlygate4sd3_1 hold2365 (.A(_06400_),
    .X(net5347));
 sg13g2_dlygate4sd3_1 hold2366 (.A(\i_i2c_peri.i_i2c.mode_stop_reg ),
    .X(net5348));
 sg13g2_dlygate4sd3_1 hold2367 (.A(\i_i2c_peri.i_i2c.phy_state_reg[3] ),
    .X(net5349));
 sg13g2_dlygate4sd3_1 hold2368 (.A(_06997_),
    .X(net5350));
 sg13g2_dlygate4sd3_1 hold2369 (.A(_01241_),
    .X(net5351));
 sg13g2_dlygate4sd3_1 hold2370 (.A(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .X(net5352));
 sg13g2_dlygate4sd3_1 hold2371 (.A(\timer_count[9] ),
    .X(net5353));
 sg13g2_dlygate4sd3_1 hold2372 (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .X(net5354));
 sg13g2_dlygate4sd3_1 hold2373 (.A(\i_tinyqv.cpu.instr_write_offset[1] ),
    .X(net5355));
 sg13g2_dlygate4sd3_1 hold2374 (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .X(net5356));
 sg13g2_dlygate4sd3_1 hold2375 (.A(\i_i2c_peri.i_i2c.delay_scl_reg ),
    .X(net5357));
 sg13g2_dlygate4sd3_1 hold2376 (.A(\i_i2c_peri.i_i2c.state_reg[0] ),
    .X(net5358));
 sg13g2_dlygate4sd3_1 hold2377 (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .X(net5359));
 sg13g2_dlygate4sd3_1 hold2378 (.A(\i_tinyqv.cpu.counter[2] ),
    .X(net5360));
 sg13g2_dlygate4sd3_1 hold2379 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .X(net5361));
 sg13g2_dlygate4sd3_1 hold2380 (.A(\i_rtc.seconds_out[0] ),
    .X(net5362));
 sg13g2_dlygate4sd3_1 hold2381 (.A(\i_tinyqv.cpu.instr_data_in[14] ),
    .X(net5363));
 sg13g2_dlygate4sd3_1 hold2382 (.A(_00551_),
    .X(net5364));
 sg13g2_dlygate4sd3_1 hold2383 (.A(\i_i2c_peri.i_i2c.s_axis_data_tready_reg ),
    .X(net5365));
 sg13g2_dlygate4sd3_1 hold2384 (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .X(net5366));
 sg13g2_dlygate4sd3_1 hold2385 (.A(_00550_),
    .X(net5367));
 sg13g2_dlygate4sd3_1 hold2386 (.A(\addr[3] ),
    .X(net5368));
 sg13g2_dlygate4sd3_1 hold2387 (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .X(net5369));
 sg13g2_dlygate4sd3_1 hold2388 (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(net5370));
 sg13g2_dlygate4sd3_1 hold2389 (.A(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .X(net5371));
 sg13g2_dlygate4sd3_1 hold2390 (.A(\i_i2c_peri.i_i2c.phy_state_reg[0] ),
    .X(net5372));
 sg13g2_dlygate4sd3_1 hold2391 (.A(\data_to_write[12] ),
    .X(net5373));
 sg13g2_dlygate4sd3_1 hold2392 (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .X(net5374));
 sg13g2_dlygate4sd3_1 hold2393 (.A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .X(net5375));
 sg13g2_dlygate4sd3_1 hold2394 (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .X(net5376));
 sg13g2_dlygate4sd3_1 hold2395 (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .X(net5377));
 sg13g2_dlygate4sd3_1 hold2396 (.A(\i_i2c_peri.i_i2c.phy_state_reg[2] ),
    .X(net5378));
 sg13g2_dlygate4sd3_1 hold2397 (.A(\i_tinyqv.cpu.alu_op[0] ),
    .X(net5379));
 sg13g2_dlygate4sd3_1 hold2398 (.A(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .X(net5380));
 sg13g2_dlygate4sd3_1 hold2399 (.A(\us_divider[4] ),
    .X(net5381));
 sg13g2_dlygate4sd3_1 hold2400 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .X(net5382));
 sg13g2_dlygate4sd3_1 hold2401 (.A(_04031_),
    .X(net5383));
 sg13g2_dlygate4sd3_1 hold2402 (.A(\i_wdt.counter[15] ),
    .X(net5384));
 sg13g2_dlygate4sd3_1 hold2403 (.A(\i_uart_rx.cycle_counter[5] ),
    .X(net5385));
 sg13g2_dlygate4sd3_1 hold2404 (.A(\i_rtc.us_count[11] ),
    .X(net5386));
 sg13g2_dlygate4sd3_1 hold2405 (.A(\timer_count[12] ),
    .X(net5387));
 sg13g2_dlygate4sd3_1 hold2406 (.A(\timer_count[0] ),
    .X(net5388));
 sg13g2_decap_4 FILLER_0_0 ();
 sg13g2_fill_2 FILLER_0_4 ();
 sg13g2_decap_8 FILLER_0_33 ();
 sg13g2_decap_8 FILLER_0_40 ();
 sg13g2_decap_4 FILLER_0_47 ();
 sg13g2_fill_1 FILLER_0_51 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_fill_2 FILLER_0_75 ();
 sg13g2_decap_8 FILLER_0_87 ();
 sg13g2_fill_2 FILLER_0_94 ();
 sg13g2_fill_1 FILLER_0_96 ();
 sg13g2_decap_4 FILLER_0_118 ();
 sg13g2_decap_4 FILLER_0_139 ();
 sg13g2_fill_1 FILLER_0_143 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_fill_2 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_fill_2 FILLER_0_203 ();
 sg13g2_fill_1 FILLER_0_205 ();
 sg13g2_fill_2 FILLER_0_209 ();
 sg13g2_fill_1 FILLER_0_211 ();
 sg13g2_decap_4 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_4 FILLER_0_266 ();
 sg13g2_fill_1 FILLER_0_270 ();
 sg13g2_fill_2 FILLER_0_299 ();
 sg13g2_fill_2 FILLER_0_369 ();
 sg13g2_fill_1 FILLER_0_371 ();
 sg13g2_fill_2 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_447 ();
 sg13g2_decap_8 FILLER_0_454 ();
 sg13g2_fill_1 FILLER_0_461 ();
 sg13g2_decap_4 FILLER_0_489 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_4 FILLER_0_511 ();
 sg13g2_fill_1 FILLER_0_515 ();
 sg13g2_decap_8 FILLER_0_544 ();
 sg13g2_fill_1 FILLER_0_551 ();
 sg13g2_fill_2 FILLER_0_580 ();
 sg13g2_fill_1 FILLER_0_582 ();
 sg13g2_decap_4 FILLER_0_611 ();
 sg13g2_fill_1 FILLER_0_615 ();
 sg13g2_fill_2 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_676 ();
 sg13g2_fill_1 FILLER_0_683 ();
 sg13g2_fill_2 FILLER_0_720 ();
 sg13g2_fill_1 FILLER_0_722 ();
 sg13g2_decap_8 FILLER_0_879 ();
 sg13g2_fill_2 FILLER_0_1041 ();
 sg13g2_fill_2 FILLER_0_1083 ();
 sg13g2_fill_1 FILLER_0_1157 ();
 sg13g2_fill_2 FILLER_0_1225 ();
 sg13g2_fill_1 FILLER_0_1227 ();
 sg13g2_fill_1 FILLER_0_1255 ();
 sg13g2_fill_2 FILLER_0_1304 ();
 sg13g2_fill_2 FILLER_0_1319 ();
 sg13g2_fill_2 FILLER_0_1357 ();
 sg13g2_fill_2 FILLER_0_1399 ();
 sg13g2_fill_1 FILLER_0_1401 ();
 sg13g2_fill_1 FILLER_0_1501 ();
 sg13g2_fill_2 FILLER_0_1538 ();
 sg13g2_fill_2 FILLER_0_1567 ();
 sg13g2_fill_2 FILLER_0_1617 ();
 sg13g2_fill_1 FILLER_0_1619 ();
 sg13g2_fill_2 FILLER_0_1633 ();
 sg13g2_fill_1 FILLER_0_1635 ();
 sg13g2_fill_2 FILLER_0_1680 ();
 sg13g2_fill_1 FILLER_0_1682 ();
 sg13g2_decap_8 FILLER_0_1716 ();
 sg13g2_decap_8 FILLER_0_1723 ();
 sg13g2_decap_8 FILLER_0_1730 ();
 sg13g2_decap_8 FILLER_0_1737 ();
 sg13g2_decap_8 FILLER_0_1744 ();
 sg13g2_decap_8 FILLER_0_1751 ();
 sg13g2_decap_8 FILLER_0_1758 ();
 sg13g2_fill_2 FILLER_0_1765 ();
 sg13g2_fill_1 FILLER_0_1767 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_fill_2 FILLER_1_14 ();
 sg13g2_fill_1 FILLER_1_16 ();
 sg13g2_decap_4 FILLER_1_152 ();
 sg13g2_fill_1 FILLER_1_156 ();
 sg13g2_decap_4 FILLER_1_161 ();
 sg13g2_fill_1 FILLER_1_170 ();
 sg13g2_fill_1 FILLER_1_226 ();
 sg13g2_decap_4 FILLER_1_230 ();
 sg13g2_fill_2 FILLER_1_242 ();
 sg13g2_fill_2 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_4 FILLER_1_294 ();
 sg13g2_fill_2 FILLER_1_345 ();
 sg13g2_fill_2 FILLER_1_374 ();
 sg13g2_fill_1 FILLER_1_404 ();
 sg13g2_fill_2 FILLER_1_409 ();
 sg13g2_decap_8 FILLER_1_415 ();
 sg13g2_decap_8 FILLER_1_422 ();
 sg13g2_fill_2 FILLER_1_429 ();
 sg13g2_fill_1 FILLER_1_431 ();
 sg13g2_fill_2 FILLER_1_477 ();
 sg13g2_fill_1 FILLER_1_526 ();
 sg13g2_fill_2 FILLER_1_531 ();
 sg13g2_fill_1 FILLER_1_533 ();
 sg13g2_decap_8 FILLER_1_548 ();
 sg13g2_fill_2 FILLER_1_555 ();
 sg13g2_decap_4 FILLER_1_561 ();
 sg13g2_fill_2 FILLER_1_565 ();
 sg13g2_decap_8 FILLER_1_572 ();
 sg13g2_fill_1 FILLER_1_579 ();
 sg13g2_decap_8 FILLER_1_594 ();
 sg13g2_decap_4 FILLER_1_605 ();
 sg13g2_fill_1 FILLER_1_609 ();
 sg13g2_fill_2 FILLER_1_619 ();
 sg13g2_decap_4 FILLER_1_625 ();
 sg13g2_fill_1 FILLER_1_629 ();
 sg13g2_fill_2 FILLER_1_659 ();
 sg13g2_decap_8 FILLER_1_687 ();
 sg13g2_fill_1 FILLER_1_694 ();
 sg13g2_fill_2 FILLER_1_704 ();
 sg13g2_decap_4 FILLER_1_753 ();
 sg13g2_fill_1 FILLER_1_819 ();
 sg13g2_fill_1 FILLER_1_927 ();
 sg13g2_fill_2 FILLER_1_986 ();
 sg13g2_fill_1 FILLER_1_988 ();
 sg13g2_fill_2 FILLER_1_1024 ();
 sg13g2_fill_2 FILLER_1_1116 ();
 sg13g2_fill_1 FILLER_1_1207 ();
 sg13g2_fill_1 FILLER_1_1377 ();
 sg13g2_fill_2 FILLER_1_1481 ();
 sg13g2_fill_2 FILLER_1_1590 ();
 sg13g2_fill_1 FILLER_1_1592 ();
 sg13g2_decap_8 FILLER_1_1727 ();
 sg13g2_decap_8 FILLER_1_1734 ();
 sg13g2_decap_8 FILLER_1_1741 ();
 sg13g2_decap_8 FILLER_1_1748 ();
 sg13g2_decap_8 FILLER_1_1755 ();
 sg13g2_decap_4 FILLER_1_1762 ();
 sg13g2_fill_2 FILLER_1_1766 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_16 ();
 sg13g2_fill_2 FILLER_2_23 ();
 sg13g2_fill_2 FILLER_2_29 ();
 sg13g2_fill_1 FILLER_2_51 ();
 sg13g2_fill_1 FILLER_2_57 ();
 sg13g2_decap_4 FILLER_2_66 ();
 sg13g2_fill_2 FILLER_2_88 ();
 sg13g2_decap_4 FILLER_2_102 ();
 sg13g2_fill_1 FILLER_2_106 ();
 sg13g2_fill_1 FILLER_2_112 ();
 sg13g2_fill_1 FILLER_2_131 ();
 sg13g2_decap_4 FILLER_2_140 ();
 sg13g2_fill_1 FILLER_2_153 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_decap_4 FILLER_2_198 ();
 sg13g2_fill_2 FILLER_2_202 ();
 sg13g2_decap_4 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_252 ();
 sg13g2_decap_4 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_fill_2 FILLER_2_291 ();
 sg13g2_fill_1 FILLER_2_293 ();
 sg13g2_decap_4 FILLER_2_298 ();
 sg13g2_fill_1 FILLER_2_302 ();
 sg13g2_fill_2 FILLER_2_322 ();
 sg13g2_fill_1 FILLER_2_324 ();
 sg13g2_fill_1 FILLER_2_351 ();
 sg13g2_fill_1 FILLER_2_398 ();
 sg13g2_decap_4 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_431 ();
 sg13g2_decap_4 FILLER_2_457 ();
 sg13g2_fill_1 FILLER_2_493 ();
 sg13g2_fill_2 FILLER_2_519 ();
 sg13g2_fill_1 FILLER_2_521 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_fill_1 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_583 ();
 sg13g2_decap_8 FILLER_2_590 ();
 sg13g2_decap_4 FILLER_2_597 ();
 sg13g2_fill_2 FILLER_2_601 ();
 sg13g2_decap_8 FILLER_2_628 ();
 sg13g2_decap_4 FILLER_2_635 ();
 sg13g2_fill_2 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_4 FILLER_2_686 ();
 sg13g2_fill_1 FILLER_2_690 ();
 sg13g2_fill_2 FILLER_2_759 ();
 sg13g2_fill_1 FILLER_2_761 ();
 sg13g2_fill_2 FILLER_2_774 ();
 sg13g2_fill_1 FILLER_2_875 ();
 sg13g2_fill_1 FILLER_2_992 ();
 sg13g2_fill_2 FILLER_2_1038 ();
 sg13g2_fill_1 FILLER_2_1040 ();
 sg13g2_fill_1 FILLER_2_1054 ();
 sg13g2_fill_2 FILLER_2_1149 ();
 sg13g2_fill_1 FILLER_2_1151 ();
 sg13g2_fill_2 FILLER_2_1182 ();
 sg13g2_fill_1 FILLER_2_1358 ();
 sg13g2_fill_1 FILLER_2_1368 ();
 sg13g2_fill_2 FILLER_2_1409 ();
 sg13g2_fill_2 FILLER_2_1424 ();
 sg13g2_fill_1 FILLER_2_1426 ();
 sg13g2_fill_2 FILLER_2_1454 ();
 sg13g2_fill_2 FILLER_2_1509 ();
 sg13g2_fill_1 FILLER_2_1511 ();
 sg13g2_fill_2 FILLER_2_1559 ();
 sg13g2_fill_1 FILLER_2_1561 ();
 sg13g2_fill_1 FILLER_2_1611 ();
 sg13g2_fill_2 FILLER_2_1625 ();
 sg13g2_fill_1 FILLER_2_1627 ();
 sg13g2_fill_2 FILLER_2_1686 ();
 sg13g2_fill_2 FILLER_2_1701 ();
 sg13g2_decap_8 FILLER_2_1735 ();
 sg13g2_decap_8 FILLER_2_1742 ();
 sg13g2_decap_8 FILLER_2_1749 ();
 sg13g2_decap_8 FILLER_2_1756 ();
 sg13g2_decap_4 FILLER_2_1763 ();
 sg13g2_fill_1 FILLER_2_1767 ();
 sg13g2_decap_4 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_4 ();
 sg13g2_fill_2 FILLER_3_14 ();
 sg13g2_fill_1 FILLER_3_16 ();
 sg13g2_fill_2 FILLER_3_30 ();
 sg13g2_fill_1 FILLER_3_32 ();
 sg13g2_fill_1 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_55 ();
 sg13g2_fill_2 FILLER_3_62 ();
 sg13g2_fill_1 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_141 ();
 sg13g2_fill_2 FILLER_3_166 ();
 sg13g2_fill_1 FILLER_3_168 ();
 sg13g2_decap_4 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_199 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_fill_1 FILLER_3_213 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_fill_2 FILLER_3_233 ();
 sg13g2_fill_1 FILLER_3_247 ();
 sg13g2_fill_2 FILLER_3_268 ();
 sg13g2_fill_1 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_fill_1 FILLER_3_287 ();
 sg13g2_fill_2 FILLER_3_316 ();
 sg13g2_fill_2 FILLER_3_387 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_412 ();
 sg13g2_decap_8 FILLER_3_426 ();
 sg13g2_fill_2 FILLER_3_437 ();
 sg13g2_fill_2 FILLER_3_460 ();
 sg13g2_decap_4 FILLER_3_471 ();
 sg13g2_fill_2 FILLER_3_488 ();
 sg13g2_fill_1 FILLER_3_495 ();
 sg13g2_fill_1 FILLER_3_501 ();
 sg13g2_decap_4 FILLER_3_510 ();
 sg13g2_fill_2 FILLER_3_528 ();
 sg13g2_fill_1 FILLER_3_530 ();
 sg13g2_fill_2 FILLER_3_536 ();
 sg13g2_fill_2 FILLER_3_543 ();
 sg13g2_fill_1 FILLER_3_558 ();
 sg13g2_fill_1 FILLER_3_630 ();
 sg13g2_fill_1 FILLER_3_664 ();
 sg13g2_fill_2 FILLER_3_685 ();
 sg13g2_fill_1 FILLER_3_687 ();
 sg13g2_fill_2 FILLER_3_693 ();
 sg13g2_fill_2 FILLER_3_700 ();
 sg13g2_fill_1 FILLER_3_702 ();
 sg13g2_decap_4 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_716 ();
 sg13g2_fill_2 FILLER_3_723 ();
 sg13g2_fill_1 FILLER_3_725 ();
 sg13g2_fill_2 FILLER_3_731 ();
 sg13g2_fill_2 FILLER_3_741 ();
 sg13g2_fill_1 FILLER_3_751 ();
 sg13g2_fill_2 FILLER_3_760 ();
 sg13g2_fill_1 FILLER_3_855 ();
 sg13g2_fill_2 FILLER_3_932 ();
 sg13g2_fill_2 FILLER_3_971 ();
 sg13g2_fill_1 FILLER_3_973 ();
 sg13g2_fill_1 FILLER_3_1010 ();
 sg13g2_fill_2 FILLER_3_1038 ();
 sg13g2_fill_1 FILLER_3_1040 ();
 sg13g2_fill_2 FILLER_3_1068 ();
 sg13g2_fill_1 FILLER_3_1208 ();
 sg13g2_fill_2 FILLER_3_1284 ();
 sg13g2_fill_1 FILLER_3_1286 ();
 sg13g2_fill_2 FILLER_3_1304 ();
 sg13g2_fill_1 FILLER_3_1306 ();
 sg13g2_fill_1 FILLER_3_1347 ();
 sg13g2_fill_2 FILLER_3_1438 ();
 sg13g2_fill_2 FILLER_3_1449 ();
 sg13g2_fill_1 FILLER_3_1451 ();
 sg13g2_fill_2 FILLER_3_1465 ();
 sg13g2_fill_1 FILLER_3_1467 ();
 sg13g2_fill_2 FILLER_3_1490 ();
 sg13g2_fill_1 FILLER_3_1492 ();
 sg13g2_fill_1 FILLER_3_1534 ();
 sg13g2_fill_2 FILLER_3_1571 ();
 sg13g2_fill_1 FILLER_3_1573 ();
 sg13g2_decap_8 FILLER_3_1741 ();
 sg13g2_decap_8 FILLER_3_1748 ();
 sg13g2_decap_8 FILLER_3_1755 ();
 sg13g2_decap_4 FILLER_3_1762 ();
 sg13g2_fill_2 FILLER_3_1766 ();
 sg13g2_fill_2 FILLER_4_34 ();
 sg13g2_fill_1 FILLER_4_43 ();
 sg13g2_decap_4 FILLER_4_61 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_fill_2 FILLER_4_78 ();
 sg13g2_fill_2 FILLER_4_85 ();
 sg13g2_decap_8 FILLER_4_99 ();
 sg13g2_fill_1 FILLER_4_106 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_170 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_decap_4 FILLER_4_184 ();
 sg13g2_fill_2 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_202 ();
 sg13g2_fill_1 FILLER_4_220 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_4 FILLER_4_252 ();
 sg13g2_fill_1 FILLER_4_256 ();
 sg13g2_decap_4 FILLER_4_261 ();
 sg13g2_fill_1 FILLER_4_265 ();
 sg13g2_fill_1 FILLER_4_315 ();
 sg13g2_fill_2 FILLER_4_410 ();
 sg13g2_fill_1 FILLER_4_412 ();
 sg13g2_fill_2 FILLER_4_439 ();
 sg13g2_fill_2 FILLER_4_456 ();
 sg13g2_fill_2 FILLER_4_490 ();
 sg13g2_fill_1 FILLER_4_492 ();
 sg13g2_fill_2 FILLER_4_508 ();
 sg13g2_fill_1 FILLER_4_528 ();
 sg13g2_decap_4 FILLER_4_553 ();
 sg13g2_fill_1 FILLER_4_557 ();
 sg13g2_fill_2 FILLER_4_568 ();
 sg13g2_fill_1 FILLER_4_575 ();
 sg13g2_decap_4 FILLER_4_598 ();
 sg13g2_fill_1 FILLER_4_602 ();
 sg13g2_fill_2 FILLER_4_607 ();
 sg13g2_fill_2 FILLER_4_629 ();
 sg13g2_decap_4 FILLER_4_651 ();
 sg13g2_fill_1 FILLER_4_659 ();
 sg13g2_fill_2 FILLER_4_664 ();
 sg13g2_fill_1 FILLER_4_666 ();
 sg13g2_fill_1 FILLER_4_703 ();
 sg13g2_fill_2 FILLER_4_716 ();
 sg13g2_fill_1 FILLER_4_751 ();
 sg13g2_fill_2 FILLER_4_770 ();
 sg13g2_fill_1 FILLER_4_772 ();
 sg13g2_fill_2 FILLER_4_833 ();
 sg13g2_decap_4 FILLER_4_874 ();
 sg13g2_fill_2 FILLER_4_887 ();
 sg13g2_fill_1 FILLER_4_889 ();
 sg13g2_fill_2 FILLER_4_925 ();
 sg13g2_fill_2 FILLER_4_944 ();
 sg13g2_fill_1 FILLER_4_946 ();
 sg13g2_fill_1 FILLER_4_983 ();
 sg13g2_fill_1 FILLER_4_1002 ();
 sg13g2_fill_2 FILLER_4_1101 ();
 sg13g2_fill_1 FILLER_4_1103 ();
 sg13g2_fill_1 FILLER_4_1140 ();
 sg13g2_fill_2 FILLER_4_1168 ();
 sg13g2_fill_1 FILLER_4_1280 ();
 sg13g2_fill_2 FILLER_4_1318 ();
 sg13g2_fill_1 FILLER_4_1320 ();
 sg13g2_fill_1 FILLER_4_1330 ();
 sg13g2_fill_1 FILLER_4_1362 ();
 sg13g2_fill_1 FILLER_4_1416 ();
 sg13g2_fill_2 FILLER_4_1448 ();
 sg13g2_fill_2 FILLER_4_1554 ();
 sg13g2_fill_1 FILLER_4_1556 ();
 sg13g2_fill_2 FILLER_4_1616 ();
 sg13g2_fill_2 FILLER_4_1676 ();
 sg13g2_fill_1 FILLER_4_1678 ();
 sg13g2_fill_2 FILLER_4_1692 ();
 sg13g2_fill_1 FILLER_4_1694 ();
 sg13g2_decap_8 FILLER_4_1752 ();
 sg13g2_decap_8 FILLER_4_1759 ();
 sg13g2_fill_2 FILLER_4_1766 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_27 ();
 sg13g2_fill_1 FILLER_5_29 ();
 sg13g2_decap_8 FILLER_5_38 ();
 sg13g2_fill_1 FILLER_5_84 ();
 sg13g2_fill_2 FILLER_5_93 ();
 sg13g2_fill_1 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_113 ();
 sg13g2_decap_4 FILLER_5_120 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_fill_2 FILLER_5_144 ();
 sg13g2_fill_2 FILLER_5_171 ();
 sg13g2_decap_4 FILLER_5_190 ();
 sg13g2_decap_4 FILLER_5_219 ();
 sg13g2_fill_1 FILLER_5_228 ();
 sg13g2_decap_4 FILLER_5_241 ();
 sg13g2_fill_1 FILLER_5_245 ();
 sg13g2_fill_2 FILLER_5_272 ();
 sg13g2_fill_1 FILLER_5_274 ();
 sg13g2_fill_2 FILLER_5_371 ();
 sg13g2_fill_2 FILLER_5_378 ();
 sg13g2_fill_1 FILLER_5_380 ();
 sg13g2_fill_2 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_decap_4 FILLER_5_429 ();
 sg13g2_fill_2 FILLER_5_433 ();
 sg13g2_decap_8 FILLER_5_444 ();
 sg13g2_fill_1 FILLER_5_451 ();
 sg13g2_fill_1 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_fill_2 FILLER_5_480 ();
 sg13g2_fill_1 FILLER_5_482 ();
 sg13g2_fill_1 FILLER_5_526 ();
 sg13g2_fill_1 FILLER_5_532 ();
 sg13g2_fill_2 FILLER_5_552 ();
 sg13g2_fill_1 FILLER_5_554 ();
 sg13g2_fill_2 FILLER_5_560 ();
 sg13g2_fill_2 FILLER_5_572 ();
 sg13g2_fill_1 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_603 ();
 sg13g2_decap_4 FILLER_5_610 ();
 sg13g2_fill_1 FILLER_5_614 ();
 sg13g2_decap_4 FILLER_5_642 ();
 sg13g2_fill_2 FILLER_5_663 ();
 sg13g2_fill_1 FILLER_5_665 ();
 sg13g2_fill_1 FILLER_5_684 ();
 sg13g2_decap_4 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_720 ();
 sg13g2_decap_8 FILLER_5_727 ();
 sg13g2_decap_8 FILLER_5_734 ();
 sg13g2_fill_2 FILLER_5_748 ();
 sg13g2_fill_2 FILLER_5_775 ();
 sg13g2_fill_1 FILLER_5_777 ();
 sg13g2_fill_2 FILLER_5_822 ();
 sg13g2_fill_1 FILLER_5_824 ();
 sg13g2_decap_4 FILLER_5_869 ();
 sg13g2_fill_1 FILLER_5_1034 ();
 sg13g2_fill_2 FILLER_5_1075 ();
 sg13g2_fill_2 FILLER_5_1153 ();
 sg13g2_fill_1 FILLER_5_1155 ();
 sg13g2_fill_1 FILLER_5_1275 ();
 sg13g2_fill_2 FILLER_5_1303 ();
 sg13g2_fill_2 FILLER_5_1395 ();
 sg13g2_fill_2 FILLER_5_1437 ();
 sg13g2_fill_1 FILLER_5_1439 ();
 sg13g2_fill_1 FILLER_5_1481 ();
 sg13g2_fill_1 FILLER_5_1504 ();
 sg13g2_fill_1 FILLER_5_1542 ();
 sg13g2_fill_2 FILLER_5_1574 ();
 sg13g2_fill_1 FILLER_5_1576 ();
 sg13g2_decap_8 FILLER_5_1756 ();
 sg13g2_decap_4 FILLER_5_1763 ();
 sg13g2_fill_1 FILLER_5_1767 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_36 ();
 sg13g2_fill_1 FILLER_6_43 ();
 sg13g2_fill_1 FILLER_6_61 ();
 sg13g2_decap_8 FILLER_6_99 ();
 sg13g2_fill_2 FILLER_6_118 ();
 sg13g2_fill_1 FILLER_6_120 ();
 sg13g2_fill_1 FILLER_6_145 ();
 sg13g2_decap_4 FILLER_6_188 ();
 sg13g2_fill_1 FILLER_6_192 ();
 sg13g2_fill_2 FILLER_6_197 ();
 sg13g2_fill_1 FILLER_6_219 ();
 sg13g2_decap_4 FILLER_6_237 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_fill_2 FILLER_6_255 ();
 sg13g2_fill_2 FILLER_6_317 ();
 sg13g2_fill_2 FILLER_6_337 ();
 sg13g2_fill_1 FILLER_6_339 ();
 sg13g2_fill_2 FILLER_6_368 ();
 sg13g2_fill_1 FILLER_6_370 ();
 sg13g2_fill_1 FILLER_6_386 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_fill_1 FILLER_6_414 ();
 sg13g2_decap_4 FILLER_6_442 ();
 sg13g2_fill_1 FILLER_6_446 ();
 sg13g2_fill_2 FILLER_6_492 ();
 sg13g2_fill_1 FILLER_6_494 ();
 sg13g2_fill_2 FILLER_6_508 ();
 sg13g2_fill_2 FILLER_6_528 ();
 sg13g2_fill_1 FILLER_6_530 ();
 sg13g2_decap_4 FILLER_6_554 ();
 sg13g2_fill_1 FILLER_6_563 ();
 sg13g2_fill_1 FILLER_6_574 ();
 sg13g2_fill_2 FILLER_6_584 ();
 sg13g2_fill_1 FILLER_6_586 ();
 sg13g2_fill_1 FILLER_6_597 ();
 sg13g2_fill_1 FILLER_6_603 ();
 sg13g2_fill_1 FILLER_6_612 ();
 sg13g2_fill_2 FILLER_6_617 ();
 sg13g2_fill_1 FILLER_6_619 ();
 sg13g2_decap_8 FILLER_6_624 ();
 sg13g2_fill_2 FILLER_6_631 ();
 sg13g2_fill_1 FILLER_6_633 ();
 sg13g2_fill_2 FILLER_6_692 ();
 sg13g2_decap_4 FILLER_6_707 ();
 sg13g2_fill_1 FILLER_6_711 ();
 sg13g2_fill_2 FILLER_6_758 ();
 sg13g2_fill_1 FILLER_6_794 ();
 sg13g2_fill_2 FILLER_6_853 ();
 sg13g2_fill_2 FILLER_6_886 ();
 sg13g2_fill_2 FILLER_6_950 ();
 sg13g2_fill_2 FILLER_6_956 ();
 sg13g2_fill_1 FILLER_6_958 ();
 sg13g2_fill_2 FILLER_6_995 ();
 sg13g2_fill_1 FILLER_6_997 ();
 sg13g2_decap_4 FILLER_6_1015 ();
 sg13g2_fill_2 FILLER_6_1019 ();
 sg13g2_decap_8 FILLER_6_1025 ();
 sg13g2_fill_2 FILLER_6_1086 ();
 sg13g2_fill_1 FILLER_6_1088 ();
 sg13g2_fill_1 FILLER_6_1138 ();
 sg13g2_fill_1 FILLER_6_1188 ();
 sg13g2_fill_2 FILLER_6_1302 ();
 sg13g2_fill_2 FILLER_6_1428 ();
 sg13g2_fill_1 FILLER_6_1518 ();
 sg13g2_fill_1 FILLER_6_1529 ();
 sg13g2_fill_2 FILLER_6_1557 ();
 sg13g2_fill_1 FILLER_6_1559 ();
 sg13g2_fill_2 FILLER_6_1698 ();
 sg13g2_fill_1 FILLER_6_1700 ();
 sg13g2_decap_8 FILLER_6_1760 ();
 sg13g2_fill_1 FILLER_6_1767 ();
 sg13g2_fill_2 FILLER_7_29 ();
 sg13g2_fill_1 FILLER_7_31 ();
 sg13g2_decap_4 FILLER_7_57 ();
 sg13g2_fill_2 FILLER_7_61 ();
 sg13g2_decap_4 FILLER_7_68 ();
 sg13g2_fill_2 FILLER_7_72 ();
 sg13g2_decap_8 FILLER_7_78 ();
 sg13g2_fill_2 FILLER_7_85 ();
 sg13g2_fill_1 FILLER_7_87 ();
 sg13g2_decap_8 FILLER_7_97 ();
 sg13g2_fill_2 FILLER_7_104 ();
 sg13g2_decap_4 FILLER_7_114 ();
 sg13g2_fill_2 FILLER_7_118 ();
 sg13g2_fill_2 FILLER_7_142 ();
 sg13g2_fill_1 FILLER_7_144 ();
 sg13g2_fill_2 FILLER_7_166 ();
 sg13g2_decap_8 FILLER_7_176 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_fill_1 FILLER_7_185 ();
 sg13g2_fill_2 FILLER_7_216 ();
 sg13g2_fill_1 FILLER_7_218 ();
 sg13g2_decap_8 FILLER_7_235 ();
 sg13g2_fill_1 FILLER_7_242 ();
 sg13g2_fill_1 FILLER_7_345 ();
 sg13g2_fill_2 FILLER_7_474 ();
 sg13g2_fill_1 FILLER_7_484 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_4 FILLER_7_497 ();
 sg13g2_fill_1 FILLER_7_501 ();
 sg13g2_fill_2 FILLER_7_507 ();
 sg13g2_fill_1 FILLER_7_509 ();
 sg13g2_fill_1 FILLER_7_515 ();
 sg13g2_fill_2 FILLER_7_526 ();
 sg13g2_fill_2 FILLER_7_536 ();
 sg13g2_fill_1 FILLER_7_549 ();
 sg13g2_fill_2 FILLER_7_560 ();
 sg13g2_fill_1 FILLER_7_562 ();
 sg13g2_decap_4 FILLER_7_566 ();
 sg13g2_fill_2 FILLER_7_570 ();
 sg13g2_fill_2 FILLER_7_586 ();
 sg13g2_fill_1 FILLER_7_598 ();
 sg13g2_fill_2 FILLER_7_649 ();
 sg13g2_fill_1 FILLER_7_651 ();
 sg13g2_decap_4 FILLER_7_656 ();
 sg13g2_fill_2 FILLER_7_660 ();
 sg13g2_decap_4 FILLER_7_665 ();
 sg13g2_fill_2 FILLER_7_669 ();
 sg13g2_fill_2 FILLER_7_702 ();
 sg13g2_fill_1 FILLER_7_704 ();
 sg13g2_decap_8 FILLER_7_724 ();
 sg13g2_decap_4 FILLER_7_731 ();
 sg13g2_decap_8 FILLER_7_754 ();
 sg13g2_decap_4 FILLER_7_761 ();
 sg13g2_fill_2 FILLER_7_765 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_fill_2 FILLER_7_791 ();
 sg13g2_fill_2 FILLER_7_810 ();
 sg13g2_fill_1 FILLER_7_812 ();
 sg13g2_fill_2 FILLER_7_858 ();
 sg13g2_fill_2 FILLER_7_887 ();
 sg13g2_fill_1 FILLER_7_889 ();
 sg13g2_decap_4 FILLER_7_903 ();
 sg13g2_fill_2 FILLER_7_938 ();
 sg13g2_fill_1 FILLER_7_949 ();
 sg13g2_fill_2 FILLER_7_981 ();
 sg13g2_fill_1 FILLER_7_983 ();
 sg13g2_fill_2 FILLER_7_1028 ();
 sg13g2_fill_2 FILLER_7_1058 ();
 sg13g2_fill_1 FILLER_7_1069 ();
 sg13g2_fill_2 FILLER_7_1165 ();
 sg13g2_fill_1 FILLER_7_1167 ();
 sg13g2_fill_1 FILLER_7_1212 ();
 sg13g2_fill_2 FILLER_7_1308 ();
 sg13g2_fill_2 FILLER_7_1337 ();
 sg13g2_fill_2 FILLER_7_1366 ();
 sg13g2_fill_2 FILLER_7_1385 ();
 sg13g2_fill_1 FILLER_7_1387 ();
 sg13g2_fill_2 FILLER_7_1483 ();
 sg13g2_fill_2 FILLER_7_1516 ();
 sg13g2_fill_1 FILLER_7_1518 ();
 sg13g2_fill_2 FILLER_7_1533 ();
 sg13g2_fill_1 FILLER_7_1535 ();
 sg13g2_fill_1 FILLER_7_1549 ();
 sg13g2_fill_1 FILLER_7_1621 ();
 sg13g2_fill_2 FILLER_7_1674 ();
 sg13g2_fill_1 FILLER_7_1725 ();
 sg13g2_fill_2 FILLER_7_1766 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_26 ();
 sg13g2_fill_2 FILLER_8_39 ();
 sg13g2_fill_1 FILLER_8_79 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_fill_1 FILLER_8_130 ();
 sg13g2_decap_4 FILLER_8_135 ();
 sg13g2_fill_1 FILLER_8_139 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_fill_2 FILLER_8_151 ();
 sg13g2_fill_1 FILLER_8_153 ();
 sg13g2_fill_1 FILLER_8_167 ();
 sg13g2_decap_8 FILLER_8_185 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_8_209 ();
 sg13g2_fill_2 FILLER_8_216 ();
 sg13g2_fill_1 FILLER_8_218 ();
 sg13g2_decap_8 FILLER_8_233 ();
 sg13g2_fill_1 FILLER_8_240 ();
 sg13g2_fill_2 FILLER_8_324 ();
 sg13g2_fill_1 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_358 ();
 sg13g2_fill_2 FILLER_8_373 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_fill_2 FILLER_8_389 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_fill_1 FILLER_8_427 ();
 sg13g2_fill_2 FILLER_8_452 ();
 sg13g2_fill_1 FILLER_8_454 ();
 sg13g2_decap_4 FILLER_8_489 ();
 sg13g2_fill_1 FILLER_8_493 ();
 sg13g2_fill_2 FILLER_8_516 ();
 sg13g2_fill_1 FILLER_8_518 ();
 sg13g2_fill_1 FILLER_8_534 ();
 sg13g2_fill_1 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_fill_2 FILLER_8_581 ();
 sg13g2_fill_2 FILLER_8_587 ();
 sg13g2_decap_4 FILLER_8_627 ();
 sg13g2_fill_2 FILLER_8_645 ();
 sg13g2_decap_4 FILLER_8_652 ();
 sg13g2_fill_2 FILLER_8_656 ();
 sg13g2_fill_2 FILLER_8_699 ();
 sg13g2_fill_1 FILLER_8_701 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_4 FILLER_8_725 ();
 sg13g2_fill_1 FILLER_8_729 ();
 sg13g2_decap_8 FILLER_8_758 ();
 sg13g2_decap_4 FILLER_8_765 ();
 sg13g2_fill_2 FILLER_8_796 ();
 sg13g2_fill_1 FILLER_8_798 ();
 sg13g2_fill_2 FILLER_8_839 ();
 sg13g2_fill_2 FILLER_8_872 ();
 sg13g2_fill_1 FILLER_8_874 ();
 sg13g2_decap_8 FILLER_8_902 ();
 sg13g2_fill_2 FILLER_8_967 ();
 sg13g2_fill_1 FILLER_8_969 ();
 sg13g2_fill_1 FILLER_8_1005 ();
 sg13g2_fill_1 FILLER_8_1133 ();
 sg13g2_fill_2 FILLER_8_1147 ();
 sg13g2_fill_1 FILLER_8_1171 ();
 sg13g2_fill_2 FILLER_8_1234 ();
 sg13g2_fill_1 FILLER_8_1268 ();
 sg13g2_fill_2 FILLER_8_1295 ();
 sg13g2_fill_2 FILLER_8_1360 ();
 sg13g2_fill_2 FILLER_8_1398 ();
 sg13g2_fill_2 FILLER_8_1501 ();
 sg13g2_fill_1 FILLER_8_1503 ();
 sg13g2_fill_2 FILLER_8_1572 ();
 sg13g2_fill_2 FILLER_8_1601 ();
 sg13g2_fill_1 FILLER_8_1603 ();
 sg13g2_fill_2 FILLER_8_1721 ();
 sg13g2_fill_2 FILLER_8_1757 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_11 ();
 sg13g2_decap_4 FILLER_9_22 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_decap_8 FILLER_9_36 ();
 sg13g2_fill_1 FILLER_9_43 ();
 sg13g2_decap_8 FILLER_9_55 ();
 sg13g2_decap_4 FILLER_9_62 ();
 sg13g2_fill_1 FILLER_9_66 ();
 sg13g2_decap_8 FILLER_9_71 ();
 sg13g2_decap_8 FILLER_9_78 ();
 sg13g2_fill_1 FILLER_9_85 ();
 sg13g2_decap_8 FILLER_9_94 ();
 sg13g2_fill_2 FILLER_9_101 ();
 sg13g2_fill_1 FILLER_9_103 ();
 sg13g2_decap_4 FILLER_9_112 ();
 sg13g2_fill_1 FILLER_9_116 ();
 sg13g2_fill_1 FILLER_9_149 ();
 sg13g2_fill_2 FILLER_9_155 ();
 sg13g2_fill_1 FILLER_9_157 ();
 sg13g2_decap_4 FILLER_9_162 ();
 sg13g2_fill_2 FILLER_9_166 ();
 sg13g2_fill_1 FILLER_9_173 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_fill_2 FILLER_9_185 ();
 sg13g2_fill_1 FILLER_9_187 ();
 sg13g2_fill_2 FILLER_9_216 ();
 sg13g2_fill_1 FILLER_9_218 ();
 sg13g2_fill_1 FILLER_9_223 ();
 sg13g2_fill_1 FILLER_9_252 ();
 sg13g2_fill_2 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_327 ();
 sg13g2_fill_1 FILLER_9_391 ();
 sg13g2_fill_2 FILLER_9_412 ();
 sg13g2_fill_2 FILLER_9_450 ();
 sg13g2_fill_1 FILLER_9_473 ();
 sg13g2_decap_4 FILLER_9_484 ();
 sg13g2_fill_1 FILLER_9_488 ();
 sg13g2_fill_2 FILLER_9_515 ();
 sg13g2_fill_2 FILLER_9_529 ();
 sg13g2_fill_1 FILLER_9_531 ();
 sg13g2_decap_4 FILLER_9_573 ();
 sg13g2_fill_1 FILLER_9_577 ();
 sg13g2_decap_4 FILLER_9_591 ();
 sg13g2_fill_2 FILLER_9_617 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_fill_1 FILLER_9_637 ();
 sg13g2_fill_2 FILLER_9_646 ();
 sg13g2_fill_1 FILLER_9_648 ();
 sg13g2_decap_8 FILLER_9_682 ();
 sg13g2_decap_4 FILLER_9_689 ();
 sg13g2_fill_1 FILLER_9_693 ();
 sg13g2_fill_1 FILLER_9_698 ();
 sg13g2_decap_4 FILLER_9_721 ();
 sg13g2_fill_2 FILLER_9_725 ();
 sg13g2_fill_1 FILLER_9_734 ();
 sg13g2_fill_2 FILLER_9_739 ();
 sg13g2_decap_4 FILLER_9_769 ();
 sg13g2_decap_8 FILLER_9_781 ();
 sg13g2_fill_2 FILLER_9_788 ();
 sg13g2_fill_1 FILLER_9_790 ();
 sg13g2_fill_2 FILLER_9_795 ();
 sg13g2_fill_1 FILLER_9_797 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_4 FILLER_9_819 ();
 sg13g2_fill_1 FILLER_9_823 ();
 sg13g2_fill_2 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_856 ();
 sg13g2_fill_2 FILLER_9_875 ();
 sg13g2_fill_1 FILLER_9_917 ();
 sg13g2_fill_2 FILLER_9_922 ();
 sg13g2_fill_1 FILLER_9_924 ();
 sg13g2_fill_2 FILLER_9_934 ();
 sg13g2_fill_1 FILLER_9_936 ();
 sg13g2_fill_1 FILLER_9_946 ();
 sg13g2_fill_2 FILLER_9_968 ();
 sg13g2_fill_1 FILLER_9_970 ();
 sg13g2_fill_2 FILLER_9_1007 ();
 sg13g2_decap_8 FILLER_9_1049 ();
 sg13g2_decap_4 FILLER_9_1056 ();
 sg13g2_fill_2 FILLER_9_1060 ();
 sg13g2_fill_1 FILLER_9_1074 ();
 sg13g2_decap_4 FILLER_9_1085 ();
 sg13g2_fill_2 FILLER_9_1115 ();
 sg13g2_fill_2 FILLER_9_1161 ();
 sg13g2_fill_2 FILLER_9_1180 ();
 sg13g2_fill_1 FILLER_9_1252 ();
 sg13g2_fill_2 FILLER_9_1326 ();
 sg13g2_fill_1 FILLER_9_1328 ();
 sg13g2_fill_2 FILLER_9_1369 ();
 sg13g2_fill_1 FILLER_9_1371 ();
 sg13g2_fill_2 FILLER_9_1421 ();
 sg13g2_fill_1 FILLER_9_1423 ();
 sg13g2_fill_2 FILLER_9_1490 ();
 sg13g2_fill_1 FILLER_9_1520 ();
 sg13g2_fill_2 FILLER_9_1609 ();
 sg13g2_fill_2 FILLER_9_1638 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_9 ();
 sg13g2_fill_2 FILLER_10_16 ();
 sg13g2_fill_1 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_36 ();
 sg13g2_decap_8 FILLER_10_66 ();
 sg13g2_decap_4 FILLER_10_73 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_fill_1 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_107 ();
 sg13g2_fill_1 FILLER_10_111 ();
 sg13g2_decap_4 FILLER_10_116 ();
 sg13g2_fill_2 FILLER_10_120 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_decap_4 FILLER_10_131 ();
 sg13g2_fill_2 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_4 FILLER_10_207 ();
 sg13g2_fill_2 FILLER_10_239 ();
 sg13g2_fill_1 FILLER_10_241 ();
 sg13g2_fill_1 FILLER_10_282 ();
 sg13g2_fill_2 FILLER_10_310 ();
 sg13g2_fill_2 FILLER_10_367 ();
 sg13g2_fill_1 FILLER_10_369 ();
 sg13g2_fill_1 FILLER_10_417 ();
 sg13g2_decap_4 FILLER_10_445 ();
 sg13g2_decap_4 FILLER_10_467 ();
 sg13g2_fill_1 FILLER_10_471 ();
 sg13g2_fill_2 FILLER_10_482 ();
 sg13g2_fill_1 FILLER_10_484 ();
 sg13g2_fill_2 FILLER_10_532 ();
 sg13g2_fill_1 FILLER_10_566 ();
 sg13g2_decap_8 FILLER_10_572 ();
 sg13g2_decap_8 FILLER_10_579 ();
 sg13g2_fill_2 FILLER_10_586 ();
 sg13g2_fill_1 FILLER_10_588 ();
 sg13g2_decap_4 FILLER_10_640 ();
 sg13g2_fill_1 FILLER_10_657 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_fill_1 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_716 ();
 sg13g2_decap_8 FILLER_10_723 ();
 sg13g2_decap_8 FILLER_10_730 ();
 sg13g2_decap_4 FILLER_10_741 ();
 sg13g2_fill_1 FILLER_10_745 ();
 sg13g2_decap_8 FILLER_10_750 ();
 sg13g2_decap_8 FILLER_10_757 ();
 sg13g2_decap_4 FILLER_10_821 ();
 sg13g2_fill_1 FILLER_10_825 ();
 sg13g2_fill_2 FILLER_10_893 ();
 sg13g2_fill_1 FILLER_10_895 ();
 sg13g2_decap_4 FILLER_10_909 ();
 sg13g2_decap_4 FILLER_10_917 ();
 sg13g2_fill_2 FILLER_10_921 ();
 sg13g2_fill_2 FILLER_10_990 ();
 sg13g2_decap_8 FILLER_10_1061 ();
 sg13g2_decap_4 FILLER_10_1068 ();
 sg13g2_fill_1 FILLER_10_1077 ();
 sg13g2_decap_8 FILLER_10_1091 ();
 sg13g2_fill_2 FILLER_10_1103 ();
 sg13g2_fill_1 FILLER_10_1113 ();
 sg13g2_fill_1 FILLER_10_1118 ();
 sg13g2_decap_4 FILLER_10_1129 ();
 sg13g2_decap_8 FILLER_10_1138 ();
 sg13g2_decap_4 FILLER_10_1145 ();
 sg13g2_fill_1 FILLER_10_1149 ();
 sg13g2_decap_4 FILLER_10_1160 ();
 sg13g2_fill_1 FILLER_10_1164 ();
 sg13g2_fill_1 FILLER_10_1229 ();
 sg13g2_fill_2 FILLER_10_1257 ();
 sg13g2_fill_1 FILLER_10_1259 ();
 sg13g2_fill_1 FILLER_10_1302 ();
 sg13g2_fill_2 FILLER_10_1343 ();
 sg13g2_fill_2 FILLER_10_1445 ();
 sg13g2_fill_2 FILLER_10_1460 ();
 sg13g2_fill_1 FILLER_10_1638 ();
 sg13g2_fill_1 FILLER_10_1730 ();
 sg13g2_fill_2 FILLER_11_36 ();
 sg13g2_fill_1 FILLER_11_77 ();
 sg13g2_fill_2 FILLER_11_112 ();
 sg13g2_fill_1 FILLER_11_114 ();
 sg13g2_decap_8 FILLER_11_134 ();
 sg13g2_decap_4 FILLER_11_163 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_fill_1 FILLER_11_197 ();
 sg13g2_fill_2 FILLER_11_237 ();
 sg13g2_fill_1 FILLER_11_239 ();
 sg13g2_fill_1 FILLER_11_276 ();
 sg13g2_fill_1 FILLER_11_325 ();
 sg13g2_decap_4 FILLER_11_358 ();
 sg13g2_decap_4 FILLER_11_465 ();
 sg13g2_fill_2 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_4 FILLER_11_497 ();
 sg13g2_fill_2 FILLER_11_514 ();
 sg13g2_fill_2 FILLER_11_544 ();
 sg13g2_fill_1 FILLER_11_555 ();
 sg13g2_fill_1 FILLER_11_597 ();
 sg13g2_decap_4 FILLER_11_624 ();
 sg13g2_decap_4 FILLER_11_633 ();
 sg13g2_fill_1 FILLER_11_637 ();
 sg13g2_fill_1 FILLER_11_645 ();
 sg13g2_fill_2 FILLER_11_655 ();
 sg13g2_fill_1 FILLER_11_657 ();
 sg13g2_decap_8 FILLER_11_673 ();
 sg13g2_fill_2 FILLER_11_680 ();
 sg13g2_fill_1 FILLER_11_682 ();
 sg13g2_fill_2 FILLER_11_726 ();
 sg13g2_fill_1 FILLER_11_728 ();
 sg13g2_fill_1 FILLER_11_804 ();
 sg13g2_fill_2 FILLER_11_855 ();
 sg13g2_fill_1 FILLER_11_857 ();
 sg13g2_fill_1 FILLER_11_866 ();
 sg13g2_decap_4 FILLER_11_876 ();
 sg13g2_fill_1 FILLER_11_907 ();
 sg13g2_fill_2 FILLER_11_944 ();
 sg13g2_fill_2 FILLER_11_1033 ();
 sg13g2_fill_1 FILLER_11_1044 ();
 sg13g2_fill_2 FILLER_11_1064 ();
 sg13g2_fill_1 FILLER_11_1066 ();
 sg13g2_fill_1 FILLER_11_1091 ();
 sg13g2_fill_1 FILLER_11_1097 ();
 sg13g2_fill_1 FILLER_11_1115 ();
 sg13g2_fill_2 FILLER_11_1123 ();
 sg13g2_fill_1 FILLER_11_1151 ();
 sg13g2_decap_4 FILLER_11_1168 ();
 sg13g2_fill_2 FILLER_11_1172 ();
 sg13g2_fill_1 FILLER_11_1319 ();
 sg13g2_fill_1 FILLER_11_1365 ();
 sg13g2_fill_2 FILLER_11_1388 ();
 sg13g2_fill_1 FILLER_11_1390 ();
 sg13g2_fill_2 FILLER_11_1491 ();
 sg13g2_fill_1 FILLER_11_1493 ();
 sg13g2_fill_2 FILLER_11_1507 ();
 sg13g2_fill_2 FILLER_11_1532 ();
 sg13g2_fill_1 FILLER_11_1551 ();
 sg13g2_fill_2 FILLER_11_1579 ();
 sg13g2_fill_1 FILLER_11_1581 ();
 sg13g2_fill_2 FILLER_11_1609 ();
 sg13g2_fill_1 FILLER_11_1638 ();
 sg13g2_fill_2 FILLER_11_1755 ();
 sg13g2_fill_2 FILLER_11_1766 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_36 ();
 sg13g2_fill_1 FILLER_12_38 ();
 sg13g2_fill_2 FILLER_12_55 ();
 sg13g2_decap_4 FILLER_12_62 ();
 sg13g2_fill_2 FILLER_12_90 ();
 sg13g2_fill_1 FILLER_12_105 ();
 sg13g2_decap_4 FILLER_12_110 ();
 sg13g2_fill_2 FILLER_12_114 ();
 sg13g2_decap_4 FILLER_12_130 ();
 sg13g2_fill_2 FILLER_12_134 ();
 sg13g2_fill_1 FILLER_12_153 ();
 sg13g2_fill_1 FILLER_12_167 ();
 sg13g2_fill_2 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_247 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_fill_1 FILLER_12_342 ();
 sg13g2_fill_1 FILLER_12_356 ();
 sg13g2_fill_2 FILLER_12_374 ();
 sg13g2_fill_1 FILLER_12_376 ();
 sg13g2_fill_2 FILLER_12_396 ();
 sg13g2_fill_1 FILLER_12_398 ();
 sg13g2_fill_1 FILLER_12_418 ();
 sg13g2_fill_2 FILLER_12_446 ();
 sg13g2_fill_2 FILLER_12_475 ();
 sg13g2_fill_1 FILLER_12_477 ();
 sg13g2_fill_1 FILLER_12_506 ();
 sg13g2_fill_1 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_578 ();
 sg13g2_fill_1 FILLER_12_585 ();
 sg13g2_fill_1 FILLER_12_599 ();
 sg13g2_fill_2 FILLER_12_619 ();
 sg13g2_fill_1 FILLER_12_621 ();
 sg13g2_decap_8 FILLER_12_666 ();
 sg13g2_decap_8 FILLER_12_673 ();
 sg13g2_fill_1 FILLER_12_696 ();
 sg13g2_decap_4 FILLER_12_710 ();
 sg13g2_fill_2 FILLER_12_727 ();
 sg13g2_fill_1 FILLER_12_729 ();
 sg13g2_decap_8 FILLER_12_745 ();
 sg13g2_fill_2 FILLER_12_752 ();
 sg13g2_fill_2 FILLER_12_771 ();
 sg13g2_fill_1 FILLER_12_773 ();
 sg13g2_fill_1 FILLER_12_799 ();
 sg13g2_fill_2 FILLER_12_827 ();
 sg13g2_fill_1 FILLER_12_856 ();
 sg13g2_decap_4 FILLER_12_889 ();
 sg13g2_fill_1 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_955 ();
 sg13g2_fill_1 FILLER_12_962 ();
 sg13g2_fill_1 FILLER_12_971 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_4 FILLER_12_1049 ();
 sg13g2_fill_2 FILLER_12_1071 ();
 sg13g2_decap_4 FILLER_12_1099 ();
 sg13g2_fill_1 FILLER_12_1103 ();
 sg13g2_decap_8 FILLER_12_1110 ();
 sg13g2_fill_1 FILLER_12_1117 ();
 sg13g2_fill_2 FILLER_12_1220 ();
 sg13g2_fill_2 FILLER_12_1298 ();
 sg13g2_fill_2 FILLER_12_1336 ();
 sg13g2_fill_1 FILLER_12_1338 ();
 sg13g2_fill_1 FILLER_12_1398 ();
 sg13g2_fill_1 FILLER_12_1487 ();
 sg13g2_fill_2 FILLER_12_1542 ();
 sg13g2_fill_2 FILLER_12_1556 ();
 sg13g2_fill_2 FILLER_12_1585 ();
 sg13g2_fill_1 FILLER_12_1618 ();
 sg13g2_fill_2 FILLER_12_1628 ();
 sg13g2_fill_1 FILLER_12_1665 ();
 sg13g2_fill_1 FILLER_12_1691 ();
 sg13g2_fill_2 FILLER_12_1710 ();
 sg13g2_fill_1 FILLER_12_1712 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_fill_1 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_37 ();
 sg13g2_fill_2 FILLER_13_44 ();
 sg13g2_fill_1 FILLER_13_46 ();
 sg13g2_fill_2 FILLER_13_52 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_decap_8 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_72 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_fill_1 FILLER_13_93 ();
 sg13g2_fill_1 FILLER_13_104 ();
 sg13g2_fill_1 FILLER_13_109 ();
 sg13g2_fill_2 FILLER_13_115 ();
 sg13g2_fill_1 FILLER_13_117 ();
 sg13g2_fill_2 FILLER_13_128 ();
 sg13g2_decap_8 FILLER_13_136 ();
 sg13g2_fill_1 FILLER_13_157 ();
 sg13g2_decap_4 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_229 ();
 sg13g2_fill_1 FILLER_13_231 ();
 sg13g2_fill_2 FILLER_13_267 ();
 sg13g2_fill_1 FILLER_13_269 ();
 sg13g2_fill_2 FILLER_13_288 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_2 FILLER_13_305 ();
 sg13g2_fill_1 FILLER_13_307 ();
 sg13g2_fill_1 FILLER_13_357 ();
 sg13g2_fill_1 FILLER_13_367 ();
 sg13g2_fill_1 FILLER_13_389 ();
 sg13g2_fill_1 FILLER_13_427 ();
 sg13g2_fill_2 FILLER_13_433 ();
 sg13g2_fill_1 FILLER_13_444 ();
 sg13g2_decap_4 FILLER_13_462 ();
 sg13g2_fill_2 FILLER_13_466 ();
 sg13g2_fill_2 FILLER_13_478 ();
 sg13g2_decap_4 FILLER_13_498 ();
 sg13g2_fill_1 FILLER_13_553 ();
 sg13g2_fill_1 FILLER_13_604 ();
 sg13g2_decap_4 FILLER_13_623 ();
 sg13g2_fill_2 FILLER_13_632 ();
 sg13g2_fill_2 FILLER_13_656 ();
 sg13g2_fill_1 FILLER_13_658 ();
 sg13g2_fill_2 FILLER_13_676 ();
 sg13g2_fill_1 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_708 ();
 sg13g2_decap_4 FILLER_13_715 ();
 sg13g2_fill_1 FILLER_13_735 ();
 sg13g2_decap_4 FILLER_13_741 ();
 sg13g2_fill_1 FILLER_13_745 ();
 sg13g2_decap_4 FILLER_13_767 ();
 sg13g2_fill_1 FILLER_13_803 ();
 sg13g2_fill_1 FILLER_13_829 ();
 sg13g2_decap_8 FILLER_13_857 ();
 sg13g2_fill_1 FILLER_13_864 ();
 sg13g2_fill_1 FILLER_13_869 ();
 sg13g2_decap_4 FILLER_13_879 ();
 sg13g2_decap_4 FILLER_13_914 ();
 sg13g2_fill_2 FILLER_13_954 ();
 sg13g2_fill_1 FILLER_13_956 ();
 sg13g2_fill_2 FILLER_13_1003 ();
 sg13g2_fill_1 FILLER_13_1032 ();
 sg13g2_fill_2 FILLER_13_1039 ();
 sg13g2_fill_1 FILLER_13_1041 ();
 sg13g2_fill_2 FILLER_13_1068 ();
 sg13g2_fill_2 FILLER_13_1095 ();
 sg13g2_fill_1 FILLER_13_1097 ();
 sg13g2_decap_8 FILLER_13_1112 ();
 sg13g2_decap_8 FILLER_13_1119 ();
 sg13g2_decap_4 FILLER_13_1141 ();
 sg13g2_fill_1 FILLER_13_1145 ();
 sg13g2_fill_2 FILLER_13_1172 ();
 sg13g2_fill_1 FILLER_13_1174 ();
 sg13g2_fill_2 FILLER_13_1252 ();
 sg13g2_fill_2 FILLER_13_1317 ();
 sg13g2_fill_2 FILLER_13_1391 ();
 sg13g2_fill_1 FILLER_13_1470 ();
 sg13g2_fill_1 FILLER_13_1590 ();
 sg13g2_fill_2 FILLER_13_1617 ();
 sg13g2_fill_1 FILLER_13_1619 ();
 sg13g2_fill_2 FILLER_13_1737 ();
 sg13g2_fill_1 FILLER_13_1739 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_1 FILLER_14_27 ();
 sg13g2_fill_1 FILLER_14_56 ();
 sg13g2_fill_1 FILLER_14_71 ();
 sg13g2_fill_2 FILLER_14_82 ();
 sg13g2_decap_8 FILLER_14_90 ();
 sg13g2_fill_2 FILLER_14_97 ();
 sg13g2_fill_1 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_118 ();
 sg13g2_fill_1 FILLER_14_125 ();
 sg13g2_decap_4 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_140 ();
 sg13g2_fill_2 FILLER_14_154 ();
 sg13g2_fill_2 FILLER_14_170 ();
 sg13g2_fill_1 FILLER_14_313 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_fill_2 FILLER_14_375 ();
 sg13g2_fill_1 FILLER_14_377 ();
 sg13g2_fill_2 FILLER_14_391 ();
 sg13g2_fill_1 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_fill_1 FILLER_14_469 ();
 sg13g2_fill_2 FILLER_14_510 ();
 sg13g2_fill_2 FILLER_14_539 ();
 sg13g2_fill_2 FILLER_14_607 ();
 sg13g2_decap_8 FILLER_14_632 ();
 sg13g2_fill_2 FILLER_14_659 ();
 sg13g2_fill_1 FILLER_14_672 ();
 sg13g2_decap_4 FILLER_14_702 ();
 sg13g2_fill_2 FILLER_14_706 ();
 sg13g2_fill_1 FILLER_14_731 ();
 sg13g2_decap_4 FILLER_14_737 ();
 sg13g2_decap_4 FILLER_14_764 ();
 sg13g2_decap_8 FILLER_14_773 ();
 sg13g2_fill_2 FILLER_14_811 ();
 sg13g2_fill_1 FILLER_14_813 ();
 sg13g2_fill_1 FILLER_14_847 ();
 sg13g2_fill_2 FILLER_14_858 ();
 sg13g2_decap_4 FILLER_14_892 ();
 sg13g2_fill_1 FILLER_14_896 ();
 sg13g2_fill_2 FILLER_14_938 ();
 sg13g2_fill_1 FILLER_14_940 ();
 sg13g2_fill_2 FILLER_14_963 ();
 sg13g2_fill_1 FILLER_14_975 ();
 sg13g2_fill_1 FILLER_14_985 ();
 sg13g2_decap_4 FILLER_14_990 ();
 sg13g2_fill_1 FILLER_14_994 ();
 sg13g2_fill_1 FILLER_14_999 ();
 sg13g2_fill_2 FILLER_14_1028 ();
 sg13g2_fill_2 FILLER_14_1065 ();
 sg13g2_fill_1 FILLER_14_1072 ();
 sg13g2_decap_8 FILLER_14_1089 ();
 sg13g2_fill_1 FILLER_14_1096 ();
 sg13g2_fill_2 FILLER_14_1109 ();
 sg13g2_fill_1 FILLER_14_1111 ();
 sg13g2_fill_2 FILLER_14_1134 ();
 sg13g2_fill_2 FILLER_14_1142 ();
 sg13g2_fill_1 FILLER_14_1144 ();
 sg13g2_fill_2 FILLER_14_1157 ();
 sg13g2_fill_1 FILLER_14_1159 ();
 sg13g2_decap_4 FILLER_14_1166 ();
 sg13g2_fill_1 FILLER_14_1170 ();
 sg13g2_decap_4 FILLER_14_1181 ();
 sg13g2_decap_8 FILLER_14_1189 ();
 sg13g2_fill_2 FILLER_14_1196 ();
 sg13g2_fill_1 FILLER_14_1250 ();
 sg13g2_fill_2 FILLER_14_1332 ();
 sg13g2_fill_2 FILLER_14_1347 ();
 sg13g2_fill_1 FILLER_14_1349 ();
 sg13g2_fill_1 FILLER_14_1399 ();
 sg13g2_fill_1 FILLER_14_1422 ();
 sg13g2_fill_1 FILLER_14_1520 ();
 sg13g2_fill_2 FILLER_14_1544 ();
 sg13g2_fill_2 FILLER_14_1574 ();
 sg13g2_fill_1 FILLER_14_1603 ();
 sg13g2_fill_2 FILLER_14_1676 ();
 sg13g2_fill_1 FILLER_14_1678 ();
 sg13g2_fill_1 FILLER_14_1697 ();
 sg13g2_fill_2 FILLER_14_1738 ();
 sg13g2_fill_2 FILLER_14_1765 ();
 sg13g2_fill_1 FILLER_14_1767 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_61 ();
 sg13g2_decap_4 FILLER_15_68 ();
 sg13g2_fill_1 FILLER_15_72 ();
 sg13g2_decap_4 FILLER_15_95 ();
 sg13g2_fill_1 FILLER_15_99 ();
 sg13g2_fill_2 FILLER_15_114 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_2 FILLER_15_229 ();
 sg13g2_fill_1 FILLER_15_250 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_266 ();
 sg13g2_fill_1 FILLER_15_341 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_fill_1 FILLER_15_372 ();
 sg13g2_fill_1 FILLER_15_378 ();
 sg13g2_fill_2 FILLER_15_389 ();
 sg13g2_decap_4 FILLER_15_422 ();
 sg13g2_fill_1 FILLER_15_445 ();
 sg13g2_decap_4 FILLER_15_459 ();
 sg13g2_fill_1 FILLER_15_463 ();
 sg13g2_fill_2 FILLER_15_564 ();
 sg13g2_fill_1 FILLER_15_566 ();
 sg13g2_fill_1 FILLER_15_580 ();
 sg13g2_fill_1 FILLER_15_619 ();
 sg13g2_fill_2 FILLER_15_625 ();
 sg13g2_fill_1 FILLER_15_627 ();
 sg13g2_fill_2 FILLER_15_640 ();
 sg13g2_fill_2 FILLER_15_666 ();
 sg13g2_fill_1 FILLER_15_668 ();
 sg13g2_fill_2 FILLER_15_674 ();
 sg13g2_decap_4 FILLER_15_694 ();
 sg13g2_fill_1 FILLER_15_698 ();
 sg13g2_decap_4 FILLER_15_708 ();
 sg13g2_fill_2 FILLER_15_712 ();
 sg13g2_fill_2 FILLER_15_730 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_fill_1 FILLER_15_749 ();
 sg13g2_fill_2 FILLER_15_755 ();
 sg13g2_fill_2 FILLER_15_770 ();
 sg13g2_fill_1 FILLER_15_772 ();
 sg13g2_fill_1 FILLER_15_790 ();
 sg13g2_fill_1 FILLER_15_815 ();
 sg13g2_fill_1 FILLER_15_821 ();
 sg13g2_fill_2 FILLER_15_893 ();
 sg13g2_fill_2 FILLER_15_927 ();
 sg13g2_fill_2 FILLER_15_957 ();
 sg13g2_fill_1 FILLER_15_959 ();
 sg13g2_fill_1 FILLER_15_990 ();
 sg13g2_fill_2 FILLER_15_995 ();
 sg13g2_fill_1 FILLER_15_997 ();
 sg13g2_fill_2 FILLER_15_1021 ();
 sg13g2_fill_1 FILLER_15_1023 ();
 sg13g2_decap_4 FILLER_15_1046 ();
 sg13g2_fill_2 FILLER_15_1050 ();
 sg13g2_decap_8 FILLER_15_1064 ();
 sg13g2_fill_1 FILLER_15_1071 ();
 sg13g2_decap_4 FILLER_15_1119 ();
 sg13g2_fill_2 FILLER_15_1145 ();
 sg13g2_fill_1 FILLER_15_1147 ();
 sg13g2_decap_4 FILLER_15_1160 ();
 sg13g2_fill_1 FILLER_15_1164 ();
 sg13g2_fill_1 FILLER_15_1205 ();
 sg13g2_fill_2 FILLER_15_1304 ();
 sg13g2_fill_2 FILLER_15_1333 ();
 sg13g2_fill_1 FILLER_15_1384 ();
 sg13g2_fill_2 FILLER_15_1417 ();
 sg13g2_fill_1 FILLER_15_1419 ();
 sg13g2_fill_1 FILLER_15_1598 ();
 sg13g2_fill_2 FILLER_15_1649 ();
 sg13g2_fill_1 FILLER_15_1651 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_31 ();
 sg13g2_fill_2 FILLER_16_65 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_decap_4 FILLER_16_81 ();
 sg13g2_fill_2 FILLER_16_85 ();
 sg13g2_fill_1 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_120 ();
 sg13g2_decap_8 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_143 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_197 ();
 sg13g2_fill_2 FILLER_16_235 ();
 sg13g2_fill_2 FILLER_16_270 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_fill_2 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_325 ();
 sg13g2_fill_2 FILLER_16_385 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_fill_2 FILLER_16_462 ();
 sg13g2_fill_1 FILLER_16_464 ();
 sg13g2_fill_1 FILLER_16_475 ();
 sg13g2_fill_1 FILLER_16_512 ();
 sg13g2_fill_2 FILLER_16_523 ();
 sg13g2_fill_1 FILLER_16_525 ();
 sg13g2_fill_2 FILLER_16_545 ();
 sg13g2_fill_2 FILLER_16_556 ();
 sg13g2_fill_1 FILLER_16_558 ();
 sg13g2_decap_4 FILLER_16_610 ();
 sg13g2_fill_2 FILLER_16_619 ();
 sg13g2_fill_1 FILLER_16_631 ();
 sg13g2_fill_1 FILLER_16_637 ();
 sg13g2_fill_1 FILLER_16_671 ();
 sg13g2_fill_1 FILLER_16_681 ();
 sg13g2_fill_2 FILLER_16_692 ();
 sg13g2_fill_2 FILLER_16_709 ();
 sg13g2_fill_1 FILLER_16_711 ();
 sg13g2_decap_8 FILLER_16_716 ();
 sg13g2_decap_8 FILLER_16_723 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_fill_2 FILLER_16_742 ();
 sg13g2_fill_1 FILLER_16_757 ();
 sg13g2_fill_2 FILLER_16_813 ();
 sg13g2_fill_1 FILLER_16_831 ();
 sg13g2_fill_2 FILLER_16_840 ();
 sg13g2_fill_1 FILLER_16_875 ();
 sg13g2_fill_2 FILLER_16_889 ();
 sg13g2_fill_2 FILLER_16_918 ();
 sg13g2_fill_1 FILLER_16_920 ();
 sg13g2_fill_1 FILLER_16_938 ();
 sg13g2_fill_2 FILLER_16_974 ();
 sg13g2_fill_2 FILLER_16_1024 ();
 sg13g2_decap_8 FILLER_16_1043 ();
 sg13g2_decap_4 FILLER_16_1050 ();
 sg13g2_decap_8 FILLER_16_1070 ();
 sg13g2_decap_4 FILLER_16_1077 ();
 sg13g2_fill_1 FILLER_16_1092 ();
 sg13g2_fill_2 FILLER_16_1141 ();
 sg13g2_fill_2 FILLER_16_1163 ();
 sg13g2_fill_1 FILLER_16_1165 ();
 sg13g2_fill_1 FILLER_16_1174 ();
 sg13g2_fill_2 FILLER_16_1184 ();
 sg13g2_fill_1 FILLER_16_1186 ();
 sg13g2_fill_1 FILLER_16_1232 ();
 sg13g2_fill_1 FILLER_16_1251 ();
 sg13g2_fill_1 FILLER_16_1321 ();
 sg13g2_fill_1 FILLER_16_1400 ();
 sg13g2_fill_2 FILLER_16_1477 ();
 sg13g2_fill_2 FILLER_16_1513 ();
 sg13g2_fill_1 FILLER_16_1565 ();
 sg13g2_fill_1 FILLER_16_1570 ();
 sg13g2_fill_2 FILLER_16_1592 ();
 sg13g2_fill_2 FILLER_16_1634 ();
 sg13g2_fill_1 FILLER_16_1707 ();
 sg13g2_fill_1 FILLER_16_1756 ();
 sg13g2_fill_2 FILLER_16_1766 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_14 ();
 sg13g2_decap_4 FILLER_17_40 ();
 sg13g2_decap_4 FILLER_17_68 ();
 sg13g2_fill_1 FILLER_17_100 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_fill_2 FILLER_17_112 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_137 ();
 sg13g2_fill_1 FILLER_17_153 ();
 sg13g2_decap_4 FILLER_17_169 ();
 sg13g2_decap_8 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_206 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_242 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_369 ();
 sg13g2_fill_2 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_388 ();
 sg13g2_fill_2 FILLER_17_395 ();
 sg13g2_fill_1 FILLER_17_397 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_521 ();
 sg13g2_fill_1 FILLER_17_546 ();
 sg13g2_fill_1 FILLER_17_575 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_fill_2 FILLER_17_630 ();
 sg13g2_decap_4 FILLER_17_642 ();
 sg13g2_decap_8 FILLER_17_654 ();
 sg13g2_fill_2 FILLER_17_661 ();
 sg13g2_decap_4 FILLER_17_686 ();
 sg13g2_fill_1 FILLER_17_690 ();
 sg13g2_fill_1 FILLER_17_697 ();
 sg13g2_fill_1 FILLER_17_735 ();
 sg13g2_fill_2 FILLER_17_757 ();
 sg13g2_fill_1 FILLER_17_773 ();
 sg13g2_fill_1 FILLER_17_833 ();
 sg13g2_fill_1 FILLER_17_856 ();
 sg13g2_fill_1 FILLER_17_866 ();
 sg13g2_fill_2 FILLER_17_875 ();
 sg13g2_fill_2 FILLER_17_918 ();
 sg13g2_fill_1 FILLER_17_920 ();
 sg13g2_decap_4 FILLER_17_966 ();
 sg13g2_fill_2 FILLER_17_979 ();
 sg13g2_fill_1 FILLER_17_981 ();
 sg13g2_decap_8 FILLER_17_1011 ();
 sg13g2_decap_4 FILLER_17_1018 ();
 sg13g2_fill_1 FILLER_17_1022 ();
 sg13g2_fill_2 FILLER_17_1064 ();
 sg13g2_fill_1 FILLER_17_1066 ();
 sg13g2_decap_4 FILLER_17_1087 ();
 sg13g2_fill_1 FILLER_17_1100 ();
 sg13g2_decap_8 FILLER_17_1113 ();
 sg13g2_decap_4 FILLER_17_1120 ();
 sg13g2_decap_8 FILLER_17_1136 ();
 sg13g2_fill_1 FILLER_17_1143 ();
 sg13g2_decap_8 FILLER_17_1158 ();
 sg13g2_fill_1 FILLER_17_1196 ();
 sg13g2_fill_1 FILLER_17_1278 ();
 sg13g2_fill_2 FILLER_17_1309 ();
 sg13g2_fill_1 FILLER_17_1311 ();
 sg13g2_fill_2 FILLER_17_1375 ();
 sg13g2_fill_1 FILLER_17_1377 ();
 sg13g2_fill_1 FILLER_17_1427 ();
 sg13g2_fill_1 FILLER_17_1445 ();
 sg13g2_fill_1 FILLER_17_1511 ();
 sg13g2_fill_2 FILLER_17_1543 ();
 sg13g2_fill_2 FILLER_17_1572 ();
 sg13g2_fill_1 FILLER_17_1601 ();
 sg13g2_fill_2 FILLER_17_1673 ();
 sg13g2_fill_1 FILLER_17_1739 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_43 ();
 sg13g2_fill_2 FILLER_18_58 ();
 sg13g2_fill_1 FILLER_18_60 ();
 sg13g2_decap_4 FILLER_18_72 ();
 sg13g2_decap_8 FILLER_18_86 ();
 sg13g2_fill_2 FILLER_18_93 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_120 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_1 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_fill_2 FILLER_18_168 ();
 sg13g2_decap_4 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_fill_2 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_fill_2 FILLER_18_241 ();
 sg13g2_fill_1 FILLER_18_243 ();
 sg13g2_fill_2 FILLER_18_342 ();
 sg13g2_fill_2 FILLER_18_404 ();
 sg13g2_fill_2 FILLER_18_431 ();
 sg13g2_decap_4 FILLER_18_437 ();
 sg13g2_fill_1 FILLER_18_441 ();
 sg13g2_fill_2 FILLER_18_446 ();
 sg13g2_decap_8 FILLER_18_461 ();
 sg13g2_fill_2 FILLER_18_468 ();
 sg13g2_fill_1 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_493 ();
 sg13g2_decap_4 FILLER_18_500 ();
 sg13g2_fill_1 FILLER_18_512 ();
 sg13g2_fill_1 FILLER_18_526 ();
 sg13g2_fill_2 FILLER_18_581 ();
 sg13g2_fill_1 FILLER_18_583 ();
 sg13g2_fill_2 FILLER_18_593 ();
 sg13g2_decap_4 FILLER_18_606 ();
 sg13g2_decap_4 FILLER_18_626 ();
 sg13g2_fill_2 FILLER_18_642 ();
 sg13g2_fill_1 FILLER_18_644 ();
 sg13g2_fill_1 FILLER_18_684 ();
 sg13g2_decap_4 FILLER_18_714 ();
 sg13g2_fill_1 FILLER_18_718 ();
 sg13g2_fill_2 FILLER_18_739 ();
 sg13g2_fill_1 FILLER_18_820 ();
 sg13g2_fill_1 FILLER_18_830 ();
 sg13g2_fill_2 FILLER_18_859 ();
 sg13g2_fill_1 FILLER_18_902 ();
 sg13g2_fill_1 FILLER_18_948 ();
 sg13g2_fill_2 FILLER_18_966 ();
 sg13g2_fill_2 FILLER_18_989 ();
 sg13g2_fill_1 FILLER_18_991 ();
 sg13g2_fill_2 FILLER_18_1085 ();
 sg13g2_decap_4 FILLER_18_1112 ();
 sg13g2_fill_2 FILLER_18_1116 ();
 sg13g2_fill_1 FILLER_18_1122 ();
 sg13g2_fill_2 FILLER_18_1168 ();
 sg13g2_fill_1 FILLER_18_1170 ();
 sg13g2_fill_1 FILLER_18_1336 ();
 sg13g2_fill_1 FILLER_18_1467 ();
 sg13g2_fill_1 FILLER_18_1482 ();
 sg13g2_fill_1 FILLER_18_1505 ();
 sg13g2_fill_1 FILLER_18_1572 ();
 sg13g2_fill_1 FILLER_18_1736 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_10 ();
 sg13g2_fill_1 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_41 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_1 FILLER_19_69 ();
 sg13g2_fill_2 FILLER_19_75 ();
 sg13g2_decap_4 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_1 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_156 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_1 FILLER_19_176 ();
 sg13g2_fill_2 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_188 ();
 sg13g2_fill_1 FILLER_19_195 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_1 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_4 FILLER_19_332 ();
 sg13g2_fill_2 FILLER_19_336 ();
 sg13g2_fill_2 FILLER_19_346 ();
 sg13g2_fill_2 FILLER_19_419 ();
 sg13g2_decap_8 FILLER_19_506 ();
 sg13g2_fill_1 FILLER_19_513 ();
 sg13g2_fill_2 FILLER_19_560 ();
 sg13g2_fill_2 FILLER_19_576 ();
 sg13g2_fill_2 FILLER_19_623 ();
 sg13g2_fill_1 FILLER_19_625 ();
 sg13g2_fill_2 FILLER_19_630 ();
 sg13g2_fill_1 FILLER_19_632 ();
 sg13g2_fill_2 FILLER_19_640 ();
 sg13g2_fill_1 FILLER_19_676 ();
 sg13g2_fill_2 FILLER_19_697 ();
 sg13g2_fill_1 FILLER_19_699 ();
 sg13g2_fill_1 FILLER_19_705 ();
 sg13g2_fill_2 FILLER_19_724 ();
 sg13g2_fill_1 FILLER_19_726 ();
 sg13g2_fill_1 FILLER_19_744 ();
 sg13g2_fill_1 FILLER_19_787 ();
 sg13g2_fill_1 FILLER_19_814 ();
 sg13g2_fill_1 FILLER_19_829 ();
 sg13g2_fill_2 FILLER_19_852 ();
 sg13g2_fill_2 FILLER_19_871 ();
 sg13g2_fill_2 FILLER_19_907 ();
 sg13g2_fill_2 FILLER_19_914 ();
 sg13g2_fill_1 FILLER_19_916 ();
 sg13g2_fill_2 FILLER_19_953 ();
 sg13g2_fill_1 FILLER_19_955 ();
 sg13g2_fill_2 FILLER_19_965 ();
 sg13g2_fill_2 FILLER_19_981 ();
 sg13g2_fill_1 FILLER_19_1001 ();
 sg13g2_fill_2 FILLER_19_1010 ();
 sg13g2_fill_2 FILLER_19_1083 ();
 sg13g2_decap_8 FILLER_19_1104 ();
 sg13g2_fill_2 FILLER_19_1111 ();
 sg13g2_fill_1 FILLER_19_1140 ();
 sg13g2_fill_1 FILLER_19_1180 ();
 sg13g2_fill_1 FILLER_19_1190 ();
 sg13g2_fill_1 FILLER_19_1249 ();
 sg13g2_fill_2 FILLER_19_1352 ();
 sg13g2_fill_1 FILLER_19_1380 ();
 sg13g2_fill_1 FILLER_19_1390 ();
 sg13g2_fill_2 FILLER_19_1440 ();
 sg13g2_fill_1 FILLER_19_1458 ();
 sg13g2_fill_1 FILLER_19_1486 ();
 sg13g2_fill_2 FILLER_19_1514 ();
 sg13g2_fill_2 FILLER_19_1556 ();
 sg13g2_fill_2 FILLER_19_1642 ();
 sg13g2_fill_1 FILLER_19_1700 ();
 sg13g2_decap_4 FILLER_19_1763 ();
 sg13g2_fill_1 FILLER_19_1767 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_93 ();
 sg13g2_fill_1 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_fill_1 FILLER_20_150 ();
 sg13g2_fill_2 FILLER_20_158 ();
 sg13g2_fill_1 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_171 ();
 sg13g2_decap_4 FILLER_20_178 ();
 sg13g2_decap_8 FILLER_20_195 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_4 FILLER_20_271 ();
 sg13g2_decap_4 FILLER_20_367 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_fill_2 FILLER_20_399 ();
 sg13g2_fill_1 FILLER_20_401 ();
 sg13g2_fill_1 FILLER_20_413 ();
 sg13g2_fill_2 FILLER_20_454 ();
 sg13g2_fill_1 FILLER_20_495 ();
 sg13g2_fill_1 FILLER_20_551 ();
 sg13g2_fill_2 FILLER_20_597 ();
 sg13g2_fill_1 FILLER_20_599 ();
 sg13g2_fill_2 FILLER_20_618 ();
 sg13g2_fill_1 FILLER_20_620 ();
 sg13g2_fill_1 FILLER_20_634 ();
 sg13g2_fill_1 FILLER_20_643 ();
 sg13g2_fill_2 FILLER_20_677 ();
 sg13g2_decap_4 FILLER_20_705 ();
 sg13g2_fill_1 FILLER_20_709 ();
 sg13g2_fill_2 FILLER_20_755 ();
 sg13g2_fill_1 FILLER_20_757 ();
 sg13g2_fill_1 FILLER_20_782 ();
 sg13g2_fill_1 FILLER_20_805 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_fill_2 FILLER_20_914 ();
 sg13g2_fill_1 FILLER_20_916 ();
 sg13g2_decap_4 FILLER_20_975 ();
 sg13g2_fill_1 FILLER_20_996 ();
 sg13g2_fill_1 FILLER_20_1092 ();
 sg13g2_fill_2 FILLER_20_1103 ();
 sg13g2_decap_8 FILLER_20_1119 ();
 sg13g2_decap_4 FILLER_20_1126 ();
 sg13g2_fill_1 FILLER_20_1130 ();
 sg13g2_fill_2 FILLER_20_1143 ();
 sg13g2_fill_1 FILLER_20_1307 ();
 sg13g2_fill_2 FILLER_20_1347 ();
 sg13g2_fill_1 FILLER_20_1428 ();
 sg13g2_fill_2 FILLER_20_1472 ();
 sg13g2_fill_1 FILLER_20_1500 ();
 sg13g2_fill_2 FILLER_20_1515 ();
 sg13g2_fill_2 FILLER_20_1525 ();
 sg13g2_fill_2 FILLER_20_1577 ();
 sg13g2_fill_1 FILLER_20_1606 ();
 sg13g2_fill_2 FILLER_20_1636 ();
 sg13g2_decap_4 FILLER_20_1755 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_4 ();
 sg13g2_decap_4 FILLER_21_10 ();
 sg13g2_fill_1 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_57 ();
 sg13g2_fill_1 FILLER_21_66 ();
 sg13g2_fill_2 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_85 ();
 sg13g2_decap_4 FILLER_21_100 ();
 sg13g2_fill_2 FILLER_21_104 ();
 sg13g2_decap_8 FILLER_21_110 ();
 sg13g2_fill_2 FILLER_21_122 ();
 sg13g2_decap_4 FILLER_21_141 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_173 ();
 sg13g2_fill_1 FILLER_21_180 ();
 sg13g2_decap_4 FILLER_21_222 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_280 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_decap_4 FILLER_21_340 ();
 sg13g2_decap_4 FILLER_21_348 ();
 sg13g2_fill_2 FILLER_21_352 ();
 sg13g2_fill_1 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_439 ();
 sg13g2_fill_1 FILLER_21_472 ();
 sg13g2_fill_2 FILLER_21_500 ();
 sg13g2_fill_1 FILLER_21_502 ();
 sg13g2_fill_1 FILLER_21_512 ();
 sg13g2_fill_2 FILLER_21_554 ();
 sg13g2_fill_1 FILLER_21_556 ();
 sg13g2_decap_8 FILLER_21_565 ();
 sg13g2_fill_2 FILLER_21_572 ();
 sg13g2_decap_8 FILLER_21_579 ();
 sg13g2_decap_8 FILLER_21_586 ();
 sg13g2_fill_2 FILLER_21_593 ();
 sg13g2_fill_1 FILLER_21_595 ();
 sg13g2_fill_2 FILLER_21_605 ();
 sg13g2_fill_1 FILLER_21_607 ();
 sg13g2_fill_2 FILLER_21_622 ();
 sg13g2_fill_1 FILLER_21_624 ();
 sg13g2_fill_2 FILLER_21_643 ();
 sg13g2_fill_1 FILLER_21_645 ();
 sg13g2_fill_2 FILLER_21_675 ();
 sg13g2_fill_1 FILLER_21_698 ();
 sg13g2_fill_2 FILLER_21_733 ();
 sg13g2_fill_2 FILLER_21_746 ();
 sg13g2_fill_1 FILLER_21_759 ();
 sg13g2_fill_2 FILLER_21_794 ();
 sg13g2_fill_1 FILLER_21_796 ();
 sg13g2_fill_1 FILLER_21_801 ();
 sg13g2_fill_2 FILLER_21_806 ();
 sg13g2_fill_2 FILLER_21_838 ();
 sg13g2_decap_4 FILLER_21_856 ();
 sg13g2_fill_2 FILLER_21_860 ();
 sg13g2_decap_4 FILLER_21_872 ();
 sg13g2_decap_8 FILLER_21_880 ();
 sg13g2_fill_2 FILLER_21_887 ();
 sg13g2_fill_1 FILLER_21_889 ();
 sg13g2_fill_2 FILLER_21_900 ();
 sg13g2_fill_1 FILLER_21_902 ();
 sg13g2_fill_2 FILLER_21_912 ();
 sg13g2_fill_1 FILLER_21_1029 ();
 sg13g2_fill_2 FILLER_21_1178 ();
 sg13g2_fill_1 FILLER_21_1180 ();
 sg13g2_fill_1 FILLER_21_1194 ();
 sg13g2_fill_2 FILLER_21_1259 ();
 sg13g2_fill_1 FILLER_21_1261 ();
 sg13g2_fill_1 FILLER_21_1280 ();
 sg13g2_fill_1 FILLER_21_1366 ();
 sg13g2_fill_1 FILLER_21_1371 ();
 sg13g2_fill_1 FILLER_21_1428 ();
 sg13g2_fill_1 FILLER_21_1462 ();
 sg13g2_fill_1 FILLER_21_1493 ();
 sg13g2_fill_2 FILLER_21_1534 ();
 sg13g2_fill_2 FILLER_21_1579 ();
 sg13g2_fill_1 FILLER_21_1590 ();
 sg13g2_fill_2 FILLER_21_1600 ();
 sg13g2_fill_2 FILLER_21_1674 ();
 sg13g2_fill_2 FILLER_21_1684 ();
 sg13g2_fill_1 FILLER_21_1686 ();
 sg13g2_fill_2 FILLER_21_1696 ();
 sg13g2_fill_1 FILLER_21_1711 ();
 sg13g2_fill_2 FILLER_21_1757 ();
 sg13g2_fill_2 FILLER_22_31 ();
 sg13g2_fill_2 FILLER_22_42 ();
 sg13g2_fill_1 FILLER_22_44 ();
 sg13g2_fill_2 FILLER_22_65 ();
 sg13g2_fill_1 FILLER_22_94 ();
 sg13g2_fill_1 FILLER_22_111 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_145 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_fill_1 FILLER_22_186 ();
 sg13g2_decap_4 FILLER_22_208 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_224 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_fill_1 FILLER_22_268 ();
 sg13g2_fill_2 FILLER_22_277 ();
 sg13g2_fill_1 FILLER_22_305 ();
 sg13g2_decap_4 FILLER_22_326 ();
 sg13g2_fill_2 FILLER_22_330 ();
 sg13g2_fill_2 FILLER_22_432 ();
 sg13g2_fill_2 FILLER_22_461 ();
 sg13g2_fill_1 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_545 ();
 sg13g2_fill_2 FILLER_22_552 ();
 sg13g2_decap_8 FILLER_22_561 ();
 sg13g2_fill_2 FILLER_22_581 ();
 sg13g2_fill_1 FILLER_22_583 ();
 sg13g2_fill_2 FILLER_22_591 ();
 sg13g2_fill_1 FILLER_22_593 ();
 sg13g2_fill_2 FILLER_22_602 ();
 sg13g2_fill_2 FILLER_22_620 ();
 sg13g2_fill_2 FILLER_22_640 ();
 sg13g2_fill_1 FILLER_22_642 ();
 sg13g2_fill_2 FILLER_22_731 ();
 sg13g2_fill_2 FILLER_22_758 ();
 sg13g2_fill_1 FILLER_22_760 ();
 sg13g2_decap_4 FILLER_22_765 ();
 sg13g2_fill_1 FILLER_22_809 ();
 sg13g2_fill_2 FILLER_22_898 ();
 sg13g2_fill_1 FILLER_22_900 ();
 sg13g2_fill_2 FILLER_22_937 ();
 sg13g2_fill_2 FILLER_22_1003 ();
 sg13g2_fill_1 FILLER_22_1005 ();
 sg13g2_fill_1 FILLER_22_1029 ();
 sg13g2_decap_4 FILLER_22_1093 ();
 sg13g2_fill_1 FILLER_22_1097 ();
 sg13g2_fill_1 FILLER_22_1135 ();
 sg13g2_fill_2 FILLER_22_1306 ();
 sg13g2_fill_2 FILLER_22_1325 ();
 sg13g2_fill_1 FILLER_22_1327 ();
 sg13g2_fill_2 FILLER_22_1341 ();
 sg13g2_fill_2 FILLER_22_1369 ();
 sg13g2_fill_2 FILLER_22_1495 ();
 sg13g2_fill_2 FILLER_22_1506 ();
 sg13g2_fill_1 FILLER_22_1521 ();
 sg13g2_fill_1 FILLER_22_1609 ();
 sg13g2_fill_1 FILLER_22_1704 ();
 sg13g2_fill_1 FILLER_22_1709 ();
 sg13g2_decap_8 FILLER_22_1761 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_fill_2 FILLER_23_17 ();
 sg13g2_fill_1 FILLER_23_19 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_fill_2 FILLER_23_58 ();
 sg13g2_fill_1 FILLER_23_60 ();
 sg13g2_decap_4 FILLER_23_100 ();
 sg13g2_fill_2 FILLER_23_107 ();
 sg13g2_fill_1 FILLER_23_127 ();
 sg13g2_decap_8 FILLER_23_141 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_150 ();
 sg13g2_fill_2 FILLER_23_222 ();
 sg13g2_decap_4 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_305 ();
 sg13g2_decap_4 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_fill_1 FILLER_23_350 ();
 sg13g2_fill_2 FILLER_23_370 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_fill_2 FILLER_23_430 ();
 sg13g2_fill_1 FILLER_23_432 ();
 sg13g2_decap_8 FILLER_23_456 ();
 sg13g2_decap_8 FILLER_23_463 ();
 sg13g2_fill_2 FILLER_23_492 ();
 sg13g2_fill_1 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_fill_2 FILLER_23_553 ();
 sg13g2_fill_1 FILLER_23_580 ();
 sg13g2_decap_4 FILLER_23_608 ();
 sg13g2_fill_1 FILLER_23_612 ();
 sg13g2_fill_2 FILLER_23_677 ();
 sg13g2_fill_1 FILLER_23_679 ();
 sg13g2_fill_2 FILLER_23_701 ();
 sg13g2_fill_1 FILLER_23_703 ();
 sg13g2_fill_1 FILLER_23_708 ();
 sg13g2_fill_2 FILLER_23_720 ();
 sg13g2_fill_2 FILLER_23_744 ();
 sg13g2_decap_8 FILLER_23_772 ();
 sg13g2_fill_1 FILLER_23_779 ();
 sg13g2_fill_2 FILLER_23_801 ();
 sg13g2_fill_2 FILLER_23_807 ();
 sg13g2_fill_1 FILLER_23_826 ();
 sg13g2_fill_1 FILLER_23_868 ();
 sg13g2_decap_4 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_896 ();
 sg13g2_decap_4 FILLER_23_903 ();
 sg13g2_decap_4 FILLER_23_911 ();
 sg13g2_fill_1 FILLER_23_915 ();
 sg13g2_fill_2 FILLER_23_969 ();
 sg13g2_fill_1 FILLER_23_971 ();
 sg13g2_fill_1 FILLER_23_976 ();
 sg13g2_decap_8 FILLER_23_1008 ();
 sg13g2_fill_1 FILLER_23_1015 ();
 sg13g2_fill_2 FILLER_23_1096 ();
 sg13g2_fill_1 FILLER_23_1151 ();
 sg13g2_fill_1 FILLER_23_1188 ();
 sg13g2_fill_1 FILLER_23_1211 ();
 sg13g2_fill_1 FILLER_23_1257 ();
 sg13g2_fill_2 FILLER_23_1287 ();
 sg13g2_fill_1 FILLER_23_1289 ();
 sg13g2_fill_2 FILLER_23_1452 ();
 sg13g2_fill_1 FILLER_23_1472 ();
 sg13g2_fill_2 FILLER_23_1546 ();
 sg13g2_fill_1 FILLER_23_1560 ();
 sg13g2_fill_1 FILLER_23_1590 ();
 sg13g2_fill_1 FILLER_23_1616 ();
 sg13g2_fill_1 FILLER_23_1693 ();
 sg13g2_fill_2 FILLER_23_1721 ();
 sg13g2_fill_2 FILLER_23_1766 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_fill_2 FILLER_24_52 ();
 sg13g2_fill_2 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_83 ();
 sg13g2_fill_1 FILLER_24_90 ();
 sg13g2_fill_1 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_121 ();
 sg13g2_fill_1 FILLER_24_138 ();
 sg13g2_fill_1 FILLER_24_149 ();
 sg13g2_fill_2 FILLER_24_155 ();
 sg13g2_decap_4 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_decap_4 FILLER_24_176 ();
 sg13g2_fill_2 FILLER_24_180 ();
 sg13g2_fill_1 FILLER_24_186 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_decap_4 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_fill_2 FILLER_24_246 ();
 sg13g2_fill_1 FILLER_24_248 ();
 sg13g2_fill_1 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_289 ();
 sg13g2_fill_1 FILLER_24_291 ();
 sg13g2_decap_4 FILLER_24_310 ();
 sg13g2_decap_4 FILLER_24_319 ();
 sg13g2_fill_2 FILLER_24_323 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_fill_2 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_370 ();
 sg13g2_decap_4 FILLER_24_398 ();
 sg13g2_fill_2 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_fill_1 FILLER_24_459 ();
 sg13g2_fill_2 FILLER_24_474 ();
 sg13g2_fill_1 FILLER_24_476 ();
 sg13g2_decap_4 FILLER_24_495 ();
 sg13g2_decap_4 FILLER_24_504 ();
 sg13g2_fill_1 FILLER_24_508 ();
 sg13g2_fill_2 FILLER_24_513 ();
 sg13g2_fill_1 FILLER_24_515 ();
 sg13g2_fill_2 FILLER_24_525 ();
 sg13g2_fill_1 FILLER_24_527 ();
 sg13g2_decap_4 FILLER_24_571 ();
 sg13g2_fill_1 FILLER_24_580 ();
 sg13g2_decap_8 FILLER_24_602 ();
 sg13g2_decap_4 FILLER_24_609 ();
 sg13g2_fill_1 FILLER_24_613 ();
 sg13g2_decap_8 FILLER_24_622 ();
 sg13g2_fill_2 FILLER_24_629 ();
 sg13g2_fill_2 FILLER_24_641 ();
 sg13g2_decap_4 FILLER_24_647 ();
 sg13g2_fill_2 FILLER_24_685 ();
 sg13g2_fill_1 FILLER_24_687 ();
 sg13g2_fill_2 FILLER_24_692 ();
 sg13g2_fill_2 FILLER_24_698 ();
 sg13g2_fill_1 FILLER_24_700 ();
 sg13g2_fill_2 FILLER_24_718 ();
 sg13g2_fill_1 FILLER_24_720 ();
 sg13g2_fill_1 FILLER_24_735 ();
 sg13g2_fill_1 FILLER_24_756 ();
 sg13g2_fill_1 FILLER_24_780 ();
 sg13g2_fill_2 FILLER_24_801 ();
 sg13g2_fill_1 FILLER_24_835 ();
 sg13g2_fill_1 FILLER_24_862 ();
 sg13g2_decap_8 FILLER_24_877 ();
 sg13g2_fill_2 FILLER_24_884 ();
 sg13g2_fill_1 FILLER_24_886 ();
 sg13g2_decap_4 FILLER_24_915 ();
 sg13g2_fill_2 FILLER_24_919 ();
 sg13g2_fill_2 FILLER_24_969 ();
 sg13g2_fill_1 FILLER_24_971 ();
 sg13g2_fill_2 FILLER_24_989 ();
 sg13g2_fill_1 FILLER_24_991 ();
 sg13g2_fill_2 FILLER_24_1072 ();
 sg13g2_fill_1 FILLER_24_1074 ();
 sg13g2_fill_1 FILLER_24_1120 ();
 sg13g2_fill_2 FILLER_24_1169 ();
 sg13g2_fill_2 FILLER_24_1225 ();
 sg13g2_fill_1 FILLER_24_1282 ();
 sg13g2_fill_1 FILLER_24_1357 ();
 sg13g2_fill_2 FILLER_24_1394 ();
 sg13g2_fill_1 FILLER_24_1457 ();
 sg13g2_fill_2 FILLER_24_1531 ();
 sg13g2_fill_1 FILLER_24_1581 ();
 sg13g2_fill_1 FILLER_24_1588 ();
 sg13g2_fill_1 FILLER_24_1616 ();
 sg13g2_fill_2 FILLER_24_1672 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_fill_1 FILLER_25_20 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_fill_2 FILLER_25_131 ();
 sg13g2_decap_4 FILLER_25_141 ();
 sg13g2_decap_4 FILLER_25_164 ();
 sg13g2_fill_1 FILLER_25_173 ();
 sg13g2_fill_1 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_251 ();
 sg13g2_fill_2 FILLER_25_258 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_287 ();
 sg13g2_fill_1 FILLER_25_312 ();
 sg13g2_fill_2 FILLER_25_336 ();
 sg13g2_fill_1 FILLER_25_338 ();
 sg13g2_fill_2 FILLER_25_346 ();
 sg13g2_fill_2 FILLER_25_379 ();
 sg13g2_fill_2 FILLER_25_385 ();
 sg13g2_fill_1 FILLER_25_387 ();
 sg13g2_decap_4 FILLER_25_393 ();
 sg13g2_fill_2 FILLER_25_397 ();
 sg13g2_fill_1 FILLER_25_421 ();
 sg13g2_fill_2 FILLER_25_450 ();
 sg13g2_fill_2 FILLER_25_484 ();
 sg13g2_fill_1 FILLER_25_583 ();
 sg13g2_decap_4 FILLER_25_604 ();
 sg13g2_fill_1 FILLER_25_608 ();
 sg13g2_fill_2 FILLER_25_641 ();
 sg13g2_fill_1 FILLER_25_643 ();
 sg13g2_fill_2 FILLER_25_657 ();
 sg13g2_fill_1 FILLER_25_664 ();
 sg13g2_decap_4 FILLER_25_669 ();
 sg13g2_fill_1 FILLER_25_718 ();
 sg13g2_fill_2 FILLER_25_746 ();
 sg13g2_fill_1 FILLER_25_748 ();
 sg13g2_fill_1 FILLER_25_795 ();
 sg13g2_fill_2 FILLER_25_817 ();
 sg13g2_fill_2 FILLER_25_870 ();
 sg13g2_fill_1 FILLER_25_876 ();
 sg13g2_decap_8 FILLER_25_886 ();
 sg13g2_fill_2 FILLER_25_974 ();
 sg13g2_fill_1 FILLER_25_976 ();
 sg13g2_fill_2 FILLER_25_1005 ();
 sg13g2_fill_1 FILLER_25_1024 ();
 sg13g2_fill_2 FILLER_25_1038 ();
 sg13g2_fill_1 FILLER_25_1040 ();
 sg13g2_fill_2 FILLER_25_1099 ();
 sg13g2_fill_1 FILLER_25_1180 ();
 sg13g2_fill_2 FILLER_25_1248 ();
 sg13g2_fill_1 FILLER_25_1336 ();
 sg13g2_fill_1 FILLER_25_1376 ();
 sg13g2_fill_2 FILLER_25_1408 ();
 sg13g2_fill_1 FILLER_25_1473 ();
 sg13g2_fill_2 FILLER_25_1504 ();
 sg13g2_fill_1 FILLER_25_1555 ();
 sg13g2_fill_1 FILLER_25_1580 ();
 sg13g2_fill_2 FILLER_25_1587 ();
 sg13g2_fill_2 FILLER_25_1605 ();
 sg13g2_fill_2 FILLER_25_1734 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_97 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_142 ();
 sg13g2_fill_1 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_168 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_fill_2 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_4 FILLER_26_328 ();
 sg13g2_fill_2 FILLER_26_350 ();
 sg13g2_fill_1 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_434 ();
 sg13g2_fill_1 FILLER_26_443 ();
 sg13g2_fill_2 FILLER_26_482 ();
 sg13g2_fill_1 FILLER_26_484 ();
 sg13g2_decap_4 FILLER_26_495 ();
 sg13g2_fill_2 FILLER_26_499 ();
 sg13g2_decap_8 FILLER_26_509 ();
 sg13g2_fill_2 FILLER_26_516 ();
 sg13g2_decap_4 FILLER_26_522 ();
 sg13g2_fill_2 FILLER_26_526 ();
 sg13g2_fill_2 FILLER_26_553 ();
 sg13g2_fill_2 FILLER_26_609 ();
 sg13g2_fill_2 FILLER_26_631 ();
 sg13g2_fill_1 FILLER_26_697 ();
 sg13g2_fill_1 FILLER_26_723 ();
 sg13g2_fill_2 FILLER_26_728 ();
 sg13g2_fill_1 FILLER_26_730 ();
 sg13g2_fill_1 FILLER_26_766 ();
 sg13g2_fill_1 FILLER_26_793 ();
 sg13g2_fill_2 FILLER_26_832 ();
 sg13g2_fill_1 FILLER_26_843 ();
 sg13g2_decap_4 FILLER_26_911 ();
 sg13g2_fill_1 FILLER_26_915 ();
 sg13g2_fill_1 FILLER_26_1001 ();
 sg13g2_fill_1 FILLER_26_1057 ();
 sg13g2_fill_2 FILLER_26_1094 ();
 sg13g2_fill_1 FILLER_26_1122 ();
 sg13g2_fill_2 FILLER_26_1141 ();
 sg13g2_fill_2 FILLER_26_1197 ();
 sg13g2_fill_1 FILLER_26_1199 ();
 sg13g2_fill_1 FILLER_26_1260 ();
 sg13g2_fill_2 FILLER_26_1282 ();
 sg13g2_fill_2 FILLER_26_1341 ();
 sg13g2_fill_1 FILLER_26_1396 ();
 sg13g2_fill_1 FILLER_26_1405 ();
 sg13g2_fill_2 FILLER_26_1473 ();
 sg13g2_fill_1 FILLER_26_1475 ();
 sg13g2_fill_1 FILLER_26_1494 ();
 sg13g2_fill_2 FILLER_26_1520 ();
 sg13g2_fill_2 FILLER_26_1554 ();
 sg13g2_fill_2 FILLER_26_1588 ();
 sg13g2_fill_1 FILLER_26_1633 ();
 sg13g2_fill_2 FILLER_26_1704 ();
 sg13g2_fill_2 FILLER_26_1744 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_63 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_2 FILLER_27_80 ();
 sg13g2_fill_1 FILLER_27_82 ();
 sg13g2_fill_2 FILLER_27_93 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_118 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_143 ();
 sg13g2_fill_1 FILLER_27_145 ();
 sg13g2_fill_1 FILLER_27_183 ();
 sg13g2_fill_2 FILLER_27_201 ();
 sg13g2_fill_1 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_230 ();
 sg13g2_decap_4 FILLER_27_243 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_decap_8 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_2 FILLER_27_285 ();
 sg13g2_fill_1 FILLER_27_287 ();
 sg13g2_decap_4 FILLER_27_316 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_decap_4 FILLER_27_356 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_decap_4 FILLER_27_384 ();
 sg13g2_fill_2 FILLER_27_388 ();
 sg13g2_fill_2 FILLER_27_424 ();
 sg13g2_decap_4 FILLER_27_489 ();
 sg13g2_decap_4 FILLER_27_511 ();
 sg13g2_fill_2 FILLER_27_515 ();
 sg13g2_fill_2 FILLER_27_661 ();
 sg13g2_fill_1 FILLER_27_663 ();
 sg13g2_decap_4 FILLER_27_668 ();
 sg13g2_fill_1 FILLER_27_672 ();
 sg13g2_fill_1 FILLER_27_695 ();
 sg13g2_fill_1 FILLER_27_716 ();
 sg13g2_decap_8 FILLER_27_730 ();
 sg13g2_fill_2 FILLER_27_737 ();
 sg13g2_decap_4 FILLER_27_748 ();
 sg13g2_fill_1 FILLER_27_752 ();
 sg13g2_fill_1 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_922 ();
 sg13g2_fill_1 FILLER_27_929 ();
 sg13g2_fill_2 FILLER_27_963 ();
 sg13g2_fill_1 FILLER_27_965 ();
 sg13g2_fill_1 FILLER_27_976 ();
 sg13g2_fill_1 FILLER_27_1025 ();
 sg13g2_fill_2 FILLER_27_1067 ();
 sg13g2_fill_1 FILLER_27_1069 ();
 sg13g2_fill_1 FILLER_27_1178 ();
 sg13g2_fill_1 FILLER_27_1269 ();
 sg13g2_fill_2 FILLER_27_1274 ();
 sg13g2_fill_1 FILLER_27_1332 ();
 sg13g2_fill_2 FILLER_27_1462 ();
 sg13g2_fill_1 FILLER_27_1512 ();
 sg13g2_fill_2 FILLER_27_1517 ();
 sg13g2_fill_1 FILLER_27_1538 ();
 sg13g2_fill_1 FILLER_27_1588 ();
 sg13g2_fill_1 FILLER_27_1616 ();
 sg13g2_fill_2 FILLER_27_1705 ();
 sg13g2_fill_2 FILLER_27_1739 ();
 sg13g2_fill_1 FILLER_28_18 ();
 sg13g2_fill_1 FILLER_28_90 ();
 sg13g2_fill_2 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_107 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_222 ();
 sg13g2_fill_1 FILLER_28_224 ();
 sg13g2_decap_4 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_257 ();
 sg13g2_decap_8 FILLER_28_286 ();
 sg13g2_decap_4 FILLER_28_293 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_fill_2 FILLER_28_356 ();
 sg13g2_fill_1 FILLER_28_394 ();
 sg13g2_fill_1 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_449 ();
 sg13g2_fill_2 FILLER_28_459 ();
 sg13g2_fill_2 FILLER_28_475 ();
 sg13g2_decap_4 FILLER_28_494 ();
 sg13g2_fill_2 FILLER_28_504 ();
 sg13g2_fill_1 FILLER_28_506 ();
 sg13g2_decap_4 FILLER_28_512 ();
 sg13g2_fill_2 FILLER_28_547 ();
 sg13g2_fill_2 FILLER_28_567 ();
 sg13g2_fill_1 FILLER_28_569 ();
 sg13g2_fill_2 FILLER_28_575 ();
 sg13g2_fill_2 FILLER_28_679 ();
 sg13g2_decap_4 FILLER_28_697 ();
 sg13g2_fill_1 FILLER_28_701 ();
 sg13g2_decap_4 FILLER_28_750 ();
 sg13g2_fill_1 FILLER_28_754 ();
 sg13g2_fill_2 FILLER_28_769 ();
 sg13g2_fill_1 FILLER_28_771 ();
 sg13g2_fill_2 FILLER_28_787 ();
 sg13g2_fill_1 FILLER_28_802 ();
 sg13g2_fill_1 FILLER_28_854 ();
 sg13g2_fill_1 FILLER_28_883 ();
 sg13g2_decap_4 FILLER_28_898 ();
 sg13g2_fill_1 FILLER_28_902 ();
 sg13g2_fill_2 FILLER_28_951 ();
 sg13g2_fill_1 FILLER_28_953 ();
 sg13g2_fill_1 FILLER_28_976 ();
 sg13g2_fill_2 FILLER_28_1053 ();
 sg13g2_fill_1 FILLER_28_1055 ();
 sg13g2_fill_1 FILLER_28_1075 ();
 sg13g2_fill_2 FILLER_28_1148 ();
 sg13g2_fill_1 FILLER_28_1150 ();
 sg13g2_fill_2 FILLER_28_1178 ();
 sg13g2_fill_1 FILLER_28_1207 ();
 sg13g2_fill_2 FILLER_28_1262 ();
 sg13g2_fill_1 FILLER_28_1264 ();
 sg13g2_fill_1 FILLER_28_1351 ();
 sg13g2_fill_1 FILLER_28_1432 ();
 sg13g2_fill_2 FILLER_28_1452 ();
 sg13g2_fill_2 FILLER_28_1467 ();
 sg13g2_fill_1 FILLER_28_1568 ();
 sg13g2_fill_1 FILLER_28_1678 ();
 sg13g2_fill_2 FILLER_28_1687 ();
 sg13g2_fill_1 FILLER_28_1702 ();
 sg13g2_decap_4 FILLER_28_1764 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_54 ();
 sg13g2_fill_1 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_75 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_212 ();
 sg13g2_fill_1 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_247 ();
 sg13g2_decap_8 FILLER_29_254 ();
 sg13g2_fill_1 FILLER_29_261 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_318 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_393 ();
 sg13g2_fill_2 FILLER_29_435 ();
 sg13g2_fill_2 FILLER_29_446 ();
 sg13g2_fill_1 FILLER_29_448 ();
 sg13g2_fill_1 FILLER_29_499 ();
 sg13g2_fill_2 FILLER_29_504 ();
 sg13g2_decap_4 FILLER_29_511 ();
 sg13g2_fill_2 FILLER_29_528 ();
 sg13g2_decap_4 FILLER_29_545 ();
 sg13g2_fill_2 FILLER_29_558 ();
 sg13g2_fill_1 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_fill_2 FILLER_29_599 ();
 sg13g2_fill_2 FILLER_29_614 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_fill_2 FILLER_29_640 ();
 sg13g2_fill_1 FILLER_29_642 ();
 sg13g2_decap_8 FILLER_29_647 ();
 sg13g2_fill_1 FILLER_29_654 ();
 sg13g2_decap_4 FILLER_29_663 ();
 sg13g2_fill_2 FILLER_29_742 ();
 sg13g2_decap_4 FILLER_29_760 ();
 sg13g2_fill_1 FILLER_29_764 ();
 sg13g2_fill_1 FILLER_29_769 ();
 sg13g2_fill_1 FILLER_29_787 ();
 sg13g2_fill_2 FILLER_29_794 ();
 sg13g2_fill_1 FILLER_29_796 ();
 sg13g2_fill_2 FILLER_29_841 ();
 sg13g2_fill_1 FILLER_29_901 ();
 sg13g2_fill_1 FILLER_29_1090 ();
 sg13g2_fill_2 FILLER_29_1233 ();
 sg13g2_fill_2 FILLER_29_1261 ();
 sg13g2_fill_1 FILLER_29_1263 ();
 sg13g2_fill_1 FILLER_29_1291 ();
 sg13g2_fill_1 FILLER_29_1333 ();
 sg13g2_fill_1 FILLER_29_1369 ();
 sg13g2_fill_2 FILLER_29_1383 ();
 sg13g2_fill_2 FILLER_29_1429 ();
 sg13g2_fill_2 FILLER_29_1557 ();
 sg13g2_fill_2 FILLER_29_1673 ();
 sg13g2_fill_2 FILLER_29_1679 ();
 sg13g2_fill_2 FILLER_29_1685 ();
 sg13g2_fill_1 FILLER_29_1739 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_82 ();
 sg13g2_fill_2 FILLER_30_117 ();
 sg13g2_fill_2 FILLER_30_129 ();
 sg13g2_fill_1 FILLER_30_131 ();
 sg13g2_fill_1 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_175 ();
 sg13g2_fill_2 FILLER_30_194 ();
 sg13g2_fill_1 FILLER_30_209 ();
 sg13g2_decap_4 FILLER_30_229 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_325 ();
 sg13g2_fill_1 FILLER_30_327 ();
 sg13g2_fill_2 FILLER_30_342 ();
 sg13g2_fill_2 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_396 ();
 sg13g2_fill_1 FILLER_30_406 ();
 sg13g2_fill_2 FILLER_30_452 ();
 sg13g2_fill_1 FILLER_30_466 ();
 sg13g2_fill_2 FILLER_30_476 ();
 sg13g2_fill_1 FILLER_30_478 ();
 sg13g2_fill_2 FILLER_30_491 ();
 sg13g2_fill_2 FILLER_30_501 ();
 sg13g2_fill_2 FILLER_30_534 ();
 sg13g2_fill_1 FILLER_30_564 ();
 sg13g2_fill_1 FILLER_30_667 ();
 sg13g2_fill_1 FILLER_30_691 ();
 sg13g2_fill_1 FILLER_30_705 ();
 sg13g2_fill_2 FILLER_30_718 ();
 sg13g2_fill_1 FILLER_30_732 ();
 sg13g2_fill_2 FILLER_30_803 ();
 sg13g2_fill_1 FILLER_30_805 ();
 sg13g2_fill_1 FILLER_30_838 ();
 sg13g2_decap_4 FILLER_30_934 ();
 sg13g2_fill_1 FILLER_30_951 ();
 sg13g2_fill_1 FILLER_30_1006 ();
 sg13g2_fill_2 FILLER_30_1021 ();
 sg13g2_fill_1 FILLER_30_1023 ();
 sg13g2_fill_2 FILLER_30_1033 ();
 sg13g2_fill_1 FILLER_30_1035 ();
 sg13g2_fill_2 FILLER_30_1087 ();
 sg13g2_fill_1 FILLER_30_1102 ();
 sg13g2_fill_2 FILLER_30_1112 ();
 sg13g2_fill_1 FILLER_30_1114 ();
 sg13g2_fill_2 FILLER_30_1155 ();
 sg13g2_fill_1 FILLER_30_1157 ();
 sg13g2_fill_1 FILLER_30_1300 ();
 sg13g2_fill_1 FILLER_30_1368 ();
 sg13g2_fill_2 FILLER_30_1434 ();
 sg13g2_fill_1 FILLER_30_1472 ();
 sg13g2_fill_1 FILLER_30_1477 ();
 sg13g2_fill_1 FILLER_30_1497 ();
 sg13g2_fill_1 FILLER_30_1536 ();
 sg13g2_fill_1 FILLER_30_1572 ();
 sg13g2_fill_2 FILLER_30_1578 ();
 sg13g2_fill_2 FILLER_30_1593 ();
 sg13g2_fill_1 FILLER_30_1608 ();
 sg13g2_fill_2 FILLER_30_1644 ();
 sg13g2_decap_8 FILLER_30_1660 ();
 sg13g2_fill_1 FILLER_30_1667 ();
 sg13g2_fill_1 FILLER_30_1751 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_fill_2 FILLER_31_30 ();
 sg13g2_fill_1 FILLER_31_32 ();
 sg13g2_fill_2 FILLER_31_80 ();
 sg13g2_fill_2 FILLER_31_96 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_decap_4 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_270 ();
 sg13g2_fill_2 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_291 ();
 sg13g2_fill_1 FILLER_31_302 ();
 sg13g2_fill_2 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_decap_4 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_fill_2 FILLER_31_399 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_fill_2 FILLER_31_425 ();
 sg13g2_fill_2 FILLER_31_435 ();
 sg13g2_fill_1 FILLER_31_441 ();
 sg13g2_fill_1 FILLER_31_448 ();
 sg13g2_decap_4 FILLER_31_470 ();
 sg13g2_decap_4 FILLER_31_485 ();
 sg13g2_decap_4 FILLER_31_506 ();
 sg13g2_fill_2 FILLER_31_518 ();
 sg13g2_fill_1 FILLER_31_520 ();
 sg13g2_fill_1 FILLER_31_531 ();
 sg13g2_fill_2 FILLER_31_537 ();
 sg13g2_fill_1 FILLER_31_539 ();
 sg13g2_fill_2 FILLER_31_543 ();
 sg13g2_fill_1 FILLER_31_545 ();
 sg13g2_fill_1 FILLER_31_550 ();
 sg13g2_fill_2 FILLER_31_565 ();
 sg13g2_fill_1 FILLER_31_567 ();
 sg13g2_fill_1 FILLER_31_580 ();
 sg13g2_fill_1 FILLER_31_594 ();
 sg13g2_fill_2 FILLER_31_623 ();
 sg13g2_fill_1 FILLER_31_625 ();
 sg13g2_fill_1 FILLER_31_643 ();
 sg13g2_fill_2 FILLER_31_648 ();
 sg13g2_fill_2 FILLER_31_682 ();
 sg13g2_fill_2 FILLER_31_725 ();
 sg13g2_fill_1 FILLER_31_727 ();
 sg13g2_fill_1 FILLER_31_735 ();
 sg13g2_fill_2 FILLER_31_746 ();
 sg13g2_fill_1 FILLER_31_780 ();
 sg13g2_fill_1 FILLER_31_798 ();
 sg13g2_fill_2 FILLER_31_803 ();
 sg13g2_fill_2 FILLER_31_828 ();
 sg13g2_fill_2 FILLER_31_870 ();
 sg13g2_fill_1 FILLER_31_872 ();
 sg13g2_fill_2 FILLER_31_913 ();
 sg13g2_fill_1 FILLER_31_957 ();
 sg13g2_fill_2 FILLER_31_995 ();
 sg13g2_fill_1 FILLER_31_997 ();
 sg13g2_fill_2 FILLER_31_1052 ();
 sg13g2_fill_1 FILLER_31_1054 ();
 sg13g2_fill_1 FILLER_31_1064 ();
 sg13g2_fill_1 FILLER_31_1138 ();
 sg13g2_fill_2 FILLER_31_1193 ();
 sg13g2_fill_1 FILLER_31_1195 ();
 sg13g2_fill_1 FILLER_31_1214 ();
 sg13g2_fill_2 FILLER_31_1232 ();
 sg13g2_fill_1 FILLER_31_1234 ();
 sg13g2_fill_2 FILLER_31_1244 ();
 sg13g2_fill_2 FILLER_31_1321 ();
 sg13g2_fill_2 FILLER_31_1335 ();
 sg13g2_fill_2 FILLER_31_1361 ();
 sg13g2_fill_1 FILLER_31_1438 ();
 sg13g2_fill_2 FILLER_31_1452 ();
 sg13g2_fill_1 FILLER_31_1489 ();
 sg13g2_fill_1 FILLER_31_1541 ();
 sg13g2_fill_1 FILLER_31_1594 ();
 sg13g2_fill_2 FILLER_31_1599 ();
 sg13g2_fill_2 FILLER_31_1648 ();
 sg13g2_decap_8 FILLER_31_1677 ();
 sg13g2_decap_8 FILLER_31_1684 ();
 sg13g2_fill_2 FILLER_31_1691 ();
 sg13g2_fill_1 FILLER_31_1693 ();
 sg13g2_fill_1 FILLER_31_1756 ();
 sg13g2_fill_2 FILLER_31_1766 ();
 sg13g2_fill_2 FILLER_32_56 ();
 sg13g2_fill_1 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_132 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_156 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_decap_4 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_225 ();
 sg13g2_fill_1 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_275 ();
 sg13g2_decap_4 FILLER_32_282 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_decap_4 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_fill_2 FILLER_32_393 ();
 sg13g2_fill_1 FILLER_32_427 ();
 sg13g2_decap_8 FILLER_32_458 ();
 sg13g2_fill_1 FILLER_32_465 ();
 sg13g2_fill_2 FILLER_32_470 ();
 sg13g2_fill_1 FILLER_32_477 ();
 sg13g2_decap_8 FILLER_32_505 ();
 sg13g2_fill_1 FILLER_32_512 ();
 sg13g2_decap_4 FILLER_32_541 ();
 sg13g2_fill_1 FILLER_32_550 ();
 sg13g2_fill_1 FILLER_32_593 ();
 sg13g2_fill_2 FILLER_32_608 ();
 sg13g2_fill_1 FILLER_32_610 ();
 sg13g2_fill_2 FILLER_32_647 ();
 sg13g2_fill_2 FILLER_32_689 ();
 sg13g2_fill_1 FILLER_32_691 ();
 sg13g2_fill_2 FILLER_32_696 ();
 sg13g2_fill_1 FILLER_32_698 ();
 sg13g2_fill_1 FILLER_32_731 ();
 sg13g2_fill_2 FILLER_32_753 ();
 sg13g2_fill_1 FILLER_32_755 ();
 sg13g2_decap_4 FILLER_32_769 ();
 sg13g2_fill_2 FILLER_32_773 ();
 sg13g2_fill_1 FILLER_32_843 ();
 sg13g2_fill_1 FILLER_32_867 ();
 sg13g2_fill_2 FILLER_32_878 ();
 sg13g2_fill_1 FILLER_32_880 ();
 sg13g2_decap_4 FILLER_32_894 ();
 sg13g2_fill_1 FILLER_32_898 ();
 sg13g2_decap_4 FILLER_32_903 ();
 sg13g2_fill_2 FILLER_32_948 ();
 sg13g2_fill_2 FILLER_32_963 ();
 sg13g2_fill_1 FILLER_32_965 ();
 sg13g2_decap_4 FILLER_32_989 ();
 sg13g2_fill_1 FILLER_32_993 ();
 sg13g2_fill_1 FILLER_32_1015 ();
 sg13g2_fill_2 FILLER_32_1020 ();
 sg13g2_fill_1 FILLER_32_1090 ();
 sg13g2_fill_2 FILLER_32_1100 ();
 sg13g2_fill_2 FILLER_32_1151 ();
 sg13g2_fill_1 FILLER_32_1346 ();
 sg13g2_fill_2 FILLER_32_1379 ();
 sg13g2_fill_1 FILLER_32_1381 ();
 sg13g2_decap_4 FILLER_32_1388 ();
 sg13g2_fill_2 FILLER_32_1455 ();
 sg13g2_fill_2 FILLER_32_1481 ();
 sg13g2_fill_1 FILLER_32_1493 ();
 sg13g2_fill_1 FILLER_32_1675 ();
 sg13g2_fill_2 FILLER_32_1685 ();
 sg13g2_fill_1 FILLER_32_1687 ();
 sg13g2_fill_2 FILLER_33_38 ();
 sg13g2_fill_2 FILLER_33_89 ();
 sg13g2_fill_2 FILLER_33_154 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_4 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_280 ();
 sg13g2_fill_1 FILLER_33_298 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_336 ();
 sg13g2_fill_2 FILLER_33_354 ();
 sg13g2_fill_1 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_375 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_412 ();
 sg13g2_fill_2 FILLER_33_419 ();
 sg13g2_fill_1 FILLER_33_454 ();
 sg13g2_decap_8 FILLER_33_481 ();
 sg13g2_decap_4 FILLER_33_510 ();
 sg13g2_fill_2 FILLER_33_514 ();
 sg13g2_fill_2 FILLER_33_520 ();
 sg13g2_fill_1 FILLER_33_522 ();
 sg13g2_fill_2 FILLER_33_541 ();
 sg13g2_fill_1 FILLER_33_543 ();
 sg13g2_fill_2 FILLER_33_567 ();
 sg13g2_fill_2 FILLER_33_573 ();
 sg13g2_fill_1 FILLER_33_575 ();
 sg13g2_fill_2 FILLER_33_598 ();
 sg13g2_fill_1 FILLER_33_615 ();
 sg13g2_decap_4 FILLER_33_620 ();
 sg13g2_fill_2 FILLER_33_637 ();
 sg13g2_decap_4 FILLER_33_736 ();
 sg13g2_decap_4 FILLER_33_777 ();
 sg13g2_fill_1 FILLER_33_781 ();
 sg13g2_decap_4 FILLER_33_817 ();
 sg13g2_fill_2 FILLER_33_821 ();
 sg13g2_fill_2 FILLER_33_855 ();
 sg13g2_fill_1 FILLER_33_857 ();
 sg13g2_fill_2 FILLER_33_944 ();
 sg13g2_fill_1 FILLER_33_1008 ();
 sg13g2_fill_1 FILLER_33_1021 ();
 sg13g2_fill_2 FILLER_33_1038 ();
 sg13g2_fill_2 FILLER_33_1079 ();
 sg13g2_fill_2 FILLER_33_1112 ();
 sg13g2_fill_1 FILLER_33_1227 ();
 sg13g2_fill_1 FILLER_33_1248 ();
 sg13g2_fill_2 FILLER_33_1267 ();
 sg13g2_fill_1 FILLER_33_1425 ();
 sg13g2_fill_1 FILLER_33_1479 ();
 sg13g2_fill_2 FILLER_33_1513 ();
 sg13g2_fill_2 FILLER_33_1535 ();
 sg13g2_fill_2 FILLER_33_1597 ();
 sg13g2_fill_2 FILLER_33_1647 ();
 sg13g2_fill_1 FILLER_33_1685 ();
 sg13g2_fill_2 FILLER_33_1690 ();
 sg13g2_fill_2 FILLER_33_1730 ();
 sg13g2_fill_1 FILLER_33_1767 ();
 sg13g2_fill_2 FILLER_34_31 ();
 sg13g2_fill_1 FILLER_34_33 ();
 sg13g2_fill_2 FILLER_34_71 ();
 sg13g2_fill_1 FILLER_34_73 ();
 sg13g2_fill_2 FILLER_34_98 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_121 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_1 FILLER_34_269 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_309 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_fill_2 FILLER_34_342 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_fill_1 FILLER_34_350 ();
 sg13g2_fill_2 FILLER_34_383 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_fill_1 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_34_430 ();
 sg13g2_fill_2 FILLER_34_448 ();
 sg13g2_decap_4 FILLER_34_492 ();
 sg13g2_decap_4 FILLER_34_504 ();
 sg13g2_decap_8 FILLER_34_518 ();
 sg13g2_decap_8 FILLER_34_525 ();
 sg13g2_decap_4 FILLER_34_532 ();
 sg13g2_fill_2 FILLER_34_536 ();
 sg13g2_fill_1 FILLER_34_557 ();
 sg13g2_decap_4 FILLER_34_567 ();
 sg13g2_fill_2 FILLER_34_598 ();
 sg13g2_fill_1 FILLER_34_619 ();
 sg13g2_decap_4 FILLER_34_723 ();
 sg13g2_fill_2 FILLER_34_727 ();
 sg13g2_decap_8 FILLER_34_750 ();
 sg13g2_fill_1 FILLER_34_757 ();
 sg13g2_fill_2 FILLER_34_770 ();
 sg13g2_fill_2 FILLER_34_782 ();
 sg13g2_fill_2 FILLER_34_825 ();
 sg13g2_fill_1 FILLER_34_827 ();
 sg13g2_fill_2 FILLER_34_832 ();
 sg13g2_decap_4 FILLER_34_869 ();
 sg13g2_fill_1 FILLER_34_881 ();
 sg13g2_fill_2 FILLER_34_886 ();
 sg13g2_fill_2 FILLER_34_896 ();
 sg13g2_fill_1 FILLER_34_898 ();
 sg13g2_fill_2 FILLER_34_940 ();
 sg13g2_decap_8 FILLER_34_970 ();
 sg13g2_decap_4 FILLER_34_977 ();
 sg13g2_fill_2 FILLER_34_1070 ();
 sg13g2_fill_2 FILLER_34_1090 ();
 sg13g2_fill_1 FILLER_34_1201 ();
 sg13g2_fill_2 FILLER_34_1302 ();
 sg13g2_fill_1 FILLER_34_1337 ();
 sg13g2_fill_1 FILLER_34_1363 ();
 sg13g2_fill_2 FILLER_34_1386 ();
 sg13g2_decap_4 FILLER_34_1424 ();
 sg13g2_fill_1 FILLER_34_1480 ();
 sg13g2_fill_1 FILLER_34_1499 ();
 sg13g2_fill_2 FILLER_34_1545 ();
 sg13g2_fill_2 FILLER_34_1560 ();
 sg13g2_fill_1 FILLER_34_1606 ();
 sg13g2_fill_2 FILLER_34_1638 ();
 sg13g2_fill_2 FILLER_34_1667 ();
 sg13g2_fill_1 FILLER_34_1669 ();
 sg13g2_fill_1 FILLER_34_1695 ();
 sg13g2_fill_1 FILLER_34_1727 ();
 sg13g2_fill_1 FILLER_34_1767 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_54 ();
 sg13g2_fill_1 FILLER_35_56 ();
 sg13g2_fill_2 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_108 ();
 sg13g2_fill_2 FILLER_35_184 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_decap_4 FILLER_35_248 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_264 ();
 sg13g2_fill_2 FILLER_35_344 ();
 sg13g2_decap_4 FILLER_35_354 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_decap_4 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_35_424 ();
 sg13g2_fill_1 FILLER_35_438 ();
 sg13g2_decap_8 FILLER_35_445 ();
 sg13g2_decap_4 FILLER_35_452 ();
 sg13g2_fill_2 FILLER_35_461 ();
 sg13g2_decap_4 FILLER_35_468 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_fill_2 FILLER_35_483 ();
 sg13g2_fill_1 FILLER_35_485 ();
 sg13g2_decap_4 FILLER_35_494 ();
 sg13g2_fill_1 FILLER_35_498 ();
 sg13g2_fill_2 FILLER_35_502 ();
 sg13g2_fill_1 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_515 ();
 sg13g2_fill_1 FILLER_35_522 ();
 sg13g2_fill_2 FILLER_35_545 ();
 sg13g2_decap_8 FILLER_35_569 ();
 sg13g2_fill_2 FILLER_35_576 ();
 sg13g2_fill_1 FILLER_35_634 ();
 sg13g2_fill_2 FILLER_35_648 ();
 sg13g2_fill_1 FILLER_35_650 ();
 sg13g2_decap_8 FILLER_35_713 ();
 sg13g2_decap_8 FILLER_35_720 ();
 sg13g2_fill_2 FILLER_35_727 ();
 sg13g2_fill_2 FILLER_35_780 ();
 sg13g2_fill_2 FILLER_35_786 ();
 sg13g2_fill_1 FILLER_35_788 ();
 sg13g2_fill_2 FILLER_35_793 ();
 sg13g2_fill_2 FILLER_35_823 ();
 sg13g2_fill_2 FILLER_35_834 ();
 sg13g2_fill_2 FILLER_35_956 ();
 sg13g2_fill_1 FILLER_35_962 ();
 sg13g2_fill_2 FILLER_35_1024 ();
 sg13g2_fill_1 FILLER_35_1026 ();
 sg13g2_fill_2 FILLER_35_1069 ();
 sg13g2_fill_1 FILLER_35_1127 ();
 sg13g2_fill_1 FILLER_35_1137 ();
 sg13g2_fill_1 FILLER_35_1156 ();
 sg13g2_fill_1 FILLER_35_1170 ();
 sg13g2_fill_1 FILLER_35_1184 ();
 sg13g2_fill_2 FILLER_35_1226 ();
 sg13g2_fill_2 FILLER_35_1247 ();
 sg13g2_fill_1 FILLER_35_1267 ();
 sg13g2_fill_2 FILLER_35_1296 ();
 sg13g2_fill_1 FILLER_35_1330 ();
 sg13g2_decap_4 FILLER_35_1398 ();
 sg13g2_fill_2 FILLER_35_1406 ();
 sg13g2_fill_1 FILLER_35_1408 ();
 sg13g2_decap_8 FILLER_35_1417 ();
 sg13g2_decap_4 FILLER_35_1424 ();
 sg13g2_fill_1 FILLER_35_1457 ();
 sg13g2_fill_2 FILLER_35_1518 ();
 sg13g2_fill_1 FILLER_35_1546 ();
 sg13g2_fill_2 FILLER_35_1609 ();
 sg13g2_fill_2 FILLER_35_1689 ();
 sg13g2_fill_1 FILLER_35_1691 ();
 sg13g2_fill_2 FILLER_35_1710 ();
 sg13g2_fill_1 FILLER_35_1712 ();
 sg13g2_fill_2 FILLER_35_1734 ();
 sg13g2_fill_1 FILLER_35_1767 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_2 FILLER_36_90 ();
 sg13g2_fill_2 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_134 ();
 sg13g2_fill_1 FILLER_36_156 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_decap_4 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_268 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_decap_8 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_405 ();
 sg13g2_fill_2 FILLER_36_450 ();
 sg13g2_decap_4 FILLER_36_484 ();
 sg13g2_fill_1 FILLER_36_488 ();
 sg13g2_fill_1 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_509 ();
 sg13g2_fill_1 FILLER_36_548 ();
 sg13g2_fill_2 FILLER_36_576 ();
 sg13g2_decap_4 FILLER_36_587 ();
 sg13g2_fill_1 FILLER_36_591 ();
 sg13g2_decap_8 FILLER_36_620 ();
 sg13g2_fill_2 FILLER_36_627 ();
 sg13g2_fill_1 FILLER_36_629 ();
 sg13g2_decap_4 FILLER_36_723 ();
 sg13g2_fill_1 FILLER_36_727 ();
 sg13g2_decap_8 FILLER_36_736 ();
 sg13g2_decap_8 FILLER_36_751 ();
 sg13g2_fill_2 FILLER_36_758 ();
 sg13g2_fill_1 FILLER_36_760 ();
 sg13g2_fill_2 FILLER_36_771 ();
 sg13g2_decap_4 FILLER_36_779 ();
 sg13g2_decap_8 FILLER_36_787 ();
 sg13g2_fill_2 FILLER_36_794 ();
 sg13g2_fill_1 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_fill_2 FILLER_36_812 ();
 sg13g2_fill_1 FILLER_36_814 ();
 sg13g2_fill_1 FILLER_36_882 ();
 sg13g2_fill_2 FILLER_36_896 ();
 sg13g2_fill_1 FILLER_36_898 ();
 sg13g2_fill_1 FILLER_36_918 ();
 sg13g2_fill_1 FILLER_36_933 ();
 sg13g2_decap_4 FILLER_36_991 ();
 sg13g2_fill_1 FILLER_36_995 ();
 sg13g2_fill_1 FILLER_36_1050 ();
 sg13g2_fill_2 FILLER_36_1065 ();
 sg13g2_fill_1 FILLER_36_1117 ();
 sg13g2_fill_1 FILLER_36_1251 ();
 sg13g2_fill_1 FILLER_36_1266 ();
 sg13g2_fill_1 FILLER_36_1341 ();
 sg13g2_fill_1 FILLER_36_1403 ();
 sg13g2_fill_2 FILLER_36_1407 ();
 sg13g2_decap_4 FILLER_36_1418 ();
 sg13g2_fill_2 FILLER_36_1458 ();
 sg13g2_fill_2 FILLER_36_1497 ();
 sg13g2_fill_2 FILLER_36_1576 ();
 sg13g2_fill_2 FILLER_36_1621 ();
 sg13g2_fill_2 FILLER_36_1666 ();
 sg13g2_fill_1 FILLER_36_1681 ();
 sg13g2_fill_1 FILLER_36_1767 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_39 ();
 sg13g2_fill_1 FILLER_37_41 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_115 ();
 sg13g2_fill_1 FILLER_37_117 ();
 sg13g2_fill_1 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_249 ();
 sg13g2_fill_1 FILLER_37_251 ();
 sg13g2_decap_4 FILLER_37_256 ();
 sg13g2_fill_2 FILLER_37_336 ();
 sg13g2_decap_4 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_fill_1 FILLER_37_455 ();
 sg13g2_fill_2 FILLER_37_464 ();
 sg13g2_fill_2 FILLER_37_476 ();
 sg13g2_fill_1 FILLER_37_478 ();
 sg13g2_decap_4 FILLER_37_515 ();
 sg13g2_fill_1 FILLER_37_559 ();
 sg13g2_decap_8 FILLER_37_618 ();
 sg13g2_decap_4 FILLER_37_625 ();
 sg13g2_fill_1 FILLER_37_690 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_fill_2 FILLER_37_752 ();
 sg13g2_fill_2 FILLER_37_820 ();
 sg13g2_fill_1 FILLER_37_822 ();
 sg13g2_decap_4 FILLER_37_833 ();
 sg13g2_fill_1 FILLER_37_837 ();
 sg13g2_fill_2 FILLER_37_865 ();
 sg13g2_fill_2 FILLER_37_877 ();
 sg13g2_fill_1 FILLER_37_879 ();
 sg13g2_fill_2 FILLER_37_894 ();
 sg13g2_fill_2 FILLER_37_909 ();
 sg13g2_fill_1 FILLER_37_937 ();
 sg13g2_fill_2 FILLER_37_943 ();
 sg13g2_fill_1 FILLER_37_945 ();
 sg13g2_fill_1 FILLER_37_968 ();
 sg13g2_fill_1 FILLER_37_983 ();
 sg13g2_decap_4 FILLER_37_997 ();
 sg13g2_fill_1 FILLER_37_1005 ();
 sg13g2_fill_1 FILLER_37_1011 ();
 sg13g2_fill_1 FILLER_37_1025 ();
 sg13g2_fill_2 FILLER_37_1031 ();
 sg13g2_fill_2 FILLER_37_1163 ();
 sg13g2_fill_1 FILLER_37_1192 ();
 sg13g2_fill_1 FILLER_37_1207 ();
 sg13g2_fill_1 FILLER_37_1356 ();
 sg13g2_fill_2 FILLER_37_1383 ();
 sg13g2_fill_2 FILLER_37_1420 ();
 sg13g2_fill_2 FILLER_37_1508 ();
 sg13g2_decap_4 FILLER_37_1537 ();
 sg13g2_fill_1 FILLER_37_1541 ();
 sg13g2_fill_2 FILLER_37_1553 ();
 sg13g2_fill_1 FILLER_37_1571 ();
 sg13g2_fill_2 FILLER_37_1616 ();
 sg13g2_fill_2 FILLER_37_1640 ();
 sg13g2_fill_1 FILLER_37_1642 ();
 sg13g2_fill_2 FILLER_37_1675 ();
 sg13g2_fill_1 FILLER_37_1677 ();
 sg13g2_decap_4 FILLER_37_1722 ();
 sg13g2_fill_2 FILLER_37_1726 ();
 sg13g2_fill_1 FILLER_37_1749 ();
 sg13g2_decap_8 FILLER_37_1760 ();
 sg13g2_fill_1 FILLER_37_1767 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_2 FILLER_38_34 ();
 sg13g2_fill_1 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_158 ();
 sg13g2_fill_1 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_274 ();
 sg13g2_fill_1 FILLER_38_276 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_395 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_1 FILLER_38_432 ();
 sg13g2_decap_4 FILLER_38_447 ();
 sg13g2_fill_2 FILLER_38_462 ();
 sg13g2_fill_2 FILLER_38_478 ();
 sg13g2_fill_2 FILLER_38_513 ();
 sg13g2_fill_1 FILLER_38_515 ();
 sg13g2_fill_2 FILLER_38_529 ();
 sg13g2_fill_1 FILLER_38_538 ();
 sg13g2_fill_2 FILLER_38_567 ();
 sg13g2_fill_2 FILLER_38_573 ();
 sg13g2_fill_1 FILLER_38_575 ();
 sg13g2_fill_1 FILLER_38_604 ();
 sg13g2_fill_2 FILLER_38_627 ();
 sg13g2_fill_1 FILLER_38_657 ();
 sg13g2_fill_2 FILLER_38_671 ();
 sg13g2_fill_1 FILLER_38_708 ();
 sg13g2_fill_2 FILLER_38_769 ();
 sg13g2_decap_8 FILLER_38_783 ();
 sg13g2_decap_8 FILLER_38_794 ();
 sg13g2_decap_4 FILLER_38_801 ();
 sg13g2_fill_2 FILLER_38_805 ();
 sg13g2_fill_2 FILLER_38_834 ();
 sg13g2_decap_4 FILLER_38_846 ();
 sg13g2_fill_2 FILLER_38_881 ();
 sg13g2_fill_1 FILLER_38_910 ();
 sg13g2_fill_1 FILLER_38_916 ();
 sg13g2_fill_2 FILLER_38_983 ();
 sg13g2_decap_4 FILLER_38_994 ();
 sg13g2_fill_1 FILLER_38_1030 ();
 sg13g2_fill_1 FILLER_38_1045 ();
 sg13g2_fill_2 FILLER_38_1059 ();
 sg13g2_fill_1 FILLER_38_1061 ();
 sg13g2_fill_1 FILLER_38_1085 ();
 sg13g2_fill_2 FILLER_38_1104 ();
 sg13g2_fill_1 FILLER_38_1115 ();
 sg13g2_fill_1 FILLER_38_1143 ();
 sg13g2_decap_4 FILLER_38_1166 ();
 sg13g2_fill_2 FILLER_38_1178 ();
 sg13g2_fill_1 FILLER_38_1232 ();
 sg13g2_fill_2 FILLER_38_1255 ();
 sg13g2_fill_1 FILLER_38_1293 ();
 sg13g2_fill_1 FILLER_38_1352 ();
 sg13g2_fill_1 FILLER_38_1357 ();
 sg13g2_fill_2 FILLER_38_1390 ();
 sg13g2_fill_1 FILLER_38_1413 ();
 sg13g2_fill_1 FILLER_38_1420 ();
 sg13g2_fill_1 FILLER_38_1460 ();
 sg13g2_fill_1 FILLER_38_1479 ();
 sg13g2_fill_1 FILLER_38_1488 ();
 sg13g2_fill_2 FILLER_38_1506 ();
 sg13g2_fill_1 FILLER_38_1508 ();
 sg13g2_decap_4 FILLER_38_1632 ();
 sg13g2_fill_2 FILLER_38_1669 ();
 sg13g2_fill_2 FILLER_38_1725 ();
 sg13g2_fill_1 FILLER_38_1737 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_57 ();
 sg13g2_fill_1 FILLER_39_152 ();
 sg13g2_fill_1 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_fill_2 FILLER_39_295 ();
 sg13g2_fill_2 FILLER_39_326 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_fill_2 FILLER_39_382 ();
 sg13g2_fill_2 FILLER_39_397 ();
 sg13g2_fill_1 FILLER_39_399 ();
 sg13g2_fill_1 FILLER_39_410 ();
 sg13g2_fill_2 FILLER_39_465 ();
 sg13g2_fill_1 FILLER_39_467 ();
 sg13g2_fill_2 FILLER_39_500 ();
 sg13g2_fill_2 FILLER_39_529 ();
 sg13g2_fill_1 FILLER_39_531 ();
 sg13g2_fill_1 FILLER_39_537 ();
 sg13g2_fill_1 FILLER_39_569 ();
 sg13g2_fill_1 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_639 ();
 sg13g2_decap_4 FILLER_39_651 ();
 sg13g2_fill_2 FILLER_39_664 ();
 sg13g2_fill_1 FILLER_39_666 ();
 sg13g2_fill_1 FILLER_39_676 ();
 sg13g2_fill_1 FILLER_39_700 ();
 sg13g2_fill_2 FILLER_39_720 ();
 sg13g2_fill_1 FILLER_39_722 ();
 sg13g2_fill_1 FILLER_39_745 ();
 sg13g2_fill_1 FILLER_39_755 ();
 sg13g2_decap_4 FILLER_39_766 ();
 sg13g2_fill_1 FILLER_39_770 ();
 sg13g2_fill_2 FILLER_39_782 ();
 sg13g2_fill_1 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_817 ();
 sg13g2_fill_2 FILLER_39_824 ();
 sg13g2_fill_1 FILLER_39_921 ();
 sg13g2_fill_2 FILLER_39_940 ();
 sg13g2_fill_2 FILLER_39_978 ();
 sg13g2_fill_1 FILLER_39_1316 ();
 sg13g2_fill_2 FILLER_39_1362 ();
 sg13g2_fill_1 FILLER_39_1393 ();
 sg13g2_fill_1 FILLER_39_1434 ();
 sg13g2_fill_2 FILLER_39_1443 ();
 sg13g2_fill_1 FILLER_39_1448 ();
 sg13g2_fill_2 FILLER_39_1484 ();
 sg13g2_fill_1 FILLER_39_1486 ();
 sg13g2_fill_1 FILLER_39_1508 ();
 sg13g2_fill_1 FILLER_39_1522 ();
 sg13g2_fill_1 FILLER_39_1614 ();
 sg13g2_fill_2 FILLER_39_1627 ();
 sg13g2_fill_2 FILLER_39_1660 ();
 sg13g2_fill_2 FILLER_39_1666 ();
 sg13g2_fill_2 FILLER_39_1698 ();
 sg13g2_fill_1 FILLER_39_1745 ();
 sg13g2_fill_1 FILLER_39_1754 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_28 ();
 sg13g2_fill_1 FILLER_40_86 ();
 sg13g2_fill_2 FILLER_40_105 ();
 sg13g2_fill_2 FILLER_40_116 ();
 sg13g2_fill_1 FILLER_40_118 ();
 sg13g2_fill_2 FILLER_40_281 ();
 sg13g2_fill_1 FILLER_40_283 ();
 sg13g2_fill_1 FILLER_40_318 ();
 sg13g2_fill_2 FILLER_40_329 ();
 sg13g2_fill_2 FILLER_40_350 ();
 sg13g2_fill_1 FILLER_40_376 ();
 sg13g2_fill_2 FILLER_40_387 ();
 sg13g2_fill_1 FILLER_40_389 ();
 sg13g2_fill_2 FILLER_40_442 ();
 sg13g2_fill_1 FILLER_40_457 ();
 sg13g2_fill_2 FILLER_40_471 ();
 sg13g2_fill_2 FILLER_40_491 ();
 sg13g2_decap_4 FILLER_40_497 ();
 sg13g2_fill_1 FILLER_40_501 ();
 sg13g2_fill_1 FILLER_40_506 ();
 sg13g2_decap_4 FILLER_40_511 ();
 sg13g2_fill_2 FILLER_40_515 ();
 sg13g2_fill_2 FILLER_40_526 ();
 sg13g2_decap_4 FILLER_40_548 ();
 sg13g2_fill_2 FILLER_40_552 ();
 sg13g2_fill_2 FILLER_40_596 ();
 sg13g2_fill_1 FILLER_40_598 ();
 sg13g2_fill_1 FILLER_40_619 ();
 sg13g2_fill_2 FILLER_40_639 ();
 sg13g2_fill_1 FILLER_40_641 ();
 sg13g2_fill_1 FILLER_40_656 ();
 sg13g2_fill_2 FILLER_40_736 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_fill_2 FILLER_40_843 ();
 sg13g2_fill_2 FILLER_40_876 ();
 sg13g2_fill_1 FILLER_40_878 ();
 sg13g2_fill_2 FILLER_40_946 ();
 sg13g2_fill_1 FILLER_40_948 ();
 sg13g2_fill_1 FILLER_40_1011 ();
 sg13g2_fill_1 FILLER_40_1029 ();
 sg13g2_fill_2 FILLER_40_1056 ();
 sg13g2_fill_2 FILLER_40_1105 ();
 sg13g2_decap_4 FILLER_40_1172 ();
 sg13g2_fill_1 FILLER_40_1176 ();
 sg13g2_fill_1 FILLER_40_1205 ();
 sg13g2_fill_2 FILLER_40_1234 ();
 sg13g2_fill_1 FILLER_40_1242 ();
 sg13g2_fill_2 FILLER_40_1260 ();
 sg13g2_fill_1 FILLER_40_1262 ();
 sg13g2_fill_2 FILLER_40_1281 ();
 sg13g2_fill_2 FILLER_40_1310 ();
 sg13g2_fill_2 FILLER_40_1315 ();
 sg13g2_fill_1 FILLER_40_1471 ();
 sg13g2_decap_4 FILLER_40_1485 ();
 sg13g2_fill_1 FILLER_40_1489 ();
 sg13g2_fill_2 FILLER_40_1512 ();
 sg13g2_fill_1 FILLER_40_1514 ();
 sg13g2_fill_1 FILLER_40_1542 ();
 sg13g2_decap_8 FILLER_40_1600 ();
 sg13g2_fill_1 FILLER_40_1627 ();
 sg13g2_fill_1 FILLER_40_1651 ();
 sg13g2_fill_2 FILLER_40_1684 ();
 sg13g2_fill_2 FILLER_40_1726 ();
 sg13g2_fill_1 FILLER_40_1767 ();
 sg13g2_fill_2 FILLER_41_0 ();
 sg13g2_fill_2 FILLER_41_52 ();
 sg13g2_fill_1 FILLER_41_94 ();
 sg13g2_fill_1 FILLER_41_163 ();
 sg13g2_fill_2 FILLER_41_191 ();
 sg13g2_fill_1 FILLER_41_215 ();
 sg13g2_fill_2 FILLER_41_249 ();
 sg13g2_fill_2 FILLER_41_306 ();
 sg13g2_fill_2 FILLER_41_318 ();
 sg13g2_fill_2 FILLER_41_324 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_fill_1 FILLER_41_340 ();
 sg13g2_fill_1 FILLER_41_377 ();
 sg13g2_fill_2 FILLER_41_405 ();
 sg13g2_fill_1 FILLER_41_422 ();
 sg13g2_fill_1 FILLER_41_441 ();
 sg13g2_fill_1 FILLER_41_447 ();
 sg13g2_fill_2 FILLER_41_465 ();
 sg13g2_fill_1 FILLER_41_481 ();
 sg13g2_fill_2 FILLER_41_525 ();
 sg13g2_fill_1 FILLER_41_527 ();
 sg13g2_fill_2 FILLER_41_565 ();
 sg13g2_fill_1 FILLER_41_576 ();
 sg13g2_fill_2 FILLER_41_586 ();
 sg13g2_fill_1 FILLER_41_588 ();
 sg13g2_fill_2 FILLER_41_616 ();
 sg13g2_fill_1 FILLER_41_618 ();
 sg13g2_decap_4 FILLER_41_652 ();
 sg13g2_fill_1 FILLER_41_656 ();
 sg13g2_fill_1 FILLER_41_670 ();
 sg13g2_fill_2 FILLER_41_680 ();
 sg13g2_fill_1 FILLER_41_682 ();
 sg13g2_fill_1 FILLER_41_712 ();
 sg13g2_fill_2 FILLER_41_722 ();
 sg13g2_decap_4 FILLER_41_737 ();
 sg13g2_fill_2 FILLER_41_741 ();
 sg13g2_fill_2 FILLER_41_758 ();
 sg13g2_fill_1 FILLER_41_760 ();
 sg13g2_fill_2 FILLER_41_765 ();
 sg13g2_fill_2 FILLER_41_775 ();
 sg13g2_fill_1 FILLER_41_777 ();
 sg13g2_decap_4 FILLER_41_841 ();
 sg13g2_fill_2 FILLER_41_845 ();
 sg13g2_fill_1 FILLER_41_875 ();
 sg13g2_fill_2 FILLER_41_907 ();
 sg13g2_fill_2 FILLER_41_923 ();
 sg13g2_fill_2 FILLER_41_962 ();
 sg13g2_fill_1 FILLER_41_1020 ();
 sg13g2_fill_1 FILLER_41_1055 ();
 sg13g2_fill_1 FILLER_41_1091 ();
 sg13g2_fill_2 FILLER_41_1142 ();
 sg13g2_fill_2 FILLER_41_1158 ();
 sg13g2_fill_1 FILLER_41_1160 ();
 sg13g2_fill_2 FILLER_41_1189 ();
 sg13g2_fill_2 FILLER_41_1200 ();
 sg13g2_fill_1 FILLER_41_1202 ();
 sg13g2_fill_2 FILLER_41_1209 ();
 sg13g2_fill_1 FILLER_41_1211 ();
 sg13g2_fill_2 FILLER_41_1220 ();
 sg13g2_fill_1 FILLER_41_1315 ();
 sg13g2_fill_2 FILLER_41_1337 ();
 sg13g2_fill_1 FILLER_41_1339 ();
 sg13g2_fill_1 FILLER_41_1349 ();
 sg13g2_fill_1 FILLER_41_1367 ();
 sg13g2_fill_2 FILLER_41_1390 ();
 sg13g2_fill_2 FILLER_41_1404 ();
 sg13g2_fill_1 FILLER_41_1416 ();
 sg13g2_fill_2 FILLER_41_1444 ();
 sg13g2_fill_1 FILLER_41_1446 ();
 sg13g2_fill_1 FILLER_41_1456 ();
 sg13g2_fill_2 FILLER_41_1505 ();
 sg13g2_fill_1 FILLER_41_1525 ();
 sg13g2_fill_2 FILLER_41_1547 ();
 sg13g2_fill_1 FILLER_41_1566 ();
 sg13g2_fill_2 FILLER_41_1576 ();
 sg13g2_fill_1 FILLER_41_1589 ();
 sg13g2_fill_1 FILLER_41_1594 ();
 sg13g2_fill_1 FILLER_41_1640 ();
 sg13g2_fill_2 FILLER_41_1657 ();
 sg13g2_fill_2 FILLER_41_1665 ();
 sg13g2_fill_2 FILLER_41_1676 ();
 sg13g2_fill_1 FILLER_41_1712 ();
 sg13g2_fill_1 FILLER_41_1729 ();
 sg13g2_fill_1 FILLER_41_1734 ();
 sg13g2_fill_2 FILLER_41_1739 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_32 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_fill_2 FILLER_42_45 ();
 sg13g2_fill_1 FILLER_42_61 ();
 sg13g2_fill_2 FILLER_42_71 ();
 sg13g2_fill_1 FILLER_42_120 ();
 sg13g2_fill_1 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_209 ();
 sg13g2_fill_2 FILLER_42_242 ();
 sg13g2_fill_2 FILLER_42_253 ();
 sg13g2_fill_1 FILLER_42_255 ();
 sg13g2_fill_1 FILLER_42_308 ();
 sg13g2_fill_1 FILLER_42_314 ();
 sg13g2_fill_1 FILLER_42_369 ();
 sg13g2_fill_2 FILLER_42_395 ();
 sg13g2_fill_1 FILLER_42_451 ();
 sg13g2_fill_2 FILLER_42_484 ();
 sg13g2_fill_1 FILLER_42_486 ();
 sg13g2_fill_2 FILLER_42_500 ();
 sg13g2_fill_2 FILLER_42_515 ();
 sg13g2_fill_1 FILLER_42_536 ();
 sg13g2_fill_2 FILLER_42_550 ();
 sg13g2_fill_1 FILLER_42_552 ();
 sg13g2_fill_2 FILLER_42_599 ();
 sg13g2_fill_1 FILLER_42_624 ();
 sg13g2_fill_1 FILLER_42_650 ();
 sg13g2_fill_2 FILLER_42_693 ();
 sg13g2_fill_1 FILLER_42_724 ();
 sg13g2_fill_2 FILLER_42_730 ();
 sg13g2_decap_4 FILLER_42_759 ();
 sg13g2_fill_1 FILLER_42_763 ();
 sg13g2_fill_2 FILLER_42_790 ();
 sg13g2_decap_4 FILLER_42_819 ();
 sg13g2_decap_4 FILLER_42_849 ();
 sg13g2_fill_1 FILLER_42_853 ();
 sg13g2_fill_1 FILLER_42_918 ();
 sg13g2_fill_2 FILLER_42_958 ();
 sg13g2_fill_1 FILLER_42_960 ();
 sg13g2_fill_2 FILLER_42_993 ();
 sg13g2_fill_1 FILLER_42_995 ();
 sg13g2_fill_1 FILLER_42_1054 ();
 sg13g2_fill_2 FILLER_42_1082 ();
 sg13g2_fill_2 FILLER_42_1100 ();
 sg13g2_decap_4 FILLER_42_1179 ();
 sg13g2_fill_2 FILLER_42_1183 ();
 sg13g2_fill_1 FILLER_42_1197 ();
 sg13g2_fill_2 FILLER_42_1241 ();
 sg13g2_fill_1 FILLER_42_1243 ();
 sg13g2_fill_1 FILLER_42_1248 ();
 sg13g2_decap_8 FILLER_42_1313 ();
 sg13g2_decap_8 FILLER_42_1320 ();
 sg13g2_fill_2 FILLER_42_1327 ();
 sg13g2_fill_1 FILLER_42_1329 ();
 sg13g2_fill_2 FILLER_42_1396 ();
 sg13g2_fill_2 FILLER_42_1429 ();
 sg13g2_fill_1 FILLER_42_1431 ();
 sg13g2_fill_1 FILLER_42_1497 ();
 sg13g2_fill_2 FILLER_42_1524 ();
 sg13g2_fill_1 FILLER_42_1593 ();
 sg13g2_fill_2 FILLER_42_1607 ();
 sg13g2_fill_2 FILLER_42_1625 ();
 sg13g2_decap_8 FILLER_42_1630 ();
 sg13g2_fill_2 FILLER_42_1717 ();
 sg13g2_fill_2 FILLER_42_1751 ();
 sg13g2_fill_2 FILLER_42_1766 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_2 ();
 sg13g2_fill_1 FILLER_43_83 ();
 sg13g2_fill_2 FILLER_43_93 ();
 sg13g2_fill_1 FILLER_43_122 ();
 sg13g2_fill_1 FILLER_43_148 ();
 sg13g2_fill_2 FILLER_43_162 ();
 sg13g2_fill_1 FILLER_43_164 ();
 sg13g2_fill_2 FILLER_43_178 ();
 sg13g2_fill_1 FILLER_43_180 ();
 sg13g2_fill_2 FILLER_43_190 ();
 sg13g2_fill_2 FILLER_43_202 ();
 sg13g2_fill_2 FILLER_43_226 ();
 sg13g2_fill_1 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_251 ();
 sg13g2_fill_1 FILLER_43_318 ();
 sg13g2_fill_2 FILLER_43_371 ();
 sg13g2_fill_2 FILLER_43_413 ();
 sg13g2_fill_1 FILLER_43_415 ();
 sg13g2_fill_2 FILLER_43_425 ();
 sg13g2_fill_2 FILLER_43_464 ();
 sg13g2_fill_2 FILLER_43_573 ();
 sg13g2_fill_2 FILLER_43_594 ();
 sg13g2_fill_1 FILLER_43_596 ();
 sg13g2_decap_4 FILLER_43_660 ();
 sg13g2_fill_2 FILLER_43_664 ();
 sg13g2_decap_8 FILLER_43_670 ();
 sg13g2_fill_2 FILLER_43_724 ();
 sg13g2_decap_4 FILLER_43_734 ();
 sg13g2_fill_1 FILLER_43_738 ();
 sg13g2_decap_4 FILLER_43_751 ();
 sg13g2_fill_2 FILLER_43_755 ();
 sg13g2_fill_2 FILLER_43_801 ();
 sg13g2_fill_1 FILLER_43_803 ();
 sg13g2_fill_2 FILLER_43_814 ();
 sg13g2_fill_1 FILLER_43_816 ();
 sg13g2_fill_2 FILLER_43_825 ();
 sg13g2_fill_1 FILLER_43_827 ();
 sg13g2_decap_8 FILLER_43_838 ();
 sg13g2_fill_1 FILLER_43_845 ();
 sg13g2_fill_2 FILLER_43_882 ();
 sg13g2_fill_1 FILLER_43_894 ();
 sg13g2_fill_2 FILLER_43_953 ();
 sg13g2_fill_1 FILLER_43_989 ();
 sg13g2_fill_2 FILLER_43_1035 ();
 sg13g2_fill_1 FILLER_43_1037 ();
 sg13g2_fill_2 FILLER_43_1047 ();
 sg13g2_fill_2 FILLER_43_1085 ();
 sg13g2_fill_1 FILLER_43_1121 ();
 sg13g2_fill_2 FILLER_43_1141 ();
 sg13g2_decap_8 FILLER_43_1175 ();
 sg13g2_decap_4 FILLER_43_1182 ();
 sg13g2_fill_2 FILLER_43_1186 ();
 sg13g2_fill_1 FILLER_43_1196 ();
 sg13g2_fill_2 FILLER_43_1220 ();
 sg13g2_fill_1 FILLER_43_1222 ();
 sg13g2_fill_2 FILLER_43_1245 ();
 sg13g2_fill_1 FILLER_43_1247 ();
 sg13g2_fill_2 FILLER_43_1291 ();
 sg13g2_decap_8 FILLER_43_1305 ();
 sg13g2_fill_2 FILLER_43_1312 ();
 sg13g2_fill_1 FILLER_43_1314 ();
 sg13g2_fill_2 FILLER_43_1357 ();
 sg13g2_fill_1 FILLER_43_1386 ();
 sg13g2_decap_4 FILLER_43_1399 ();
 sg13g2_fill_2 FILLER_43_1403 ();
 sg13g2_fill_2 FILLER_43_1410 ();
 sg13g2_fill_1 FILLER_43_1424 ();
 sg13g2_fill_2 FILLER_43_1428 ();
 sg13g2_fill_1 FILLER_43_1443 ();
 sg13g2_fill_1 FILLER_43_1451 ();
 sg13g2_fill_1 FILLER_43_1474 ();
 sg13g2_fill_2 FILLER_43_1481 ();
 sg13g2_fill_1 FILLER_43_1496 ();
 sg13g2_decap_4 FILLER_43_1617 ();
 sg13g2_fill_2 FILLER_43_1621 ();
 sg13g2_fill_2 FILLER_43_1632 ();
 sg13g2_fill_2 FILLER_43_1637 ();
 sg13g2_fill_1 FILLER_43_1639 ();
 sg13g2_fill_2 FILLER_43_1694 ();
 sg13g2_fill_2 FILLER_43_1705 ();
 sg13g2_fill_1 FILLER_43_1711 ();
 sg13g2_fill_2 FILLER_43_1750 ();
 sg13g2_fill_1 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_33 ();
 sg13g2_fill_1 FILLER_44_35 ();
 sg13g2_fill_1 FILLER_44_63 ();
 sg13g2_fill_2 FILLER_44_141 ();
 sg13g2_fill_1 FILLER_44_180 ();
 sg13g2_fill_2 FILLER_44_258 ();
 sg13g2_fill_2 FILLER_44_341 ();
 sg13g2_fill_2 FILLER_44_352 ();
 sg13g2_fill_1 FILLER_44_427 ();
 sg13g2_fill_2 FILLER_44_464 ();
 sg13g2_fill_1 FILLER_44_466 ();
 sg13g2_fill_2 FILLER_44_570 ();
 sg13g2_fill_1 FILLER_44_588 ();
 sg13g2_fill_2 FILLER_44_617 ();
 sg13g2_fill_2 FILLER_44_629 ();
 sg13g2_fill_2 FILLER_44_695 ();
 sg13g2_fill_1 FILLER_44_706 ();
 sg13g2_fill_2 FILLER_44_722 ();
 sg13g2_fill_2 FILLER_44_729 ();
 sg13g2_decap_4 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_743 ();
 sg13g2_decap_8 FILLER_44_750 ();
 sg13g2_fill_2 FILLER_44_757 ();
 sg13g2_fill_1 FILLER_44_799 ();
 sg13g2_fill_2 FILLER_44_809 ();
 sg13g2_decap_4 FILLER_44_816 ();
 sg13g2_fill_2 FILLER_44_831 ();
 sg13g2_fill_1 FILLER_44_833 ();
 sg13g2_fill_1 FILLER_44_847 ();
 sg13g2_fill_1 FILLER_44_882 ();
 sg13g2_decap_4 FILLER_44_896 ();
 sg13g2_fill_1 FILLER_44_900 ();
 sg13g2_fill_2 FILLER_44_967 ();
 sg13g2_fill_2 FILLER_44_982 ();
 sg13g2_fill_2 FILLER_44_1018 ();
 sg13g2_fill_1 FILLER_44_1066 ();
 sg13g2_fill_1 FILLER_44_1111 ();
 sg13g2_fill_1 FILLER_44_1185 ();
 sg13g2_fill_2 FILLER_44_1190 ();
 sg13g2_fill_1 FILLER_44_1192 ();
 sg13g2_fill_1 FILLER_44_1233 ();
 sg13g2_fill_1 FILLER_44_1247 ();
 sg13g2_fill_1 FILLER_44_1302 ();
 sg13g2_fill_1 FILLER_44_1307 ();
 sg13g2_fill_2 FILLER_44_1343 ();
 sg13g2_fill_1 FILLER_44_1438 ();
 sg13g2_decap_4 FILLER_44_1448 ();
 sg13g2_fill_2 FILLER_44_1452 ();
 sg13g2_decap_8 FILLER_44_1496 ();
 sg13g2_fill_2 FILLER_44_1503 ();
 sg13g2_fill_2 FILLER_44_1647 ();
 sg13g2_fill_2 FILLER_44_1734 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_1 FILLER_45_2 ();
 sg13g2_fill_2 FILLER_45_30 ();
 sg13g2_fill_1 FILLER_45_32 ();
 sg13g2_fill_1 FILLER_45_82 ();
 sg13g2_fill_1 FILLER_45_138 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_185 ();
 sg13g2_fill_2 FILLER_45_253 ();
 sg13g2_fill_2 FILLER_45_286 ();
 sg13g2_fill_2 FILLER_45_348 ();
 sg13g2_fill_2 FILLER_45_377 ();
 sg13g2_fill_1 FILLER_45_490 ();
 sg13g2_fill_1 FILLER_45_504 ();
 sg13g2_fill_2 FILLER_45_553 ();
 sg13g2_fill_1 FILLER_45_581 ();
 sg13g2_fill_2 FILLER_45_664 ();
 sg13g2_fill_1 FILLER_45_666 ();
 sg13g2_fill_2 FILLER_45_721 ();
 sg13g2_decap_4 FILLER_45_770 ();
 sg13g2_fill_1 FILLER_45_774 ();
 sg13g2_fill_1 FILLER_45_816 ();
 sg13g2_fill_2 FILLER_45_832 ();
 sg13g2_fill_1 FILLER_45_889 ();
 sg13g2_fill_2 FILLER_45_922 ();
 sg13g2_fill_1 FILLER_45_924 ();
 sg13g2_fill_2 FILLER_45_935 ();
 sg13g2_fill_2 FILLER_45_951 ();
 sg13g2_fill_1 FILLER_45_953 ();
 sg13g2_decap_8 FILLER_45_1002 ();
 sg13g2_fill_2 FILLER_45_1009 ();
 sg13g2_decap_4 FILLER_45_1018 ();
 sg13g2_fill_2 FILLER_45_1022 ();
 sg13g2_fill_1 FILLER_45_1056 ();
 sg13g2_fill_1 FILLER_45_1107 ();
 sg13g2_fill_2 FILLER_45_1150 ();
 sg13g2_fill_1 FILLER_45_1152 ();
 sg13g2_fill_1 FILLER_45_1194 ();
 sg13g2_decap_4 FILLER_45_1203 ();
 sg13g2_decap_4 FILLER_45_1216 ();
 sg13g2_fill_2 FILLER_45_1296 ();
 sg13g2_decap_8 FILLER_45_1358 ();
 sg13g2_decap_8 FILLER_45_1365 ();
 sg13g2_decap_8 FILLER_45_1372 ();
 sg13g2_decap_8 FILLER_45_1379 ();
 sg13g2_fill_2 FILLER_45_1386 ();
 sg13g2_decap_4 FILLER_45_1396 ();
 sg13g2_fill_2 FILLER_45_1400 ();
 sg13g2_decap_4 FILLER_45_1411 ();
 sg13g2_fill_2 FILLER_45_1432 ();
 sg13g2_fill_1 FILLER_45_1434 ();
 sg13g2_fill_2 FILLER_45_1468 ();
 sg13g2_decap_8 FILLER_45_1496 ();
 sg13g2_fill_1 FILLER_45_1503 ();
 sg13g2_fill_2 FILLER_45_1579 ();
 sg13g2_fill_2 FILLER_45_1598 ();
 sg13g2_fill_1 FILLER_45_1670 ();
 sg13g2_fill_2 FILLER_45_1680 ();
 sg13g2_fill_2 FILLER_45_1730 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_37 ();
 sg13g2_fill_1 FILLER_46_68 ();
 sg13g2_fill_1 FILLER_46_92 ();
 sg13g2_fill_1 FILLER_46_169 ();
 sg13g2_fill_1 FILLER_46_183 ();
 sg13g2_fill_2 FILLER_46_242 ();
 sg13g2_fill_2 FILLER_46_256 ();
 sg13g2_fill_2 FILLER_46_343 ();
 sg13g2_fill_1 FILLER_46_345 ();
 sg13g2_fill_1 FILLER_46_416 ();
 sg13g2_fill_1 FILLER_46_446 ();
 sg13g2_fill_2 FILLER_46_489 ();
 sg13g2_fill_2 FILLER_46_539 ();
 sg13g2_fill_1 FILLER_46_550 ();
 sg13g2_fill_2 FILLER_46_588 ();
 sg13g2_fill_2 FILLER_46_630 ();
 sg13g2_fill_2 FILLER_46_671 ();
 sg13g2_fill_1 FILLER_46_673 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_fill_2 FILLER_46_738 ();
 sg13g2_fill_1 FILLER_46_740 ();
 sg13g2_fill_2 FILLER_46_769 ();
 sg13g2_fill_1 FILLER_46_771 ();
 sg13g2_decap_8 FILLER_46_776 ();
 sg13g2_decap_4 FILLER_46_783 ();
 sg13g2_fill_2 FILLER_46_787 ();
 sg13g2_fill_1 FILLER_46_793 ();
 sg13g2_fill_2 FILLER_46_803 ();
 sg13g2_fill_1 FILLER_46_805 ();
 sg13g2_decap_4 FILLER_46_825 ();
 sg13g2_fill_1 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_846 ();
 sg13g2_fill_2 FILLER_46_853 ();
 sg13g2_fill_2 FILLER_46_867 ();
 sg13g2_fill_1 FILLER_46_869 ();
 sg13g2_decap_4 FILLER_46_879 ();
 sg13g2_fill_2 FILLER_46_896 ();
 sg13g2_fill_1 FILLER_46_920 ();
 sg13g2_fill_2 FILLER_46_930 ();
 sg13g2_fill_1 FILLER_46_959 ();
 sg13g2_fill_1 FILLER_46_992 ();
 sg13g2_fill_1 FILLER_46_1003 ();
 sg13g2_fill_1 FILLER_46_1098 ();
 sg13g2_fill_2 FILLER_46_1137 ();
 sg13g2_fill_2 FILLER_46_1157 ();
 sg13g2_fill_2 FILLER_46_1199 ();
 sg13g2_fill_1 FILLER_46_1283 ();
 sg13g2_decap_4 FILLER_46_1371 ();
 sg13g2_fill_2 FILLER_46_1375 ();
 sg13g2_fill_1 FILLER_46_1431 ();
 sg13g2_decap_4 FILLER_46_1461 ();
 sg13g2_fill_2 FILLER_46_1537 ();
 sg13g2_fill_2 FILLER_46_1566 ();
 sg13g2_fill_1 FILLER_46_1640 ();
 sg13g2_fill_2 FILLER_46_1702 ();
 sg13g2_fill_1 FILLER_46_1713 ();
 sg13g2_fill_1 FILLER_46_1740 ();
 sg13g2_fill_2 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_2 ();
 sg13g2_fill_2 FILLER_47_38 ();
 sg13g2_fill_1 FILLER_47_40 ();
 sg13g2_fill_2 FILLER_47_132 ();
 sg13g2_fill_2 FILLER_47_266 ();
 sg13g2_fill_1 FILLER_47_268 ();
 sg13g2_fill_2 FILLER_47_379 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_47_459 ();
 sg13g2_fill_1 FILLER_47_524 ();
 sg13g2_fill_1 FILLER_47_535 ();
 sg13g2_fill_1 FILLER_47_550 ();
 sg13g2_fill_2 FILLER_47_556 ();
 sg13g2_fill_1 FILLER_47_558 ();
 sg13g2_fill_2 FILLER_47_564 ();
 sg13g2_fill_1 FILLER_47_566 ();
 sg13g2_fill_1 FILLER_47_600 ();
 sg13g2_fill_2 FILLER_47_637 ();
 sg13g2_fill_2 FILLER_47_657 ();
 sg13g2_fill_2 FILLER_47_671 ();
 sg13g2_fill_2 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_679 ();
 sg13g2_fill_1 FILLER_47_717 ();
 sg13g2_decap_4 FILLER_47_722 ();
 sg13g2_decap_8 FILLER_47_732 ();
 sg13g2_fill_1 FILLER_47_739 ();
 sg13g2_decap_8 FILLER_47_754 ();
 sg13g2_fill_2 FILLER_47_761 ();
 sg13g2_decap_4 FILLER_47_809 ();
 sg13g2_fill_1 FILLER_47_819 ();
 sg13g2_fill_2 FILLER_47_868 ();
 sg13g2_fill_1 FILLER_47_870 ();
 sg13g2_fill_1 FILLER_47_879 ();
 sg13g2_fill_2 FILLER_47_911 ();
 sg13g2_fill_1 FILLER_47_940 ();
 sg13g2_fill_1 FILLER_47_959 ();
 sg13g2_fill_2 FILLER_47_988 ();
 sg13g2_fill_1 FILLER_47_990 ();
 sg13g2_fill_2 FILLER_47_1008 ();
 sg13g2_fill_1 FILLER_47_1022 ();
 sg13g2_fill_2 FILLER_47_1068 ();
 sg13g2_fill_1 FILLER_47_1070 ();
 sg13g2_fill_2 FILLER_47_1084 ();
 sg13g2_fill_1 FILLER_47_1086 ();
 sg13g2_fill_2 FILLER_47_1093 ();
 sg13g2_fill_1 FILLER_47_1127 ();
 sg13g2_fill_2 FILLER_47_1207 ();
 sg13g2_fill_1 FILLER_47_1209 ();
 sg13g2_decap_8 FILLER_47_1219 ();
 sg13g2_decap_4 FILLER_47_1226 ();
 sg13g2_fill_2 FILLER_47_1230 ();
 sg13g2_decap_4 FILLER_47_1240 ();
 sg13g2_fill_1 FILLER_47_1251 ();
 sg13g2_fill_2 FILLER_47_1265 ();
 sg13g2_fill_1 FILLER_47_1318 ();
 sg13g2_fill_1 FILLER_47_1341 ();
 sg13g2_fill_2 FILLER_47_1351 ();
 sg13g2_fill_1 FILLER_47_1353 ();
 sg13g2_fill_2 FILLER_47_1381 ();
 sg13g2_fill_2 FILLER_47_1397 ();
 sg13g2_fill_1 FILLER_47_1399 ();
 sg13g2_fill_1 FILLER_47_1409 ();
 sg13g2_fill_1 FILLER_47_1422 ();
 sg13g2_fill_2 FILLER_47_1437 ();
 sg13g2_fill_1 FILLER_47_1439 ();
 sg13g2_fill_2 FILLER_47_1478 ();
 sg13g2_fill_2 FILLER_47_1484 ();
 sg13g2_fill_1 FILLER_47_1498 ();
 sg13g2_fill_1 FILLER_47_1559 ();
 sg13g2_fill_2 FILLER_47_1591 ();
 sg13g2_decap_4 FILLER_47_1636 ();
 sg13g2_fill_1 FILLER_47_1672 ();
 sg13g2_fill_2 FILLER_47_1711 ();
 sg13g2_fill_2 FILLER_47_1745 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_2 FILLER_48_45 ();
 sg13g2_fill_1 FILLER_48_47 ();
 sg13g2_fill_2 FILLER_48_58 ();
 sg13g2_fill_2 FILLER_48_88 ();
 sg13g2_fill_2 FILLER_48_120 ();
 sg13g2_fill_2 FILLER_48_173 ();
 sg13g2_fill_1 FILLER_48_175 ();
 sg13g2_fill_1 FILLER_48_186 ();
 sg13g2_fill_1 FILLER_48_318 ();
 sg13g2_fill_2 FILLER_48_378 ();
 sg13g2_fill_2 FILLER_48_393 ();
 sg13g2_fill_2 FILLER_48_431 ();
 sg13g2_fill_2 FILLER_48_485 ();
 sg13g2_fill_1 FILLER_48_487 ();
 sg13g2_fill_2 FILLER_48_498 ();
 sg13g2_fill_1 FILLER_48_527 ();
 sg13g2_fill_1 FILLER_48_547 ();
 sg13g2_fill_2 FILLER_48_710 ();
 sg13g2_fill_2 FILLER_48_740 ();
 sg13g2_fill_1 FILLER_48_742 ();
 sg13g2_decap_4 FILLER_48_755 ();
 sg13g2_fill_1 FILLER_48_775 ();
 sg13g2_decap_4 FILLER_48_780 ();
 sg13g2_fill_2 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_4 FILLER_48_826 ();
 sg13g2_fill_1 FILLER_48_830 ();
 sg13g2_fill_1 FILLER_48_885 ();
 sg13g2_fill_1 FILLER_48_912 ();
 sg13g2_fill_1 FILLER_48_977 ();
 sg13g2_fill_2 FILLER_48_1012 ();
 sg13g2_fill_1 FILLER_48_1014 ();
 sg13g2_fill_2 FILLER_48_1043 ();
 sg13g2_fill_2 FILLER_48_1098 ();
 sg13g2_fill_2 FILLER_48_1130 ();
 sg13g2_fill_2 FILLER_48_1155 ();
 sg13g2_fill_1 FILLER_48_1189 ();
 sg13g2_decap_8 FILLER_48_1198 ();
 sg13g2_decap_4 FILLER_48_1205 ();
 sg13g2_fill_2 FILLER_48_1209 ();
 sg13g2_fill_1 FILLER_48_1216 ();
 sg13g2_decap_8 FILLER_48_1221 ();
 sg13g2_decap_8 FILLER_48_1228 ();
 sg13g2_fill_1 FILLER_48_1263 ();
 sg13g2_decap_4 FILLER_48_1395 ();
 sg13g2_fill_2 FILLER_48_1404 ();
 sg13g2_fill_1 FILLER_48_1406 ();
 sg13g2_fill_2 FILLER_48_1455 ();
 sg13g2_fill_1 FILLER_48_1466 ();
 sg13g2_fill_1 FILLER_48_1504 ();
 sg13g2_fill_2 FILLER_48_1562 ();
 sg13g2_fill_2 FILLER_48_1656 ();
 sg13g2_fill_2 FILLER_48_1685 ();
 sg13g2_fill_2 FILLER_48_1698 ();
 sg13g2_fill_1 FILLER_48_1767 ();
 sg13g2_fill_2 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_57 ();
 sg13g2_fill_2 FILLER_49_129 ();
 sg13g2_fill_2 FILLER_49_166 ();
 sg13g2_fill_1 FILLER_49_168 ();
 sg13g2_fill_2 FILLER_49_240 ();
 sg13g2_fill_1 FILLER_49_242 ();
 sg13g2_fill_1 FILLER_49_252 ();
 sg13g2_fill_1 FILLER_49_262 ();
 sg13g2_fill_1 FILLER_49_290 ();
 sg13g2_fill_2 FILLER_49_324 ();
 sg13g2_fill_2 FILLER_49_358 ();
 sg13g2_fill_1 FILLER_49_360 ();
 sg13g2_fill_1 FILLER_49_462 ();
 sg13g2_fill_2 FILLER_49_472 ();
 sg13g2_fill_1 FILLER_49_474 ();
 sg13g2_fill_2 FILLER_49_511 ();
 sg13g2_fill_2 FILLER_49_535 ();
 sg13g2_fill_1 FILLER_49_653 ();
 sg13g2_fill_1 FILLER_49_671 ();
 sg13g2_fill_2 FILLER_49_707 ();
 sg13g2_decap_4 FILLER_49_713 ();
 sg13g2_fill_1 FILLER_49_717 ();
 sg13g2_decap_4 FILLER_49_722 ();
 sg13g2_fill_2 FILLER_49_732 ();
 sg13g2_fill_1 FILLER_49_753 ();
 sg13g2_fill_1 FILLER_49_785 ();
 sg13g2_fill_1 FILLER_49_803 ();
 sg13g2_decap_4 FILLER_49_849 ();
 sg13g2_fill_2 FILLER_49_853 ();
 sg13g2_fill_2 FILLER_49_864 ();
 sg13g2_fill_2 FILLER_49_887 ();
 sg13g2_fill_1 FILLER_49_889 ();
 sg13g2_fill_1 FILLER_49_917 ();
 sg13g2_fill_2 FILLER_49_955 ();
 sg13g2_fill_1 FILLER_49_957 ();
 sg13g2_fill_2 FILLER_49_1002 ();
 sg13g2_fill_1 FILLER_49_1102 ();
 sg13g2_decap_4 FILLER_49_1181 ();
 sg13g2_fill_1 FILLER_49_1185 ();
 sg13g2_fill_1 FILLER_49_1247 ();
 sg13g2_fill_1 FILLER_49_1271 ();
 sg13g2_fill_1 FILLER_49_1299 ();
 sg13g2_fill_1 FILLER_49_1327 ();
 sg13g2_fill_1 FILLER_49_1338 ();
 sg13g2_decap_4 FILLER_49_1418 ();
 sg13g2_fill_1 FILLER_49_1500 ();
 sg13g2_fill_1 FILLER_49_1538 ();
 sg13g2_fill_1 FILLER_49_1574 ();
 sg13g2_fill_1 FILLER_49_1584 ();
 sg13g2_fill_2 FILLER_49_1597 ();
 sg13g2_fill_1 FILLER_49_1612 ();
 sg13g2_fill_1 FILLER_49_1626 ();
 sg13g2_fill_1 FILLER_49_1671 ();
 sg13g2_fill_1 FILLER_49_1675 ();
 sg13g2_fill_2 FILLER_49_1700 ();
 sg13g2_fill_2 FILLER_49_1725 ();
 sg13g2_fill_2 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_2 ();
 sg13g2_fill_1 FILLER_50_74 ();
 sg13g2_fill_2 FILLER_50_108 ();
 sg13g2_fill_1 FILLER_50_110 ();
 sg13g2_fill_2 FILLER_50_151 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_fill_1 FILLER_50_210 ();
 sg13g2_fill_2 FILLER_50_238 ();
 sg13g2_fill_1 FILLER_50_240 ();
 sg13g2_fill_2 FILLER_50_278 ();
 sg13g2_fill_1 FILLER_50_329 ();
 sg13g2_fill_1 FILLER_50_401 ();
 sg13g2_fill_1 FILLER_50_415 ();
 sg13g2_fill_1 FILLER_50_444 ();
 sg13g2_fill_2 FILLER_50_484 ();
 sg13g2_fill_1 FILLER_50_530 ();
 sg13g2_fill_1 FILLER_50_539 ();
 sg13g2_fill_1 FILLER_50_558 ();
 sg13g2_fill_2 FILLER_50_572 ();
 sg13g2_fill_1 FILLER_50_574 ();
 sg13g2_fill_2 FILLER_50_615 ();
 sg13g2_fill_1 FILLER_50_617 ();
 sg13g2_fill_1 FILLER_50_631 ();
 sg13g2_fill_2 FILLER_50_718 ();
 sg13g2_decap_4 FILLER_50_746 ();
 sg13g2_fill_2 FILLER_50_758 ();
 sg13g2_fill_2 FILLER_50_778 ();
 sg13g2_fill_1 FILLER_50_780 ();
 sg13g2_decap_8 FILLER_50_813 ();
 sg13g2_decap_8 FILLER_50_820 ();
 sg13g2_decap_4 FILLER_50_859 ();
 sg13g2_fill_1 FILLER_50_863 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_fill_2 FILLER_50_895 ();
 sg13g2_fill_2 FILLER_50_921 ();
 sg13g2_fill_2 FILLER_50_932 ();
 sg13g2_fill_2 FILLER_50_978 ();
 sg13g2_fill_1 FILLER_50_980 ();
 sg13g2_fill_2 FILLER_50_998 ();
 sg13g2_fill_1 FILLER_50_1000 ();
 sg13g2_fill_1 FILLER_50_1036 ();
 sg13g2_fill_1 FILLER_50_1066 ();
 sg13g2_fill_1 FILLER_50_1097 ();
 sg13g2_fill_1 FILLER_50_1152 ();
 sg13g2_fill_1 FILLER_50_1170 ();
 sg13g2_fill_1 FILLER_50_1179 ();
 sg13g2_fill_1 FILLER_50_1233 ();
 sg13g2_fill_2 FILLER_50_1248 ();
 sg13g2_fill_2 FILLER_50_1300 ();
 sg13g2_fill_1 FILLER_50_1307 ();
 sg13g2_fill_2 FILLER_50_1322 ();
 sg13g2_fill_1 FILLER_50_1324 ();
 sg13g2_fill_2 FILLER_50_1339 ();
 sg13g2_fill_1 FILLER_50_1341 ();
 sg13g2_fill_2 FILLER_50_1350 ();
 sg13g2_fill_2 FILLER_50_1419 ();
 sg13g2_fill_2 FILLER_50_1461 ();
 sg13g2_fill_1 FILLER_50_1472 ();
 sg13g2_fill_2 FILLER_50_1502 ();
 sg13g2_fill_2 FILLER_50_1517 ();
 sg13g2_fill_1 FILLER_50_1559 ();
 sg13g2_fill_1 FILLER_50_1579 ();
 sg13g2_fill_1 FILLER_50_1628 ();
 sg13g2_fill_1 FILLER_50_1674 ();
 sg13g2_fill_2 FILLER_50_1718 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_29 ();
 sg13g2_fill_2 FILLER_51_120 ();
 sg13g2_fill_1 FILLER_51_122 ();
 sg13g2_fill_2 FILLER_51_144 ();
 sg13g2_fill_2 FILLER_51_190 ();
 sg13g2_fill_1 FILLER_51_192 ();
 sg13g2_fill_2 FILLER_51_269 ();
 sg13g2_fill_1 FILLER_51_280 ();
 sg13g2_fill_1 FILLER_51_303 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_fill_2 FILLER_51_328 ();
 sg13g2_fill_2 FILLER_51_335 ();
 sg13g2_fill_1 FILLER_51_410 ();
 sg13g2_fill_1 FILLER_51_466 ();
 sg13g2_fill_2 FILLER_51_557 ();
 sg13g2_fill_1 FILLER_51_559 ();
 sg13g2_fill_1 FILLER_51_606 ();
 sg13g2_fill_1 FILLER_51_647 ();
 sg13g2_fill_2 FILLER_51_661 ();
 sg13g2_fill_1 FILLER_51_672 ();
 sg13g2_fill_2 FILLER_51_686 ();
 sg13g2_fill_1 FILLER_51_688 ();
 sg13g2_fill_1 FILLER_51_722 ();
 sg13g2_fill_2 FILLER_51_739 ();
 sg13g2_fill_1 FILLER_51_741 ();
 sg13g2_decap_4 FILLER_51_746 ();
 sg13g2_fill_2 FILLER_51_782 ();
 sg13g2_fill_1 FILLER_51_784 ();
 sg13g2_fill_2 FILLER_51_790 ();
 sg13g2_fill_1 FILLER_51_792 ();
 sg13g2_decap_4 FILLER_51_858 ();
 sg13g2_fill_2 FILLER_51_866 ();
 sg13g2_fill_2 FILLER_51_901 ();
 sg13g2_fill_2 FILLER_51_959 ();
 sg13g2_fill_2 FILLER_51_1087 ();
 sg13g2_fill_2 FILLER_51_1114 ();
 sg13g2_fill_2 FILLER_51_1137 ();
 sg13g2_fill_2 FILLER_51_1148 ();
 sg13g2_fill_2 FILLER_51_1194 ();
 sg13g2_fill_2 FILLER_51_1200 ();
 sg13g2_decap_8 FILLER_51_1246 ();
 sg13g2_fill_2 FILLER_51_1253 ();
 sg13g2_decap_4 FILLER_51_1258 ();
 sg13g2_fill_1 FILLER_51_1262 ();
 sg13g2_fill_1 FILLER_51_1290 ();
 sg13g2_fill_1 FILLER_51_1312 ();
 sg13g2_fill_2 FILLER_51_1394 ();
 sg13g2_fill_1 FILLER_51_1401 ();
 sg13g2_fill_1 FILLER_51_1410 ();
 sg13g2_decap_8 FILLER_51_1424 ();
 sg13g2_fill_1 FILLER_51_1431 ();
 sg13g2_fill_2 FILLER_51_1441 ();
 sg13g2_fill_2 FILLER_51_1463 ();
 sg13g2_fill_1 FILLER_51_1481 ();
 sg13g2_fill_1 FILLER_51_1494 ();
 sg13g2_fill_2 FILLER_51_1522 ();
 sg13g2_fill_2 FILLER_51_1576 ();
 sg13g2_fill_1 FILLER_51_1591 ();
 sg13g2_fill_1 FILLER_51_1601 ();
 sg13g2_fill_2 FILLER_51_1615 ();
 sg13g2_fill_1 FILLER_51_1617 ();
 sg13g2_fill_1 FILLER_51_1673 ();
 sg13g2_fill_2 FILLER_51_1686 ();
 sg13g2_fill_2 FILLER_51_1712 ();
 sg13g2_fill_1 FILLER_51_1748 ();
 sg13g2_fill_2 FILLER_51_1766 ();
 sg13g2_fill_1 FILLER_52_153 ();
 sg13g2_fill_1 FILLER_52_204 ();
 sg13g2_fill_2 FILLER_52_218 ();
 sg13g2_fill_1 FILLER_52_220 ();
 sg13g2_fill_2 FILLER_52_304 ();
 sg13g2_fill_1 FILLER_52_315 ();
 sg13g2_fill_2 FILLER_52_345 ();
 sg13g2_fill_2 FILLER_52_493 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_2 FILLER_52_505 ();
 sg13g2_fill_2 FILLER_52_618 ();
 sg13g2_fill_1 FILLER_52_620 ();
 sg13g2_fill_1 FILLER_52_652 ();
 sg13g2_fill_2 FILLER_52_677 ();
 sg13g2_decap_4 FILLER_52_706 ();
 sg13g2_fill_1 FILLER_52_710 ();
 sg13g2_fill_1 FILLER_52_715 ();
 sg13g2_fill_1 FILLER_52_721 ();
 sg13g2_fill_2 FILLER_52_751 ();
 sg13g2_fill_1 FILLER_52_753 ();
 sg13g2_fill_2 FILLER_52_775 ();
 sg13g2_decap_8 FILLER_52_786 ();
 sg13g2_fill_2 FILLER_52_793 ();
 sg13g2_fill_1 FILLER_52_795 ();
 sg13g2_decap_8 FILLER_52_813 ();
 sg13g2_decap_4 FILLER_52_820 ();
 sg13g2_fill_1 FILLER_52_824 ();
 sg13g2_fill_2 FILLER_52_835 ();
 sg13g2_decap_4 FILLER_52_843 ();
 sg13g2_fill_1 FILLER_52_879 ();
 sg13g2_fill_2 FILLER_52_886 ();
 sg13g2_fill_1 FILLER_52_888 ();
 sg13g2_fill_2 FILLER_52_902 ();
 sg13g2_fill_2 FILLER_52_974 ();
 sg13g2_fill_1 FILLER_52_990 ();
 sg13g2_fill_2 FILLER_52_1024 ();
 sg13g2_fill_1 FILLER_52_1038 ();
 sg13g2_fill_2 FILLER_52_1051 ();
 sg13g2_fill_2 FILLER_52_1059 ();
 sg13g2_fill_1 FILLER_52_1061 ();
 sg13g2_fill_1 FILLER_52_1102 ();
 sg13g2_fill_2 FILLER_52_1127 ();
 sg13g2_fill_1 FILLER_52_1183 ();
 sg13g2_fill_2 FILLER_52_1221 ();
 sg13g2_fill_2 FILLER_52_1340 ();
 sg13g2_fill_1 FILLER_52_1342 ();
 sg13g2_fill_2 FILLER_52_1402 ();
 sg13g2_fill_1 FILLER_52_1495 ();
 sg13g2_fill_2 FILLER_52_1509 ();
 sg13g2_fill_1 FILLER_52_1563 ();
 sg13g2_fill_1 FILLER_52_1576 ();
 sg13g2_fill_1 FILLER_52_1616 ();
 sg13g2_fill_1 FILLER_52_1656 ();
 sg13g2_fill_2 FILLER_52_1663 ();
 sg13g2_fill_2 FILLER_52_1705 ();
 sg13g2_fill_2 FILLER_52_1734 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_29 ();
 sg13g2_fill_2 FILLER_53_77 ();
 sg13g2_fill_1 FILLER_53_79 ();
 sg13g2_fill_2 FILLER_53_113 ();
 sg13g2_fill_1 FILLER_53_115 ();
 sg13g2_fill_2 FILLER_53_129 ();
 sg13g2_fill_2 FILLER_53_141 ();
 sg13g2_fill_1 FILLER_53_178 ();
 sg13g2_fill_2 FILLER_53_188 ();
 sg13g2_fill_1 FILLER_53_190 ();
 sg13g2_fill_2 FILLER_53_222 ();
 sg13g2_fill_2 FILLER_53_237 ();
 sg13g2_fill_1 FILLER_53_256 ();
 sg13g2_fill_2 FILLER_53_276 ();
 sg13g2_fill_1 FILLER_53_302 ();
 sg13g2_fill_2 FILLER_53_320 ();
 sg13g2_fill_1 FILLER_53_335 ();
 sg13g2_fill_1 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_421 ();
 sg13g2_fill_1 FILLER_53_445 ();
 sg13g2_fill_2 FILLER_53_473 ();
 sg13g2_fill_1 FILLER_53_479 ();
 sg13g2_fill_2 FILLER_53_574 ();
 sg13g2_fill_1 FILLER_53_576 ();
 sg13g2_fill_1 FILLER_53_613 ();
 sg13g2_fill_2 FILLER_53_646 ();
 sg13g2_fill_1 FILLER_53_648 ();
 sg13g2_fill_1 FILLER_53_686 ();
 sg13g2_fill_1 FILLER_53_700 ();
 sg13g2_fill_1 FILLER_53_718 ();
 sg13g2_fill_1 FILLER_53_724 ();
 sg13g2_fill_2 FILLER_53_756 ();
 sg13g2_decap_8 FILLER_53_784 ();
 sg13g2_fill_2 FILLER_53_791 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_fill_1 FILLER_53_879 ();
 sg13g2_fill_2 FILLER_53_911 ();
 sg13g2_fill_2 FILLER_53_940 ();
 sg13g2_fill_2 FILLER_53_977 ();
 sg13g2_fill_1 FILLER_53_979 ();
 sg13g2_fill_1 FILLER_53_1003 ();
 sg13g2_fill_1 FILLER_53_1018 ();
 sg13g2_fill_2 FILLER_53_1030 ();
 sg13g2_fill_1 FILLER_53_1087 ();
 sg13g2_fill_2 FILLER_53_1109 ();
 sg13g2_fill_2 FILLER_53_1180 ();
 sg13g2_decap_4 FILLER_53_1230 ();
 sg13g2_fill_2 FILLER_53_1234 ();
 sg13g2_fill_1 FILLER_53_1277 ();
 sg13g2_fill_1 FILLER_53_1321 ();
 sg13g2_fill_2 FILLER_53_1349 ();
 sg13g2_fill_1 FILLER_53_1378 ();
 sg13g2_fill_1 FILLER_53_1394 ();
 sg13g2_fill_2 FILLER_53_1442 ();
 sg13g2_fill_2 FILLER_53_1458 ();
 sg13g2_fill_2 FILLER_53_1473 ();
 sg13g2_fill_1 FILLER_53_1475 ();
 sg13g2_fill_1 FILLER_53_1494 ();
 sg13g2_fill_1 FILLER_53_1501 ();
 sg13g2_fill_2 FILLER_53_1646 ();
 sg13g2_fill_1 FILLER_53_1648 ();
 sg13g2_fill_2 FILLER_53_1681 ();
 sg13g2_fill_2 FILLER_53_1710 ();
 sg13g2_fill_2 FILLER_53_1716 ();
 sg13g2_fill_1 FILLER_53_1767 ();
 sg13g2_fill_1 FILLER_54_103 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_fill_2 FILLER_54_168 ();
 sg13g2_fill_1 FILLER_54_201 ();
 sg13g2_fill_2 FILLER_54_322 ();
 sg13g2_fill_1 FILLER_54_324 ();
 sg13g2_fill_2 FILLER_54_343 ();
 sg13g2_fill_2 FILLER_54_376 ();
 sg13g2_fill_1 FILLER_54_378 ();
 sg13g2_fill_2 FILLER_54_424 ();
 sg13g2_fill_2 FILLER_54_486 ();
 sg13g2_fill_1 FILLER_54_514 ();
 sg13g2_fill_1 FILLER_54_628 ();
 sg13g2_fill_2 FILLER_54_661 ();
 sg13g2_fill_2 FILLER_54_677 ();
 sg13g2_fill_1 FILLER_54_679 ();
 sg13g2_fill_1 FILLER_54_695 ();
 sg13g2_fill_2 FILLER_54_714 ();
 sg13g2_decap_8 FILLER_54_725 ();
 sg13g2_decap_8 FILLER_54_732 ();
 sg13g2_fill_1 FILLER_54_739 ();
 sg13g2_fill_2 FILLER_54_744 ();
 sg13g2_fill_1 FILLER_54_746 ();
 sg13g2_decap_4 FILLER_54_791 ();
 sg13g2_fill_2 FILLER_54_795 ();
 sg13g2_fill_2 FILLER_54_871 ();
 sg13g2_fill_1 FILLER_54_873 ();
 sg13g2_fill_2 FILLER_54_891 ();
 sg13g2_fill_1 FILLER_54_893 ();
 sg13g2_fill_2 FILLER_54_912 ();
 sg13g2_fill_2 FILLER_54_1002 ();
 sg13g2_fill_1 FILLER_54_1004 ();
 sg13g2_fill_2 FILLER_54_1018 ();
 sg13g2_fill_1 FILLER_54_1033 ();
 sg13g2_fill_2 FILLER_54_1039 ();
 sg13g2_fill_1 FILLER_54_1046 ();
 sg13g2_fill_1 FILLER_54_1100 ();
 sg13g2_fill_1 FILLER_54_1155 ();
 sg13g2_fill_2 FILLER_54_1184 ();
 sg13g2_fill_1 FILLER_54_1186 ();
 sg13g2_fill_2 FILLER_54_1256 ();
 sg13g2_fill_1 FILLER_54_1263 ();
 sg13g2_fill_1 FILLER_54_1333 ();
 sg13g2_fill_1 FILLER_54_1337 ();
 sg13g2_fill_2 FILLER_54_1366 ();
 sg13g2_fill_1 FILLER_54_1409 ();
 sg13g2_fill_2 FILLER_54_1480 ();
 sg13g2_fill_1 FILLER_54_1513 ();
 sg13g2_fill_1 FILLER_54_1527 ();
 sg13g2_fill_1 FILLER_54_1567 ();
 sg13g2_fill_1 FILLER_54_1643 ();
 sg13g2_fill_1 FILLER_54_1665 ();
 sg13g2_fill_1 FILLER_54_1684 ();
 sg13g2_fill_1 FILLER_54_1712 ();
 sg13g2_fill_2 FILLER_54_1718 ();
 sg13g2_fill_2 FILLER_54_1731 ();
 sg13g2_fill_1 FILLER_54_1767 ();
 sg13g2_fill_2 FILLER_55_31 ();
 sg13g2_fill_2 FILLER_55_68 ();
 sg13g2_fill_1 FILLER_55_70 ();
 sg13g2_fill_2 FILLER_55_86 ();
 sg13g2_fill_2 FILLER_55_160 ();
 sg13g2_fill_2 FILLER_55_171 ();
 sg13g2_fill_1 FILLER_55_173 ();
 sg13g2_fill_2 FILLER_55_188 ();
 sg13g2_fill_1 FILLER_55_190 ();
 sg13g2_fill_2 FILLER_55_250 ();
 sg13g2_fill_1 FILLER_55_252 ();
 sg13g2_fill_1 FILLER_55_349 ();
 sg13g2_fill_1 FILLER_55_356 ();
 sg13g2_fill_2 FILLER_55_372 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_fill_2 FILLER_55_387 ();
 sg13g2_fill_1 FILLER_55_389 ();
 sg13g2_fill_2 FILLER_55_419 ();
 sg13g2_fill_2 FILLER_55_430 ();
 sg13g2_fill_1 FILLER_55_432 ();
 sg13g2_fill_1 FILLER_55_555 ();
 sg13g2_fill_2 FILLER_55_569 ();
 sg13g2_fill_1 FILLER_55_649 ();
 sg13g2_fill_1 FILLER_55_659 ();
 sg13g2_fill_2 FILLER_55_700 ();
 sg13g2_decap_4 FILLER_55_801 ();
 sg13g2_fill_1 FILLER_55_805 ();
 sg13g2_fill_1 FILLER_55_841 ();
 sg13g2_fill_2 FILLER_55_877 ();
 sg13g2_fill_1 FILLER_55_879 ();
 sg13g2_fill_2 FILLER_55_917 ();
 sg13g2_fill_1 FILLER_55_919 ();
 sg13g2_fill_2 FILLER_55_948 ();
 sg13g2_fill_2 FILLER_55_978 ();
 sg13g2_fill_2 FILLER_55_1086 ();
 sg13g2_fill_2 FILLER_55_1155 ();
 sg13g2_decap_8 FILLER_55_1197 ();
 sg13g2_fill_2 FILLER_55_1219 ();
 sg13g2_decap_8 FILLER_55_1234 ();
 sg13g2_decap_4 FILLER_55_1241 ();
 sg13g2_fill_1 FILLER_55_1245 ();
 sg13g2_fill_2 FILLER_55_1284 ();
 sg13g2_fill_2 FILLER_55_1291 ();
 sg13g2_fill_1 FILLER_55_1339 ();
 sg13g2_fill_2 FILLER_55_1345 ();
 sg13g2_fill_2 FILLER_55_1360 ();
 sg13g2_fill_2 FILLER_55_1366 ();
 sg13g2_fill_2 FILLER_55_1430 ();
 sg13g2_fill_2 FILLER_55_1462 ();
 sg13g2_fill_1 FILLER_55_1486 ();
 sg13g2_fill_1 FILLER_55_1495 ();
 sg13g2_fill_1 FILLER_55_1508 ();
 sg13g2_fill_1 FILLER_55_1545 ();
 sg13g2_fill_2 FILLER_55_1565 ();
 sg13g2_fill_2 FILLER_55_1602 ();
 sg13g2_fill_1 FILLER_55_1617 ();
 sg13g2_fill_1 FILLER_55_1651 ();
 sg13g2_fill_2 FILLER_55_1711 ();
 sg13g2_fill_2 FILLER_55_1766 ();
 sg13g2_fill_2 FILLER_56_27 ();
 sg13g2_fill_1 FILLER_56_29 ();
 sg13g2_fill_2 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_78 ();
 sg13g2_fill_2 FILLER_56_106 ();
 sg13g2_fill_1 FILLER_56_108 ();
 sg13g2_fill_1 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_156 ();
 sg13g2_fill_1 FILLER_56_158 ();
 sg13g2_fill_2 FILLER_56_191 ();
 sg13g2_fill_1 FILLER_56_210 ();
 sg13g2_fill_1 FILLER_56_244 ();
 sg13g2_fill_2 FILLER_56_267 ();
 sg13g2_fill_2 FILLER_56_296 ();
 sg13g2_fill_1 FILLER_56_298 ();
 sg13g2_fill_1 FILLER_56_311 ();
 sg13g2_fill_2 FILLER_56_321 ();
 sg13g2_fill_2 FILLER_56_341 ();
 sg13g2_fill_1 FILLER_56_343 ();
 sg13g2_fill_2 FILLER_56_368 ();
 sg13g2_fill_2 FILLER_56_415 ();
 sg13g2_fill_1 FILLER_56_417 ();
 sg13g2_fill_2 FILLER_56_445 ();
 sg13g2_fill_2 FILLER_56_456 ();
 sg13g2_fill_1 FILLER_56_458 ();
 sg13g2_fill_2 FILLER_56_492 ();
 sg13g2_fill_2 FILLER_56_549 ();
 sg13g2_fill_2 FILLER_56_601 ();
 sg13g2_fill_1 FILLER_56_603 ();
 sg13g2_fill_2 FILLER_56_636 ();
 sg13g2_fill_2 FILLER_56_673 ();
 sg13g2_fill_1 FILLER_56_675 ();
 sg13g2_fill_2 FILLER_56_683 ();
 sg13g2_decap_8 FILLER_56_726 ();
 sg13g2_fill_2 FILLER_56_733 ();
 sg13g2_fill_1 FILLER_56_735 ();
 sg13g2_fill_2 FILLER_56_740 ();
 sg13g2_fill_1 FILLER_56_742 ();
 sg13g2_fill_2 FILLER_56_784 ();
 sg13g2_fill_1 FILLER_56_786 ();
 sg13g2_fill_2 FILLER_56_815 ();
 sg13g2_fill_2 FILLER_56_843 ();
 sg13g2_fill_1 FILLER_56_845 ();
 sg13g2_fill_2 FILLER_56_890 ();
 sg13g2_fill_1 FILLER_56_892 ();
 sg13g2_fill_1 FILLER_56_902 ();
 sg13g2_fill_1 FILLER_56_922 ();
 sg13g2_fill_1 FILLER_56_949 ();
 sg13g2_fill_2 FILLER_56_1027 ();
 sg13g2_fill_2 FILLER_56_1128 ();
 sg13g2_decap_4 FILLER_56_1183 ();
 sg13g2_decap_8 FILLER_56_1193 ();
 sg13g2_decap_4 FILLER_56_1200 ();
 sg13g2_fill_1 FILLER_56_1331 ();
 sg13g2_fill_2 FILLER_56_1502 ();
 sg13g2_fill_1 FILLER_56_1530 ();
 sg13g2_fill_2 FILLER_56_1582 ();
 sg13g2_fill_2 FILLER_56_1636 ();
 sg13g2_fill_1 FILLER_56_1662 ();
 sg13g2_fill_1 FILLER_56_1694 ();
 sg13g2_fill_2 FILLER_57_72 ();
 sg13g2_fill_2 FILLER_57_173 ();
 sg13g2_fill_2 FILLER_57_179 ();
 sg13g2_fill_1 FILLER_57_230 ();
 sg13g2_fill_2 FILLER_57_315 ();
 sg13g2_fill_1 FILLER_57_317 ();
 sg13g2_fill_2 FILLER_57_345 ();
 sg13g2_fill_1 FILLER_57_347 ();
 sg13g2_fill_2 FILLER_57_362 ();
 sg13g2_fill_1 FILLER_57_364 ();
 sg13g2_fill_2 FILLER_57_374 ();
 sg13g2_fill_1 FILLER_57_376 ();
 sg13g2_fill_1 FILLER_57_396 ();
 sg13g2_fill_2 FILLER_57_543 ();
 sg13g2_fill_1 FILLER_57_577 ();
 sg13g2_fill_1 FILLER_57_600 ();
 sg13g2_fill_2 FILLER_57_614 ();
 sg13g2_fill_1 FILLER_57_616 ();
 sg13g2_fill_2 FILLER_57_657 ();
 sg13g2_fill_2 FILLER_57_713 ();
 sg13g2_fill_1 FILLER_57_715 ();
 sg13g2_decap_8 FILLER_57_729 ();
 sg13g2_fill_1 FILLER_57_736 ();
 sg13g2_fill_2 FILLER_57_789 ();
 sg13g2_fill_1 FILLER_57_791 ();
 sg13g2_fill_1 FILLER_57_803 ();
 sg13g2_fill_1 FILLER_57_813 ();
 sg13g2_fill_1 FILLER_57_825 ();
 sg13g2_fill_1 FILLER_57_839 ();
 sg13g2_fill_2 FILLER_57_896 ();
 sg13g2_fill_1 FILLER_57_898 ();
 sg13g2_fill_1 FILLER_57_912 ();
 sg13g2_fill_2 FILLER_57_1078 ();
 sg13g2_decap_8 FILLER_57_1230 ();
 sg13g2_fill_1 FILLER_57_1279 ();
 sg13g2_fill_1 FILLER_57_1325 ();
 sg13g2_fill_1 FILLER_57_1331 ();
 sg13g2_fill_1 FILLER_57_1421 ();
 sg13g2_decap_4 FILLER_57_1443 ();
 sg13g2_fill_2 FILLER_57_1458 ();
 sg13g2_fill_1 FILLER_57_1506 ();
 sg13g2_fill_1 FILLER_57_1547 ();
 sg13g2_fill_2 FILLER_57_1553 ();
 sg13g2_fill_2 FILLER_57_1575 ();
 sg13g2_fill_1 FILLER_57_1614 ();
 sg13g2_fill_2 FILLER_57_1628 ();
 sg13g2_fill_2 FILLER_57_1643 ();
 sg13g2_fill_1 FILLER_57_1645 ();
 sg13g2_fill_1 FILLER_57_1731 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_29 ();
 sg13g2_fill_2 FILLER_58_44 ();
 sg13g2_fill_1 FILLER_58_110 ();
 sg13g2_fill_2 FILLER_58_120 ();
 sg13g2_fill_1 FILLER_58_135 ();
 sg13g2_fill_1 FILLER_58_154 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_fill_2 FILLER_58_207 ();
 sg13g2_fill_2 FILLER_58_222 ();
 sg13g2_fill_1 FILLER_58_260 ();
 sg13g2_fill_2 FILLER_58_270 ();
 sg13g2_fill_1 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_310 ();
 sg13g2_fill_2 FILLER_58_355 ();
 sg13g2_fill_1 FILLER_58_367 ();
 sg13g2_fill_2 FILLER_58_409 ();
 sg13g2_fill_2 FILLER_58_425 ();
 sg13g2_fill_1 FILLER_58_427 ();
 sg13g2_fill_2 FILLER_58_441 ();
 sg13g2_fill_1 FILLER_58_443 ();
 sg13g2_fill_2 FILLER_58_452 ();
 sg13g2_fill_2 FILLER_58_467 ();
 sg13g2_fill_1 FILLER_58_469 ();
 sg13g2_fill_2 FILLER_58_517 ();
 sg13g2_fill_1 FILLER_58_564 ();
 sg13g2_fill_2 FILLER_58_638 ();
 sg13g2_fill_1 FILLER_58_671 ();
 sg13g2_fill_2 FILLER_58_709 ();
 sg13g2_fill_2 FILLER_58_765 ();
 sg13g2_fill_1 FILLER_58_767 ();
 sg13g2_decap_8 FILLER_58_808 ();
 sg13g2_decap_4 FILLER_58_815 ();
 sg13g2_fill_2 FILLER_58_819 ();
 sg13g2_fill_2 FILLER_58_827 ();
 sg13g2_fill_1 FILLER_58_829 ();
 sg13g2_fill_2 FILLER_58_836 ();
 sg13g2_fill_1 FILLER_58_838 ();
 sg13g2_fill_1 FILLER_58_859 ();
 sg13g2_fill_1 FILLER_58_875 ();
 sg13g2_fill_1 FILLER_58_907 ();
 sg13g2_fill_2 FILLER_58_937 ();
 sg13g2_fill_2 FILLER_58_958 ();
 sg13g2_fill_2 FILLER_58_1011 ();
 sg13g2_fill_1 FILLER_58_1065 ();
 sg13g2_fill_1 FILLER_58_1093 ();
 sg13g2_decap_4 FILLER_58_1200 ();
 sg13g2_fill_1 FILLER_58_1204 ();
 sg13g2_fill_1 FILLER_58_1222 ();
 sg13g2_fill_1 FILLER_58_1254 ();
 sg13g2_fill_2 FILLER_58_1312 ();
 sg13g2_fill_2 FILLER_58_1341 ();
 sg13g2_fill_1 FILLER_58_1396 ();
 sg13g2_fill_2 FILLER_58_1442 ();
 sg13g2_fill_2 FILLER_58_1448 ();
 sg13g2_fill_2 FILLER_58_1577 ();
 sg13g2_fill_2 FILLER_58_1616 ();
 sg13g2_fill_1 FILLER_58_1704 ();
 sg13g2_fill_1 FILLER_58_1767 ();
 sg13g2_fill_2 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_79 ();
 sg13g2_fill_1 FILLER_59_130 ();
 sg13g2_fill_1 FILLER_59_226 ();
 sg13g2_fill_2 FILLER_59_260 ();
 sg13g2_fill_1 FILLER_59_262 ();
 sg13g2_fill_2 FILLER_59_292 ();
 sg13g2_fill_2 FILLER_59_342 ();
 sg13g2_fill_1 FILLER_59_381 ();
 sg13g2_fill_1 FILLER_59_432 ();
 sg13g2_fill_2 FILLER_59_460 ();
 sg13g2_fill_2 FILLER_59_579 ();
 sg13g2_fill_1 FILLER_59_581 ();
 sg13g2_fill_1 FILLER_59_591 ();
 sg13g2_fill_2 FILLER_59_600 ();
 sg13g2_fill_2 FILLER_59_611 ();
 sg13g2_fill_1 FILLER_59_617 ();
 sg13g2_fill_2 FILLER_59_622 ();
 sg13g2_fill_2 FILLER_59_646 ();
 sg13g2_fill_1 FILLER_59_648 ();
 sg13g2_fill_1 FILLER_59_666 ();
 sg13g2_fill_2 FILLER_59_672 ();
 sg13g2_fill_2 FILLER_59_701 ();
 sg13g2_fill_1 FILLER_59_703 ();
 sg13g2_fill_2 FILLER_59_763 ();
 sg13g2_decap_8 FILLER_59_805 ();
 sg13g2_fill_2 FILLER_59_862 ();
 sg13g2_fill_1 FILLER_59_864 ();
 sg13g2_fill_1 FILLER_59_874 ();
 sg13g2_fill_2 FILLER_59_892 ();
 sg13g2_fill_1 FILLER_59_926 ();
 sg13g2_fill_1 FILLER_59_931 ();
 sg13g2_fill_2 FILLER_59_999 ();
 sg13g2_fill_2 FILLER_59_1222 ();
 sg13g2_fill_1 FILLER_59_1328 ();
 sg13g2_fill_2 FILLER_59_1471 ();
 sg13g2_fill_2 FILLER_59_1490 ();
 sg13g2_fill_1 FILLER_59_1538 ();
 sg13g2_fill_1 FILLER_59_1560 ();
 sg13g2_fill_2 FILLER_59_1630 ();
 sg13g2_fill_1 FILLER_59_1670 ();
 sg13g2_fill_1 FILLER_59_1712 ();
 sg13g2_fill_2 FILLER_59_1739 ();
 sg13g2_fill_2 FILLER_60_47 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_fill_2 FILLER_60_96 ();
 sg13g2_fill_1 FILLER_60_158 ();
 sg13g2_fill_2 FILLER_60_236 ();
 sg13g2_fill_1 FILLER_60_238 ();
 sg13g2_fill_2 FILLER_60_398 ();
 sg13g2_fill_2 FILLER_60_414 ();
 sg13g2_fill_2 FILLER_60_421 ();
 sg13g2_fill_2 FILLER_60_491 ();
 sg13g2_fill_2 FILLER_60_510 ();
 sg13g2_fill_2 FILLER_60_526 ();
 sg13g2_fill_1 FILLER_60_528 ();
 sg13g2_fill_2 FILLER_60_555 ();
 sg13g2_fill_1 FILLER_60_673 ();
 sg13g2_fill_2 FILLER_60_696 ();
 sg13g2_fill_2 FILLER_60_715 ();
 sg13g2_fill_2 FILLER_60_768 ();
 sg13g2_fill_1 FILLER_60_770 ();
 sg13g2_fill_2 FILLER_60_799 ();
 sg13g2_fill_1 FILLER_60_801 ();
 sg13g2_fill_2 FILLER_60_827 ();
 sg13g2_fill_1 FILLER_60_829 ();
 sg13g2_fill_1 FILLER_60_844 ();
 sg13g2_fill_2 FILLER_60_909 ();
 sg13g2_fill_1 FILLER_60_911 ();
 sg13g2_fill_2 FILLER_60_921 ();
 sg13g2_fill_1 FILLER_60_923 ();
 sg13g2_fill_2 FILLER_60_968 ();
 sg13g2_fill_1 FILLER_60_998 ();
 sg13g2_fill_1 FILLER_60_1026 ();
 sg13g2_fill_1 FILLER_60_1054 ();
 sg13g2_fill_2 FILLER_60_1068 ();
 sg13g2_fill_1 FILLER_60_1201 ();
 sg13g2_fill_1 FILLER_60_1215 ();
 sg13g2_fill_1 FILLER_60_1234 ();
 sg13g2_fill_1 FILLER_60_1259 ();
 sg13g2_fill_2 FILLER_60_1265 ();
 sg13g2_fill_1 FILLER_60_1287 ();
 sg13g2_fill_1 FILLER_60_1327 ();
 sg13g2_fill_2 FILLER_60_1427 ();
 sg13g2_fill_1 FILLER_60_1456 ();
 sg13g2_fill_1 FILLER_60_1610 ();
 sg13g2_fill_1 FILLER_60_1617 ();
 sg13g2_fill_1 FILLER_60_1645 ();
 sg13g2_fill_1 FILLER_60_1713 ();
 sg13g2_fill_2 FILLER_60_1756 ();
 sg13g2_fill_2 FILLER_60_1766 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_30 ();
 sg13g2_fill_1 FILLER_61_107 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_2 FILLER_61_199 ();
 sg13g2_fill_2 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_298 ();
 sg13g2_fill_1 FILLER_61_300 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_fill_2 FILLER_61_361 ();
 sg13g2_fill_1 FILLER_61_434 ();
 sg13g2_fill_1 FILLER_61_455 ();
 sg13g2_fill_2 FILLER_61_498 ();
 sg13g2_fill_2 FILLER_61_510 ();
 sg13g2_fill_1 FILLER_61_522 ();
 sg13g2_fill_1 FILLER_61_552 ();
 sg13g2_fill_1 FILLER_61_593 ();
 sg13g2_fill_2 FILLER_61_670 ();
 sg13g2_fill_1 FILLER_61_672 ();
 sg13g2_fill_2 FILLER_61_761 ();
 sg13g2_fill_1 FILLER_61_763 ();
 sg13g2_fill_1 FILLER_61_803 ();
 sg13g2_fill_2 FILLER_61_810 ();
 sg13g2_fill_1 FILLER_61_852 ();
 sg13g2_fill_2 FILLER_61_881 ();
 sg13g2_fill_1 FILLER_61_883 ();
 sg13g2_fill_2 FILLER_61_942 ();
 sg13g2_fill_2 FILLER_61_967 ();
 sg13g2_fill_2 FILLER_61_995 ();
 sg13g2_fill_2 FILLER_61_1011 ();
 sg13g2_fill_1 FILLER_61_1027 ();
 sg13g2_fill_1 FILLER_61_1079 ();
 sg13g2_fill_2 FILLER_61_1151 ();
 sg13g2_fill_1 FILLER_61_1153 ();
 sg13g2_fill_1 FILLER_61_1190 ();
 sg13g2_fill_2 FILLER_61_1218 ();
 sg13g2_fill_1 FILLER_61_1220 ();
 sg13g2_fill_1 FILLER_61_1249 ();
 sg13g2_fill_2 FILLER_61_1274 ();
 sg13g2_fill_1 FILLER_61_1306 ();
 sg13g2_fill_2 FILLER_61_1329 ();
 sg13g2_fill_1 FILLER_61_1340 ();
 sg13g2_fill_1 FILLER_61_1351 ();
 sg13g2_fill_1 FILLER_61_1394 ();
 sg13g2_fill_2 FILLER_61_1423 ();
 sg13g2_fill_2 FILLER_61_1467 ();
 sg13g2_fill_1 FILLER_61_1469 ();
 sg13g2_fill_1 FILLER_61_1475 ();
 sg13g2_fill_1 FILLER_61_1494 ();
 sg13g2_fill_2 FILLER_61_1538 ();
 sg13g2_fill_2 FILLER_61_1546 ();
 sg13g2_fill_1 FILLER_61_1629 ();
 sg13g2_fill_1 FILLER_61_1643 ();
 sg13g2_fill_2 FILLER_61_1671 ();
 sg13g2_decap_8 FILLER_61_1676 ();
 sg13g2_fill_2 FILLER_61_1683 ();
 sg13g2_fill_1 FILLER_61_1685 ();
 sg13g2_fill_2 FILLER_61_1690 ();
 sg13g2_fill_2 FILLER_61_1707 ();
 sg13g2_fill_1 FILLER_61_1727 ();
 sg13g2_fill_1 FILLER_61_1767 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_1 FILLER_62_109 ();
 sg13g2_fill_2 FILLER_62_119 ();
 sg13g2_fill_1 FILLER_62_121 ();
 sg13g2_fill_1 FILLER_62_159 ();
 sg13g2_fill_1 FILLER_62_203 ();
 sg13g2_fill_2 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_316 ();
 sg13g2_fill_2 FILLER_62_330 ();
 sg13g2_fill_1 FILLER_62_363 ();
 sg13g2_fill_1 FILLER_62_373 ();
 sg13g2_fill_2 FILLER_62_482 ();
 sg13g2_fill_2 FILLER_62_533 ();
 sg13g2_fill_1 FILLER_62_576 ();
 sg13g2_fill_2 FILLER_62_630 ();
 sg13g2_fill_2 FILLER_62_680 ();
 sg13g2_fill_1 FILLER_62_701 ();
 sg13g2_fill_1 FILLER_62_738 ();
 sg13g2_fill_2 FILLER_62_811 ();
 sg13g2_fill_1 FILLER_62_813 ();
 sg13g2_fill_1 FILLER_62_820 ();
 sg13g2_fill_1 FILLER_62_845 ();
 sg13g2_fill_2 FILLER_62_882 ();
 sg13g2_fill_2 FILLER_62_889 ();
 sg13g2_fill_1 FILLER_62_1031 ();
 sg13g2_fill_1 FILLER_62_1047 ();
 sg13g2_fill_1 FILLER_62_1056 ();
 sg13g2_fill_2 FILLER_62_1100 ();
 sg13g2_fill_1 FILLER_62_1106 ();
 sg13g2_fill_2 FILLER_62_1162 ();
 sg13g2_fill_1 FILLER_62_1181 ();
 sg13g2_fill_1 FILLER_62_1205 ();
 sg13g2_fill_1 FILLER_62_1223 ();
 sg13g2_fill_1 FILLER_62_1279 ();
 sg13g2_fill_2 FILLER_62_1471 ();
 sg13g2_decap_4 FILLER_62_1673 ();
 sg13g2_fill_2 FILLER_62_1715 ();
 sg13g2_fill_1 FILLER_62_1758 ();
 sg13g2_fill_1 FILLER_62_1762 ();
 sg13g2_fill_2 FILLER_62_1766 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_46 ();
 sg13g2_fill_1 FILLER_63_79 ();
 sg13g2_fill_1 FILLER_63_94 ();
 sg13g2_fill_2 FILLER_63_132 ();
 sg13g2_fill_1 FILLER_63_134 ();
 sg13g2_fill_1 FILLER_63_196 ();
 sg13g2_fill_2 FILLER_63_242 ();
 sg13g2_fill_2 FILLER_63_272 ();
 sg13g2_fill_1 FILLER_63_348 ();
 sg13g2_fill_1 FILLER_63_379 ();
 sg13g2_fill_2 FILLER_63_397 ();
 sg13g2_fill_1 FILLER_63_399 ();
 sg13g2_fill_2 FILLER_63_463 ();
 sg13g2_fill_2 FILLER_63_487 ();
 sg13g2_fill_2 FILLER_63_509 ();
 sg13g2_fill_1 FILLER_63_519 ();
 sg13g2_fill_1 FILLER_63_578 ();
 sg13g2_fill_2 FILLER_63_594 ();
 sg13g2_fill_2 FILLER_63_629 ();
 sg13g2_fill_1 FILLER_63_650 ();
 sg13g2_fill_2 FILLER_63_676 ();
 sg13g2_fill_1 FILLER_63_678 ();
 sg13g2_fill_2 FILLER_63_712 ();
 sg13g2_fill_1 FILLER_63_782 ();
 sg13g2_fill_2 FILLER_63_801 ();
 sg13g2_fill_2 FILLER_63_809 ();
 sg13g2_fill_2 FILLER_63_856 ();
 sg13g2_fill_1 FILLER_63_858 ();
 sg13g2_fill_2 FILLER_63_887 ();
 sg13g2_fill_2 FILLER_63_950 ();
 sg13g2_fill_1 FILLER_63_952 ();
 sg13g2_fill_2 FILLER_63_977 ();
 sg13g2_fill_1 FILLER_63_979 ();
 sg13g2_fill_2 FILLER_63_1010 ();
 sg13g2_fill_1 FILLER_63_1079 ();
 sg13g2_fill_1 FILLER_63_1112 ();
 sg13g2_fill_2 FILLER_63_1122 ();
 sg13g2_fill_1 FILLER_63_1133 ();
 sg13g2_fill_2 FILLER_63_1167 ();
 sg13g2_fill_2 FILLER_63_1268 ();
 sg13g2_fill_1 FILLER_63_1310 ();
 sg13g2_fill_2 FILLER_63_1343 ();
 sg13g2_fill_1 FILLER_63_1381 ();
 sg13g2_fill_1 FILLER_63_1424 ();
 sg13g2_fill_1 FILLER_63_1511 ();
 sg13g2_fill_1 FILLER_63_1523 ();
 sg13g2_fill_2 FILLER_63_1541 ();
 sg13g2_fill_2 FILLER_63_1587 ();
 sg13g2_fill_1 FILLER_63_1651 ();
 sg13g2_decap_4 FILLER_63_1682 ();
 sg13g2_fill_1 FILLER_63_1686 ();
 sg13g2_fill_1 FILLER_63_1713 ();
 sg13g2_fill_1 FILLER_64_0 ();
 sg13g2_fill_2 FILLER_64_34 ();
 sg13g2_fill_2 FILLER_64_45 ();
 sg13g2_fill_2 FILLER_64_84 ();
 sg13g2_fill_1 FILLER_64_91 ();
 sg13g2_fill_2 FILLER_64_97 ();
 sg13g2_fill_1 FILLER_64_99 ();
 sg13g2_fill_2 FILLER_64_144 ();
 sg13g2_fill_1 FILLER_64_325 ();
 sg13g2_fill_1 FILLER_64_341 ();
 sg13g2_fill_1 FILLER_64_360 ();
 sg13g2_fill_2 FILLER_64_437 ();
 sg13g2_fill_2 FILLER_64_475 ();
 sg13g2_fill_2 FILLER_64_576 ();
 sg13g2_fill_1 FILLER_64_669 ();
 sg13g2_fill_2 FILLER_64_756 ();
 sg13g2_fill_1 FILLER_64_758 ();
 sg13g2_fill_2 FILLER_64_812 ();
 sg13g2_fill_2 FILLER_64_829 ();
 sg13g2_fill_1 FILLER_64_831 ();
 sg13g2_fill_2 FILLER_64_851 ();
 sg13g2_fill_1 FILLER_64_853 ();
 sg13g2_fill_1 FILLER_64_872 ();
 sg13g2_fill_1 FILLER_64_915 ();
 sg13g2_fill_1 FILLER_64_925 ();
 sg13g2_fill_1 FILLER_64_948 ();
 sg13g2_fill_2 FILLER_64_1004 ();
 sg13g2_fill_2 FILLER_64_1063 ();
 sg13g2_fill_2 FILLER_64_1111 ();
 sg13g2_fill_1 FILLER_64_1127 ();
 sg13g2_fill_2 FILLER_64_1142 ();
 sg13g2_fill_1 FILLER_64_1365 ();
 sg13g2_fill_1 FILLER_64_1409 ();
 sg13g2_fill_2 FILLER_64_1518 ();
 sg13g2_fill_1 FILLER_64_1551 ();
 sg13g2_fill_2 FILLER_64_1579 ();
 sg13g2_fill_2 FILLER_64_1608 ();
 sg13g2_fill_2 FILLER_64_1628 ();
 sg13g2_fill_1 FILLER_64_1634 ();
 sg13g2_fill_1 FILLER_64_1678 ();
 sg13g2_fill_1 FILLER_64_1718 ();
 sg13g2_fill_2 FILLER_64_1732 ();
 sg13g2_fill_2 FILLER_64_1751 ();
 sg13g2_fill_2 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_2 ();
 sg13g2_fill_2 FILLER_65_31 ();
 sg13g2_fill_1 FILLER_65_43 ();
 sg13g2_fill_2 FILLER_65_91 ();
 sg13g2_fill_1 FILLER_65_93 ();
 sg13g2_fill_1 FILLER_65_112 ();
 sg13g2_fill_1 FILLER_65_137 ();
 sg13g2_fill_2 FILLER_65_155 ();
 sg13g2_fill_2 FILLER_65_186 ();
 sg13g2_fill_2 FILLER_65_202 ();
 sg13g2_fill_2 FILLER_65_224 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_fill_2 FILLER_65_273 ();
 sg13g2_fill_2 FILLER_65_320 ();
 sg13g2_fill_2 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_347 ();
 sg13g2_fill_2 FILLER_65_375 ();
 sg13g2_fill_2 FILLER_65_390 ();
 sg13g2_fill_2 FILLER_65_414 ();
 sg13g2_fill_1 FILLER_65_430 ();
 sg13g2_fill_1 FILLER_65_509 ();
 sg13g2_fill_2 FILLER_65_524 ();
 sg13g2_fill_1 FILLER_65_540 ();
 sg13g2_fill_2 FILLER_65_560 ();
 sg13g2_fill_2 FILLER_65_571 ();
 sg13g2_fill_1 FILLER_65_590 ();
 sg13g2_fill_1 FILLER_65_605 ();
 sg13g2_fill_2 FILLER_65_643 ();
 sg13g2_fill_1 FILLER_65_812 ();
 sg13g2_fill_2 FILLER_65_841 ();
 sg13g2_fill_1 FILLER_65_843 ();
 sg13g2_fill_2 FILLER_65_924 ();
 sg13g2_fill_1 FILLER_65_926 ();
 sg13g2_fill_2 FILLER_65_959 ();
 sg13g2_fill_1 FILLER_65_1007 ();
 sg13g2_fill_2 FILLER_65_1022 ();
 sg13g2_fill_1 FILLER_65_1024 ();
 sg13g2_fill_2 FILLER_65_1070 ();
 sg13g2_fill_1 FILLER_65_1072 ();
 sg13g2_fill_1 FILLER_65_1172 ();
 sg13g2_fill_2 FILLER_65_1195 ();
 sg13g2_fill_1 FILLER_65_1218 ();
 sg13g2_fill_2 FILLER_65_1261 ();
 sg13g2_fill_1 FILLER_65_1291 ();
 sg13g2_fill_2 FILLER_65_1387 ();
 sg13g2_fill_2 FILLER_65_1433 ();
 sg13g2_fill_1 FILLER_65_1480 ();
 sg13g2_fill_1 FILLER_65_1596 ();
 sg13g2_fill_1 FILLER_65_1606 ();
 sg13g2_fill_1 FILLER_65_1679 ();
 sg13g2_decap_8 FILLER_65_1684 ();
 sg13g2_fill_2 FILLER_65_1691 ();
 sg13g2_fill_1 FILLER_65_1697 ();
 sg13g2_decap_8 FILLER_65_1711 ();
 sg13g2_decap_8 FILLER_65_1718 ();
 sg13g2_fill_2 FILLER_65_1725 ();
 sg13g2_fill_1 FILLER_65_1727 ();
 sg13g2_decap_8 FILLER_65_1735 ();
 sg13g2_decap_8 FILLER_65_1742 ();
 sg13g2_fill_2 FILLER_65_1749 ();
 sg13g2_fill_1 FILLER_65_1751 ();
 sg13g2_decap_8 FILLER_65_1761 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_1 FILLER_66_32 ();
 sg13g2_fill_2 FILLER_66_73 ();
 sg13g2_fill_2 FILLER_66_84 ();
 sg13g2_fill_2 FILLER_66_96 ();
 sg13g2_fill_2 FILLER_66_117 ();
 sg13g2_fill_1 FILLER_66_162 ();
 sg13g2_fill_1 FILLER_66_172 ();
 sg13g2_fill_1 FILLER_66_185 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_fill_1 FILLER_66_214 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_fill_1 FILLER_66_282 ();
 sg13g2_fill_1 FILLER_66_316 ();
 sg13g2_fill_2 FILLER_66_325 ();
 sg13g2_fill_2 FILLER_66_336 ();
 sg13g2_fill_2 FILLER_66_367 ();
 sg13g2_fill_2 FILLER_66_406 ();
 sg13g2_fill_1 FILLER_66_481 ();
 sg13g2_fill_1 FILLER_66_591 ();
 sg13g2_fill_2 FILLER_66_615 ();
 sg13g2_fill_1 FILLER_66_666 ();
 sg13g2_fill_2 FILLER_66_728 ();
 sg13g2_fill_2 FILLER_66_770 ();
 sg13g2_fill_1 FILLER_66_772 ();
 sg13g2_fill_1 FILLER_66_800 ();
 sg13g2_fill_2 FILLER_66_832 ();
 sg13g2_fill_1 FILLER_66_834 ();
 sg13g2_fill_2 FILLER_66_852 ();
 sg13g2_fill_1 FILLER_66_876 ();
 sg13g2_fill_1 FILLER_66_891 ();
 sg13g2_fill_2 FILLER_66_911 ();
 sg13g2_fill_2 FILLER_66_932 ();
 sg13g2_fill_1 FILLER_66_934 ();
 sg13g2_fill_2 FILLER_66_979 ();
 sg13g2_fill_2 FILLER_66_990 ();
 sg13g2_fill_1 FILLER_66_992 ();
 sg13g2_fill_2 FILLER_66_1034 ();
 sg13g2_fill_1 FILLER_66_1045 ();
 sg13g2_fill_2 FILLER_66_1090 ();
 sg13g2_fill_1 FILLER_66_1119 ();
 sg13g2_fill_1 FILLER_66_1143 ();
 sg13g2_fill_2 FILLER_66_1223 ();
 sg13g2_fill_2 FILLER_66_1275 ();
 sg13g2_fill_1 FILLER_66_1304 ();
 sg13g2_fill_2 FILLER_66_1674 ();
 sg13g2_fill_2 FILLER_66_1709 ();
 sg13g2_decap_8 FILLER_66_1724 ();
 sg13g2_decap_8 FILLER_66_1731 ();
 sg13g2_decap_8 FILLER_66_1738 ();
 sg13g2_decap_8 FILLER_66_1745 ();
 sg13g2_decap_8 FILLER_66_1752 ();
 sg13g2_decap_8 FILLER_66_1759 ();
 sg13g2_fill_2 FILLER_66_1766 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_54 ();
 sg13g2_fill_1 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_124 ();
 sg13g2_fill_1 FILLER_67_150 ();
 sg13g2_fill_1 FILLER_67_174 ();
 sg13g2_fill_1 FILLER_67_181 ();
 sg13g2_fill_2 FILLER_67_198 ();
 sg13g2_fill_2 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_267 ();
 sg13g2_fill_1 FILLER_67_446 ();
 sg13g2_fill_1 FILLER_67_470 ();
 sg13g2_fill_2 FILLER_67_510 ();
 sg13g2_fill_2 FILLER_67_603 ();
 sg13g2_fill_2 FILLER_67_637 ();
 sg13g2_fill_1 FILLER_67_658 ();
 sg13g2_fill_1 FILLER_67_673 ();
 sg13g2_fill_1 FILLER_67_701 ();
 sg13g2_fill_2 FILLER_67_724 ();
 sg13g2_fill_1 FILLER_67_739 ();
 sg13g2_fill_1 FILLER_67_749 ();
 sg13g2_fill_1 FILLER_67_776 ();
 sg13g2_fill_2 FILLER_67_814 ();
 sg13g2_fill_1 FILLER_67_816 ();
 sg13g2_fill_2 FILLER_67_889 ();
 sg13g2_fill_2 FILLER_67_948 ();
 sg13g2_fill_1 FILLER_67_950 ();
 sg13g2_fill_1 FILLER_67_960 ();
 sg13g2_fill_2 FILLER_67_967 ();
 sg13g2_fill_1 FILLER_67_969 ();
 sg13g2_fill_2 FILLER_67_1007 ();
 sg13g2_fill_1 FILLER_67_1009 ();
 sg13g2_fill_2 FILLER_67_1026 ();
 sg13g2_fill_1 FILLER_67_1145 ();
 sg13g2_fill_1 FILLER_67_1228 ();
 sg13g2_fill_2 FILLER_67_1267 ();
 sg13g2_fill_1 FILLER_67_1278 ();
 sg13g2_fill_1 FILLER_67_1301 ();
 sg13g2_fill_1 FILLER_67_1373 ();
 sg13g2_fill_2 FILLER_67_1391 ();
 sg13g2_fill_2 FILLER_67_1402 ();
 sg13g2_fill_1 FILLER_67_1474 ();
 sg13g2_fill_1 FILLER_67_1536 ();
 sg13g2_fill_2 FILLER_67_1542 ();
 sg13g2_fill_2 FILLER_67_1561 ();
 sg13g2_fill_1 FILLER_67_1586 ();
 sg13g2_fill_1 FILLER_67_1690 ();
 sg13g2_decap_8 FILLER_67_1703 ();
 sg13g2_decap_8 FILLER_67_1710 ();
 sg13g2_decap_8 FILLER_67_1717 ();
 sg13g2_decap_4 FILLER_67_1724 ();
 sg13g2_decap_8 FILLER_67_1731 ();
 sg13g2_decap_8 FILLER_67_1738 ();
 sg13g2_decap_8 FILLER_67_1745 ();
 sg13g2_decap_8 FILLER_67_1752 ();
 sg13g2_decap_8 FILLER_67_1759 ();
 sg13g2_fill_2 FILLER_67_1766 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_2 FILLER_68_91 ();
 sg13g2_fill_2 FILLER_68_111 ();
 sg13g2_fill_2 FILLER_68_123 ();
 sg13g2_fill_2 FILLER_68_134 ();
 sg13g2_fill_1 FILLER_68_178 ();
 sg13g2_fill_1 FILLER_68_212 ();
 sg13g2_fill_2 FILLER_68_385 ();
 sg13g2_fill_1 FILLER_68_446 ();
 sg13g2_fill_1 FILLER_68_530 ();
 sg13g2_fill_1 FILLER_68_589 ();
 sg13g2_fill_2 FILLER_68_626 ();
 sg13g2_fill_1 FILLER_68_637 ();
 sg13g2_fill_2 FILLER_68_657 ();
 sg13g2_fill_2 FILLER_68_677 ();
 sg13g2_fill_1 FILLER_68_683 ();
 sg13g2_fill_2 FILLER_68_739 ();
 sg13g2_fill_1 FILLER_68_794 ();
 sg13g2_fill_2 FILLER_68_816 ();
 sg13g2_fill_1 FILLER_68_818 ();
 sg13g2_fill_1 FILLER_68_875 ();
 sg13g2_fill_2 FILLER_68_890 ();
 sg13g2_fill_1 FILLER_68_892 ();
 sg13g2_fill_2 FILLER_68_901 ();
 sg13g2_fill_1 FILLER_68_903 ();
 sg13g2_fill_1 FILLER_68_940 ();
 sg13g2_fill_2 FILLER_68_987 ();
 sg13g2_fill_1 FILLER_68_989 ();
 sg13g2_fill_1 FILLER_68_999 ();
 sg13g2_fill_2 FILLER_68_1028 ();
 sg13g2_fill_2 FILLER_68_1047 ();
 sg13g2_fill_1 FILLER_68_1073 ();
 sg13g2_fill_2 FILLER_68_1116 ();
 sg13g2_fill_1 FILLER_68_1123 ();
 sg13g2_fill_1 FILLER_68_1256 ();
 sg13g2_fill_1 FILLER_68_1292 ();
 sg13g2_fill_1 FILLER_68_1409 ();
 sg13g2_fill_1 FILLER_68_1432 ();
 sg13g2_fill_2 FILLER_68_1459 ();
 sg13g2_fill_2 FILLER_68_1503 ();
 sg13g2_fill_2 FILLER_68_1515 ();
 sg13g2_fill_1 FILLER_68_1605 ();
 sg13g2_fill_1 FILLER_68_1614 ();
 sg13g2_fill_1 FILLER_68_1624 ();
 sg13g2_fill_2 FILLER_68_1661 ();
 sg13g2_fill_2 FILLER_68_1686 ();
 sg13g2_decap_8 FILLER_68_1695 ();
 sg13g2_decap_8 FILLER_68_1702 ();
 sg13g2_decap_8 FILLER_68_1709 ();
 sg13g2_decap_8 FILLER_68_1744 ();
 sg13g2_decap_8 FILLER_68_1751 ();
 sg13g2_decap_8 FILLER_68_1758 ();
 sg13g2_fill_2 FILLER_68_1765 ();
 sg13g2_fill_1 FILLER_68_1767 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_14 ();
 sg13g2_fill_2 FILLER_69_38 ();
 sg13g2_fill_1 FILLER_69_67 ();
 sg13g2_fill_2 FILLER_69_120 ();
 sg13g2_fill_2 FILLER_69_138 ();
 sg13g2_fill_1 FILLER_69_140 ();
 sg13g2_fill_2 FILLER_69_203 ();
 sg13g2_fill_2 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_263 ();
 sg13g2_fill_1 FILLER_69_313 ();
 sg13g2_fill_2 FILLER_69_350 ();
 sg13g2_fill_1 FILLER_69_384 ();
 sg13g2_fill_2 FILLER_69_390 ();
 sg13g2_fill_1 FILLER_69_413 ();
 sg13g2_fill_1 FILLER_69_428 ();
 sg13g2_fill_1 FILLER_69_467 ();
 sg13g2_fill_1 FILLER_69_496 ();
 sg13g2_fill_1 FILLER_69_548 ();
 sg13g2_fill_1 FILLER_69_576 ();
 sg13g2_fill_1 FILLER_69_583 ();
 sg13g2_fill_2 FILLER_69_673 ();
 sg13g2_fill_1 FILLER_69_721 ();
 sg13g2_fill_2 FILLER_69_768 ();
 sg13g2_fill_2 FILLER_69_824 ();
 sg13g2_fill_1 FILLER_69_840 ();
 sg13g2_fill_2 FILLER_69_879 ();
 sg13g2_fill_1 FILLER_69_890 ();
 sg13g2_fill_2 FILLER_69_907 ();
 sg13g2_fill_1 FILLER_69_930 ();
 sg13g2_fill_1 FILLER_69_939 ();
 sg13g2_fill_2 FILLER_69_949 ();
 sg13g2_fill_2 FILLER_69_1002 ();
 sg13g2_fill_1 FILLER_69_1137 ();
 sg13g2_fill_2 FILLER_69_1203 ();
 sg13g2_fill_2 FILLER_69_1257 ();
 sg13g2_fill_2 FILLER_69_1270 ();
 sg13g2_fill_2 FILLER_69_1378 ();
 sg13g2_fill_1 FILLER_69_1452 ();
 sg13g2_fill_2 FILLER_69_1494 ();
 sg13g2_fill_1 FILLER_69_1531 ();
 sg13g2_fill_1 FILLER_69_1584 ();
 sg13g2_fill_2 FILLER_69_1668 ();
 sg13g2_decap_4 FILLER_69_1700 ();
 sg13g2_fill_1 FILLER_69_1704 ();
 sg13g2_fill_1 FILLER_69_1733 ();
 sg13g2_fill_1 FILLER_70_0 ();
 sg13g2_fill_2 FILLER_70_45 ();
 sg13g2_fill_2 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_103 ();
 sg13g2_fill_1 FILLER_70_159 ();
 sg13g2_fill_1 FILLER_70_166 ();
 sg13g2_fill_2 FILLER_70_197 ();
 sg13g2_fill_1 FILLER_70_240 ();
 sg13g2_fill_1 FILLER_70_355 ();
 sg13g2_fill_2 FILLER_70_440 ();
 sg13g2_fill_1 FILLER_70_511 ();
 sg13g2_fill_2 FILLER_70_553 ();
 sg13g2_fill_2 FILLER_70_580 ();
 sg13g2_fill_1 FILLER_70_664 ();
 sg13g2_fill_1 FILLER_70_671 ();
 sg13g2_fill_1 FILLER_70_698 ();
 sg13g2_fill_2 FILLER_70_712 ();
 sg13g2_fill_1 FILLER_70_714 ();
 sg13g2_fill_1 FILLER_70_781 ();
 sg13g2_fill_1 FILLER_70_816 ();
 sg13g2_fill_2 FILLER_70_830 ();
 sg13g2_fill_2 FILLER_70_867 ();
 sg13g2_fill_2 FILLER_70_873 ();
 sg13g2_fill_1 FILLER_70_875 ();
 sg13g2_fill_2 FILLER_70_896 ();
 sg13g2_fill_2 FILLER_70_924 ();
 sg13g2_fill_1 FILLER_70_926 ();
 sg13g2_fill_2 FILLER_70_953 ();
 sg13g2_fill_1 FILLER_70_973 ();
 sg13g2_fill_2 FILLER_70_987 ();
 sg13g2_fill_1 FILLER_70_989 ();
 sg13g2_fill_1 FILLER_70_1058 ();
 sg13g2_fill_2 FILLER_70_1068 ();
 sg13g2_fill_1 FILLER_70_1070 ();
 sg13g2_fill_2 FILLER_70_1092 ();
 sg13g2_fill_2 FILLER_70_1113 ();
 sg13g2_fill_1 FILLER_70_1124 ();
 sg13g2_fill_1 FILLER_70_1166 ();
 sg13g2_fill_1 FILLER_70_1206 ();
 sg13g2_fill_1 FILLER_70_1251 ();
 sg13g2_fill_2 FILLER_70_1275 ();
 sg13g2_fill_2 FILLER_70_1295 ();
 sg13g2_fill_2 FILLER_70_1330 ();
 sg13g2_fill_1 FILLER_70_1397 ();
 sg13g2_fill_1 FILLER_70_1489 ();
 sg13g2_fill_2 FILLER_70_1555 ();
 sg13g2_fill_2 FILLER_70_1571 ();
 sg13g2_fill_1 FILLER_70_1612 ();
 sg13g2_fill_1 FILLER_70_1635 ();
 sg13g2_fill_1 FILLER_70_1654 ();
 sg13g2_fill_1 FILLER_70_1659 ();
 sg13g2_decap_4 FILLER_70_1752 ();
 sg13g2_fill_2 FILLER_70_1765 ();
 sg13g2_fill_1 FILLER_70_1767 ();
 sg13g2_fill_2 FILLER_71_45 ();
 sg13g2_fill_2 FILLER_71_75 ();
 sg13g2_fill_1 FILLER_71_138 ();
 sg13g2_fill_2 FILLER_71_200 ();
 sg13g2_fill_1 FILLER_71_309 ();
 sg13g2_fill_1 FILLER_71_336 ();
 sg13g2_fill_1 FILLER_71_350 ();
 sg13g2_fill_1 FILLER_71_474 ();
 sg13g2_fill_1 FILLER_71_578 ();
 sg13g2_fill_2 FILLER_71_595 ();
 sg13g2_fill_2 FILLER_71_657 ();
 sg13g2_fill_2 FILLER_71_776 ();
 sg13g2_fill_1 FILLER_71_790 ();
 sg13g2_fill_2 FILLER_71_859 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_fill_1 FILLER_71_890 ();
 sg13g2_fill_2 FILLER_71_900 ();
 sg13g2_fill_1 FILLER_71_902 ();
 sg13g2_fill_1 FILLER_71_920 ();
 sg13g2_fill_2 FILLER_71_938 ();
 sg13g2_fill_1 FILLER_71_940 ();
 sg13g2_fill_2 FILLER_71_1036 ();
 sg13g2_fill_1 FILLER_71_1150 ();
 sg13g2_fill_1 FILLER_71_1246 ();
 sg13g2_fill_2 FILLER_71_1266 ();
 sg13g2_fill_1 FILLER_71_1292 ();
 sg13g2_fill_1 FILLER_71_1303 ();
 sg13g2_fill_1 FILLER_71_1313 ();
 sg13g2_fill_1 FILLER_71_1349 ();
 sg13g2_fill_1 FILLER_71_1379 ();
 sg13g2_fill_2 FILLER_71_1454 ();
 sg13g2_fill_2 FILLER_71_1553 ();
 sg13g2_fill_1 FILLER_71_1588 ();
 sg13g2_fill_1 FILLER_71_1603 ();
 sg13g2_fill_2 FILLER_71_1626 ();
 sg13g2_fill_1 FILLER_71_1665 ();
 sg13g2_fill_2 FILLER_71_1678 ();
 sg13g2_fill_1 FILLER_72_0 ();
 sg13g2_fill_2 FILLER_72_148 ();
 sg13g2_fill_1 FILLER_72_236 ();
 sg13g2_fill_2 FILLER_72_260 ();
 sg13g2_fill_2 FILLER_72_308 ();
 sg13g2_fill_1 FILLER_72_331 ();
 sg13g2_fill_2 FILLER_72_392 ();
 sg13g2_fill_1 FILLER_72_548 ();
 sg13g2_fill_1 FILLER_72_689 ();
 sg13g2_fill_1 FILLER_72_703 ();
 sg13g2_fill_2 FILLER_72_727 ();
 sg13g2_fill_1 FILLER_72_729 ();
 sg13g2_fill_1 FILLER_72_808 ();
 sg13g2_fill_2 FILLER_72_841 ();
 sg13g2_fill_1 FILLER_72_843 ();
 sg13g2_fill_2 FILLER_72_873 ();
 sg13g2_fill_1 FILLER_72_875 ();
 sg13g2_fill_2 FILLER_72_920 ();
 sg13g2_fill_1 FILLER_72_922 ();
 sg13g2_fill_2 FILLER_72_960 ();
 sg13g2_fill_2 FILLER_72_984 ();
 sg13g2_fill_1 FILLER_72_1000 ();
 sg13g2_fill_1 FILLER_72_1006 ();
 sg13g2_fill_2 FILLER_72_1032 ();
 sg13g2_fill_1 FILLER_72_1043 ();
 sg13g2_fill_2 FILLER_72_1048 ();
 sg13g2_fill_1 FILLER_72_1050 ();
 sg13g2_fill_2 FILLER_72_1220 ();
 sg13g2_fill_1 FILLER_72_1237 ();
 sg13g2_fill_1 FILLER_72_1274 ();
 sg13g2_fill_2 FILLER_72_1367 ();
 sg13g2_fill_2 FILLER_72_1545 ();
 sg13g2_fill_2 FILLER_72_1614 ();
 sg13g2_fill_1 FILLER_72_1730 ();
 sg13g2_fill_1 FILLER_72_1767 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_56 ();
 sg13g2_fill_2 FILLER_73_79 ();
 sg13g2_fill_2 FILLER_73_108 ();
 sg13g2_fill_2 FILLER_73_124 ();
 sg13g2_fill_2 FILLER_73_148 ();
 sg13g2_fill_1 FILLER_73_186 ();
 sg13g2_fill_1 FILLER_73_286 ();
 sg13g2_fill_1 FILLER_73_320 ();
 sg13g2_fill_2 FILLER_73_375 ();
 sg13g2_fill_1 FILLER_73_391 ();
 sg13g2_fill_1 FILLER_73_398 ();
 sg13g2_fill_1 FILLER_73_432 ();
 sg13g2_fill_2 FILLER_73_447 ();
 sg13g2_fill_1 FILLER_73_490 ();
 sg13g2_fill_2 FILLER_73_515 ();
 sg13g2_fill_2 FILLER_73_523 ();
 sg13g2_fill_1 FILLER_73_535 ();
 sg13g2_fill_2 FILLER_73_555 ();
 sg13g2_fill_1 FILLER_73_571 ();
 sg13g2_fill_2 FILLER_73_628 ();
 sg13g2_fill_2 FILLER_73_667 ();
 sg13g2_fill_1 FILLER_73_697 ();
 sg13g2_fill_1 FILLER_73_718 ();
 sg13g2_fill_1 FILLER_73_804 ();
 sg13g2_fill_2 FILLER_73_811 ();
 sg13g2_fill_1 FILLER_73_846 ();
 sg13g2_fill_1 FILLER_73_872 ();
 sg13g2_fill_2 FILLER_73_886 ();
 sg13g2_fill_1 FILLER_73_897 ();
 sg13g2_fill_2 FILLER_73_933 ();
 sg13g2_fill_2 FILLER_73_956 ();
 sg13g2_fill_1 FILLER_73_967 ();
 sg13g2_fill_2 FILLER_73_1022 ();
 sg13g2_fill_2 FILLER_73_1043 ();
 sg13g2_fill_2 FILLER_73_1055 ();
 sg13g2_fill_2 FILLER_73_1097 ();
 sg13g2_fill_1 FILLER_73_1099 ();
 sg13g2_fill_1 FILLER_73_1113 ();
 sg13g2_fill_2 FILLER_73_1202 ();
 sg13g2_fill_2 FILLER_73_1249 ();
 sg13g2_fill_1 FILLER_73_1274 ();
 sg13g2_fill_1 FILLER_73_1281 ();
 sg13g2_fill_2 FILLER_73_1291 ();
 sg13g2_fill_1 FILLER_73_1301 ();
 sg13g2_fill_2 FILLER_73_1330 ();
 sg13g2_fill_1 FILLER_73_1482 ();
 sg13g2_fill_1 FILLER_73_1518 ();
 sg13g2_fill_1 FILLER_73_1572 ();
 sg13g2_fill_2 FILLER_73_1734 ();
 sg13g2_fill_1 FILLER_74_72 ();
 sg13g2_fill_1 FILLER_74_103 ();
 sg13g2_fill_1 FILLER_74_144 ();
 sg13g2_fill_2 FILLER_74_285 ();
 sg13g2_fill_2 FILLER_74_396 ();
 sg13g2_fill_1 FILLER_74_441 ();
 sg13g2_fill_2 FILLER_74_447 ();
 sg13g2_fill_2 FILLER_74_552 ();
 sg13g2_fill_1 FILLER_74_554 ();
 sg13g2_fill_2 FILLER_74_559 ();
 sg13g2_fill_2 FILLER_74_597 ();
 sg13g2_fill_2 FILLER_74_654 ();
 sg13g2_fill_1 FILLER_74_656 ();
 sg13g2_fill_1 FILLER_74_682 ();
 sg13g2_fill_1 FILLER_74_728 ();
 sg13g2_fill_2 FILLER_74_738 ();
 sg13g2_fill_1 FILLER_74_740 ();
 sg13g2_fill_2 FILLER_74_751 ();
 sg13g2_fill_1 FILLER_74_759 ();
 sg13g2_fill_2 FILLER_74_797 ();
 sg13g2_fill_2 FILLER_74_879 ();
 sg13g2_fill_1 FILLER_74_898 ();
 sg13g2_fill_1 FILLER_74_908 ();
 sg13g2_fill_1 FILLER_74_1004 ();
 sg13g2_fill_1 FILLER_74_1042 ();
 sg13g2_fill_2 FILLER_74_1052 ();
 sg13g2_fill_1 FILLER_74_1054 ();
 sg13g2_fill_1 FILLER_74_1081 ();
 sg13g2_fill_1 FILLER_74_1127 ();
 sg13g2_fill_1 FILLER_74_1141 ();
 sg13g2_fill_1 FILLER_74_1194 ();
 sg13g2_fill_2 FILLER_74_1200 ();
 sg13g2_fill_1 FILLER_74_1249 ();
 sg13g2_fill_1 FILLER_74_1317 ();
 sg13g2_fill_1 FILLER_74_1333 ();
 sg13g2_fill_1 FILLER_74_1417 ();
 sg13g2_fill_2 FILLER_74_1423 ();
 sg13g2_fill_1 FILLER_74_1466 ();
 sg13g2_fill_2 FILLER_74_1644 ();
 sg13g2_fill_1 FILLER_74_1683 ();
 sg13g2_fill_1 FILLER_74_1755 ();
 sg13g2_fill_2 FILLER_74_1765 ();
 sg13g2_fill_1 FILLER_74_1767 ();
 sg13g2_fill_1 FILLER_75_118 ();
 sg13g2_fill_2 FILLER_75_128 ();
 sg13g2_fill_2 FILLER_75_170 ();
 sg13g2_fill_1 FILLER_75_301 ();
 sg13g2_fill_2 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_349 ();
 sg13g2_fill_1 FILLER_75_393 ();
 sg13g2_fill_2 FILLER_75_416 ();
 sg13g2_fill_2 FILLER_75_465 ();
 sg13g2_fill_1 FILLER_75_467 ();
 sg13g2_fill_1 FILLER_75_486 ();
 sg13g2_fill_1 FILLER_75_509 ();
 sg13g2_fill_1 FILLER_75_528 ();
 sg13g2_fill_2 FILLER_75_542 ();
 sg13g2_fill_2 FILLER_75_569 ();
 sg13g2_fill_1 FILLER_75_598 ();
 sg13g2_fill_2 FILLER_75_608 ();
 sg13g2_fill_2 FILLER_75_623 ();
 sg13g2_fill_2 FILLER_75_679 ();
 sg13g2_fill_2 FILLER_75_745 ();
 sg13g2_fill_1 FILLER_75_747 ();
 sg13g2_fill_2 FILLER_75_775 ();
 sg13g2_fill_2 FILLER_75_809 ();
 sg13g2_fill_1 FILLER_75_876 ();
 sg13g2_fill_1 FILLER_75_914 ();
 sg13g2_fill_1 FILLER_75_919 ();
 sg13g2_fill_2 FILLER_75_945 ();
 sg13g2_fill_1 FILLER_75_947 ();
 sg13g2_fill_1 FILLER_75_974 ();
 sg13g2_fill_1 FILLER_75_990 ();
 sg13g2_fill_1 FILLER_75_996 ();
 sg13g2_fill_2 FILLER_75_1019 ();
 sg13g2_fill_1 FILLER_75_1056 ();
 sg13g2_fill_2 FILLER_75_1076 ();
 sg13g2_fill_1 FILLER_75_1078 ();
 sg13g2_fill_1 FILLER_75_1097 ();
 sg13g2_fill_1 FILLER_75_1122 ();
 sg13g2_fill_2 FILLER_75_1136 ();
 sg13g2_fill_2 FILLER_75_1151 ();
 sg13g2_fill_2 FILLER_75_1160 ();
 sg13g2_fill_2 FILLER_75_1258 ();
 sg13g2_fill_1 FILLER_75_1260 ();
 sg13g2_fill_1 FILLER_75_1287 ();
 sg13g2_fill_2 FILLER_75_1371 ();
 sg13g2_fill_1 FILLER_75_1450 ();
 sg13g2_fill_1 FILLER_75_1532 ();
 sg13g2_fill_1 FILLER_75_1569 ();
 sg13g2_fill_2 FILLER_75_1610 ();
 sg13g2_fill_2 FILLER_75_1622 ();
 sg13g2_fill_1 FILLER_75_1658 ();
 sg13g2_fill_1 FILLER_75_1689 ();
 sg13g2_fill_2 FILLER_75_1765 ();
 sg13g2_fill_1 FILLER_75_1767 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_58 ();
 sg13g2_fill_1 FILLER_76_89 ();
 sg13g2_fill_1 FILLER_76_98 ();
 sg13g2_fill_1 FILLER_76_136 ();
 sg13g2_fill_2 FILLER_76_187 ();
 sg13g2_fill_1 FILLER_76_239 ();
 sg13g2_fill_1 FILLER_76_254 ();
 sg13g2_fill_2 FILLER_76_268 ();
 sg13g2_fill_1 FILLER_76_335 ();
 sg13g2_fill_1 FILLER_76_342 ();
 sg13g2_fill_1 FILLER_76_355 ();
 sg13g2_fill_1 FILLER_76_439 ();
 sg13g2_fill_1 FILLER_76_458 ();
 sg13g2_fill_2 FILLER_76_494 ();
 sg13g2_fill_2 FILLER_76_574 ();
 sg13g2_fill_1 FILLER_76_576 ();
 sg13g2_fill_1 FILLER_76_586 ();
 sg13g2_fill_2 FILLER_76_596 ();
 sg13g2_fill_2 FILLER_76_679 ();
 sg13g2_fill_1 FILLER_76_681 ();
 sg13g2_fill_1 FILLER_76_687 ();
 sg13g2_fill_2 FILLER_76_710 ();
 sg13g2_fill_1 FILLER_76_712 ();
 sg13g2_fill_2 FILLER_76_759 ();
 sg13g2_fill_1 FILLER_76_766 ();
 sg13g2_fill_2 FILLER_76_777 ();
 sg13g2_fill_2 FILLER_76_792 ();
 sg13g2_fill_1 FILLER_76_803 ();
 sg13g2_fill_2 FILLER_76_841 ();
 sg13g2_fill_1 FILLER_76_843 ();
 sg13g2_fill_2 FILLER_76_900 ();
 sg13g2_fill_1 FILLER_76_902 ();
 sg13g2_fill_1 FILLER_76_912 ();
 sg13g2_fill_1 FILLER_76_1118 ();
 sg13g2_fill_2 FILLER_76_1181 ();
 sg13g2_fill_1 FILLER_76_1226 ();
 sg13g2_fill_1 FILLER_76_1242 ();
 sg13g2_fill_1 FILLER_76_1300 ();
 sg13g2_fill_1 FILLER_76_1307 ();
 sg13g2_fill_2 FILLER_76_1327 ();
 sg13g2_fill_2 FILLER_76_1338 ();
 sg13g2_fill_1 FILLER_76_1389 ();
 sg13g2_fill_2 FILLER_76_1399 ();
 sg13g2_fill_1 FILLER_76_1437 ();
 sg13g2_fill_1 FILLER_76_1483 ();
 sg13g2_fill_1 FILLER_76_1515 ();
 sg13g2_fill_2 FILLER_76_1588 ();
 sg13g2_fill_1 FILLER_76_1612 ();
 sg13g2_fill_1 FILLER_76_1618 ();
 sg13g2_fill_1 FILLER_76_1728 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_40 ();
 sg13g2_fill_2 FILLER_77_76 ();
 sg13g2_fill_2 FILLER_77_332 ();
 sg13g2_fill_1 FILLER_77_340 ();
 sg13g2_fill_2 FILLER_77_350 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_fill_1 FILLER_77_389 ();
 sg13g2_fill_2 FILLER_77_485 ();
 sg13g2_fill_1 FILLER_77_493 ();
 sg13g2_fill_1 FILLER_77_533 ();
 sg13g2_fill_1 FILLER_77_570 ();
 sg13g2_fill_2 FILLER_77_603 ();
 sg13g2_fill_1 FILLER_77_605 ();
 sg13g2_fill_1 FILLER_77_691 ();
 sg13g2_fill_2 FILLER_77_743 ();
 sg13g2_fill_1 FILLER_77_783 ();
 sg13g2_fill_2 FILLER_77_793 ();
 sg13g2_fill_2 FILLER_77_829 ();
 sg13g2_fill_1 FILLER_77_831 ();
 sg13g2_fill_1 FILLER_77_845 ();
 sg13g2_fill_2 FILLER_77_855 ();
 sg13g2_fill_1 FILLER_77_857 ();
 sg13g2_fill_2 FILLER_77_895 ();
 sg13g2_fill_2 FILLER_77_911 ();
 sg13g2_fill_2 FILLER_77_926 ();
 sg13g2_fill_1 FILLER_77_969 ();
 sg13g2_fill_2 FILLER_77_1003 ();
 sg13g2_fill_1 FILLER_77_1018 ();
 sg13g2_fill_1 FILLER_77_1033 ();
 sg13g2_fill_1 FILLER_77_1049 ();
 sg13g2_fill_1 FILLER_77_1063 ();
 sg13g2_fill_1 FILLER_77_1197 ();
 sg13g2_fill_2 FILLER_77_1238 ();
 sg13g2_fill_2 FILLER_77_1278 ();
 sg13g2_fill_2 FILLER_77_1317 ();
 sg13g2_fill_2 FILLER_77_1361 ();
 sg13g2_fill_1 FILLER_77_1400 ();
 sg13g2_fill_1 FILLER_77_1521 ();
 sg13g2_fill_2 FILLER_77_1554 ();
 sg13g2_fill_1 FILLER_77_1635 ();
 sg13g2_fill_2 FILLER_77_1693 ();
 sg13g2_fill_2 FILLER_77_1723 ();
 sg13g2_fill_1 FILLER_78_88 ();
 sg13g2_fill_2 FILLER_78_137 ();
 sg13g2_fill_2 FILLER_78_156 ();
 sg13g2_fill_2 FILLER_78_171 ();
 sg13g2_fill_1 FILLER_78_191 ();
 sg13g2_fill_2 FILLER_78_201 ();
 sg13g2_fill_1 FILLER_78_215 ();
 sg13g2_fill_2 FILLER_78_270 ();
 sg13g2_fill_1 FILLER_78_313 ();
 sg13g2_fill_2 FILLER_78_433 ();
 sg13g2_fill_1 FILLER_78_449 ();
 sg13g2_fill_2 FILLER_78_468 ();
 sg13g2_fill_2 FILLER_78_506 ();
 sg13g2_fill_2 FILLER_78_557 ();
 sg13g2_fill_2 FILLER_78_622 ();
 sg13g2_fill_1 FILLER_78_661 ();
 sg13g2_fill_1 FILLER_78_693 ();
 sg13g2_fill_2 FILLER_78_703 ();
 sg13g2_fill_1 FILLER_78_705 ();
 sg13g2_fill_1 FILLER_78_725 ();
 sg13g2_fill_2 FILLER_78_748 ();
 sg13g2_fill_2 FILLER_78_767 ();
 sg13g2_fill_1 FILLER_78_769 ();
 sg13g2_fill_2 FILLER_78_780 ();
 sg13g2_fill_1 FILLER_78_782 ();
 sg13g2_fill_2 FILLER_78_810 ();
 sg13g2_fill_1 FILLER_78_812 ();
 sg13g2_fill_1 FILLER_78_818 ();
 sg13g2_fill_2 FILLER_78_921 ();
 sg13g2_fill_1 FILLER_78_923 ();
 sg13g2_fill_1 FILLER_78_932 ();
 sg13g2_fill_2 FILLER_78_983 ();
 sg13g2_fill_1 FILLER_78_1014 ();
 sg13g2_fill_1 FILLER_78_1129 ();
 sg13g2_fill_1 FILLER_78_1141 ();
 sg13g2_fill_2 FILLER_78_1182 ();
 sg13g2_fill_1 FILLER_78_1264 ();
 sg13g2_fill_1 FILLER_78_1297 ();
 sg13g2_fill_1 FILLER_78_1325 ();
 sg13g2_fill_2 FILLER_78_1335 ();
 sg13g2_fill_2 FILLER_78_1386 ();
 sg13g2_fill_1 FILLER_78_1415 ();
 sg13g2_fill_2 FILLER_78_1550 ();
 sg13g2_fill_1 FILLER_78_1584 ();
 sg13g2_fill_1 FILLER_78_1617 ();
 sg13g2_fill_2 FILLER_78_1766 ();
 sg13g2_fill_2 FILLER_79_24 ();
 sg13g2_fill_1 FILLER_79_62 ();
 sg13g2_fill_1 FILLER_79_72 ();
 sg13g2_fill_1 FILLER_79_155 ();
 sg13g2_fill_1 FILLER_79_254 ();
 sg13g2_fill_2 FILLER_79_332 ();
 sg13g2_fill_1 FILLER_79_351 ();
 sg13g2_fill_2 FILLER_79_397 ();
 sg13g2_fill_2 FILLER_79_557 ();
 sg13g2_fill_2 FILLER_79_568 ();
 sg13g2_fill_1 FILLER_79_584 ();
 sg13g2_fill_2 FILLER_79_599 ();
 sg13g2_fill_1 FILLER_79_601 ();
 sg13g2_fill_1 FILLER_79_615 ();
 sg13g2_fill_1 FILLER_79_639 ();
 sg13g2_fill_2 FILLER_79_672 ();
 sg13g2_fill_1 FILLER_79_674 ();
 sg13g2_fill_2 FILLER_79_712 ();
 sg13g2_fill_2 FILLER_79_821 ();
 sg13g2_fill_1 FILLER_79_823 ();
 sg13g2_fill_2 FILLER_79_828 ();
 sg13g2_fill_1 FILLER_79_830 ();
 sg13g2_fill_2 FILLER_79_868 ();
 sg13g2_fill_2 FILLER_79_906 ();
 sg13g2_fill_2 FILLER_79_912 ();
 sg13g2_fill_1 FILLER_79_914 ();
 sg13g2_fill_2 FILLER_79_978 ();
 sg13g2_fill_2 FILLER_79_989 ();
 sg13g2_fill_2 FILLER_79_1000 ();
 sg13g2_fill_2 FILLER_79_1010 ();
 sg13g2_fill_1 FILLER_79_1039 ();
 sg13g2_fill_2 FILLER_79_1098 ();
 sg13g2_fill_1 FILLER_79_1127 ();
 sg13g2_fill_2 FILLER_79_1151 ();
 sg13g2_fill_2 FILLER_79_1234 ();
 sg13g2_fill_1 FILLER_79_1282 ();
 sg13g2_fill_2 FILLER_79_1314 ();
 sg13g2_fill_1 FILLER_79_1403 ();
 sg13g2_fill_2 FILLER_79_1606 ();
 sg13g2_fill_2 FILLER_79_1648 ();
 sg13g2_fill_2 FILLER_79_1699 ();
 sg13g2_decap_4 FILLER_79_1763 ();
 sg13g2_fill_1 FILLER_79_1767 ();
 sg13g2_fill_2 FILLER_80_115 ();
 sg13g2_fill_1 FILLER_80_130 ();
 sg13g2_fill_2 FILLER_80_152 ();
 sg13g2_fill_1 FILLER_80_207 ();
 sg13g2_fill_2 FILLER_80_321 ();
 sg13g2_fill_2 FILLER_80_480 ();
 sg13g2_fill_1 FILLER_80_529 ();
 sg13g2_fill_1 FILLER_80_575 ();
 sg13g2_fill_2 FILLER_80_604 ();
 sg13g2_fill_2 FILLER_80_637 ();
 sg13g2_fill_2 FILLER_80_676 ();
 sg13g2_fill_2 FILLER_80_738 ();
 sg13g2_fill_1 FILLER_80_740 ();
 sg13g2_fill_1 FILLER_80_768 ();
 sg13g2_fill_2 FILLER_80_783 ();
 sg13g2_fill_1 FILLER_80_812 ();
 sg13g2_fill_2 FILLER_80_863 ();
 sg13g2_fill_1 FILLER_80_873 ();
 sg13g2_fill_2 FILLER_80_886 ();
 sg13g2_fill_1 FILLER_80_888 ();
 sg13g2_decap_4 FILLER_80_897 ();
 sg13g2_fill_2 FILLER_80_901 ();
 sg13g2_fill_2 FILLER_80_931 ();
 sg13g2_fill_1 FILLER_80_969 ();
 sg13g2_fill_1 FILLER_80_1046 ();
 sg13g2_fill_1 FILLER_80_1364 ();
 sg13g2_fill_1 FILLER_80_1448 ();
 sg13g2_fill_2 FILLER_80_1458 ();
 sg13g2_fill_1 FILLER_80_1485 ();
 sg13g2_fill_1 FILLER_80_1538 ();
 sg13g2_fill_1 FILLER_80_1567 ();
 sg13g2_fill_2 FILLER_80_1717 ();
 sg13g2_fill_2 FILLER_80_1733 ();
 sg13g2_fill_1 FILLER_80_1735 ();
 sg13g2_fill_2 FILLER_80_1766 ();
endmodule
