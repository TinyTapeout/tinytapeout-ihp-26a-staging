VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tinymoa_ihp26a
  CLASS BLOCK ;
  FOREIGN tt_um_tinymoa_ihp26a ;
  ORIGIN 0.000 0.000 ;
  SIZE 1724.160 BY 313.740 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 21.580 3.150 23.780 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 60.450 3.150 62.650 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 99.320 3.150 101.520 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 138.190 3.150 140.390 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 177.060 3.150 179.260 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 215.930 3.150 218.130 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 254.800 3.150 257.000 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 293.670 3.150 295.870 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 332.540 3.150 334.740 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 371.410 3.150 373.610 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 410.280 3.150 412.480 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 449.150 3.150 451.350 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 488.020 3.150 490.220 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 526.890 3.150 529.090 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 565.760 3.150 567.960 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 604.630 3.150 606.830 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 643.500 3.150 645.700 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 682.370 3.150 684.570 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 721.240 3.150 723.440 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 760.110 3.150 762.310 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 798.980 3.150 801.180 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 837.850 3.150 840.050 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 876.720 3.150 878.920 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 915.590 3.150 917.790 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 954.460 3.150 956.660 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 993.330 3.150 995.530 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1032.200 3.150 1034.400 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1071.070 3.150 1073.270 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1109.940 3.150 1112.140 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1148.810 3.150 1151.010 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1187.680 3.150 1189.880 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1226.550 3.150 1228.750 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1265.420 3.150 1267.620 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1304.290 3.150 1306.490 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1343.160 3.150 1345.360 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1382.030 3.150 1384.230 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1420.900 3.150 1423.100 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1459.770 3.150 1461.970 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1498.640 3.150 1500.840 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1537.510 3.150 1539.710 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1576.380 3.150 1578.580 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1615.250 3.150 1617.450 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1654.120 3.150 1656.320 310.180 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1692.990 3.150 1695.190 310.180 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 15.380 3.560 17.580 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 54.250 3.560 56.450 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 93.120 3.560 95.320 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 131.990 3.560 134.190 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 170.860 3.560 173.060 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 209.730 3.560 211.930 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 248.600 3.560 250.800 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 287.470 3.560 289.670 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 326.340 3.560 328.540 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 365.210 3.560 367.410 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 404.080 3.560 406.280 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 442.950 3.560 445.150 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 481.820 3.560 484.020 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 520.690 3.560 522.890 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 559.560 3.560 561.760 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 598.430 3.560 600.630 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 637.300 3.560 639.500 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 676.170 3.560 678.370 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 715.040 3.560 717.240 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 753.910 3.560 756.110 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 792.780 3.560 794.980 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 831.650 3.560 833.850 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 870.520 3.560 872.720 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 909.390 3.560 911.590 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 948.260 3.560 950.460 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 987.130 3.560 989.330 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1026.000 3.560 1028.200 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1064.870 3.560 1067.070 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1103.740 3.560 1105.940 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1142.610 3.560 1144.810 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1181.480 3.560 1183.680 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1220.350 3.560 1222.550 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1259.220 3.560 1261.420 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1298.090 3.560 1300.290 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1336.960 3.560 1339.160 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1375.830 3.560 1378.030 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1414.700 3.560 1416.900 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1453.570 3.560 1455.770 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1492.440 3.560 1494.640 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1531.310 3.560 1533.510 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1570.180 3.560 1572.380 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1609.050 3.560 1611.250 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1647.920 3.560 1650.120 310.590 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 1686.790 3.560 1688.990 310.590 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal4 ;
        RECT 187.050 312.740 187.350 313.740 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 190.890 312.740 191.190 313.740 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal4 ;
        RECT 183.210 312.740 183.510 313.740 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal4 ;
        RECT 179.370 312.740 179.670 313.740 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal4 ;
        RECT 175.530 312.740 175.830 313.740 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 171.690 312.740 171.990 313.740 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 167.850 312.740 168.150 313.740 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 164.010 312.740 164.310 313.740 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 160.170 312.740 160.470 313.740 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 156.330 312.740 156.630 313.740 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 152.490 312.740 152.790 313.740 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 148.650 312.740 148.950 313.740 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 144.810 312.740 145.110 313.740 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 140.970 312.740 141.270 313.740 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 137.130 312.740 137.430 313.740 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 133.290 312.740 133.590 313.740 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 129.450 312.740 129.750 313.740 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 125.610 312.740 125.910 313.740 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal4 ;
        RECT 121.770 312.740 122.070 313.740 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 56.490 312.740 56.790 313.740 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 52.650 312.740 52.950 313.740 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 48.810 312.740 49.110 313.740 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 44.970 312.740 45.270 313.740 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 41.130 312.740 41.430 313.740 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 37.290 312.740 37.590 313.740 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 33.450 312.740 33.750 313.740 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 29.610 312.740 29.910 313.740 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 87.210 312.740 87.510 313.740 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 83.370 312.740 83.670 313.740 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 79.530 312.740 79.830 313.740 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 75.690 312.740 75.990 313.740 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 71.850 312.740 72.150 313.740 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 68.010 312.740 68.310 313.740 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 64.170 312.740 64.470 313.740 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal4 ;
        RECT 60.330 312.740 60.630 313.740 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.109200 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 117.930 312.740 118.230 313.740 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.109200 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 114.090 312.740 114.390 313.740 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.601400 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 110.250 312.740 110.550 313.740 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388200 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 106.410 312.740 106.710 313.740 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.289900 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 102.570 312.740 102.870 313.740 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.351000 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 98.730 312.740 99.030 313.740 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.109200 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 94.890 312.740 95.190 313.740 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.109200 ;
    ANTENNADIFFAREA 0.716100 ;
    PORT
      LAYER Metal4 ;
        RECT 91.050 312.740 91.350 313.740 ;
    END
  END uo_out[7]
  OBS
      LAYER GatPoly ;
        RECT 2.880 3.630 1721.280 310.110 ;
      LAYER Metal1 ;
        RECT 2.880 3.560 1721.280 310.180 ;
      LAYER Metal2 ;
        RECT 15.560 3.635 1695.010 310.105 ;
      LAYER Metal3 ;
        RECT 15.515 3.680 1695.055 310.060 ;
      LAYER Metal4 ;
        RECT 15.560 312.530 29.400 312.740 ;
        RECT 30.120 312.530 33.240 312.740 ;
        RECT 33.960 312.530 37.080 312.740 ;
        RECT 37.800 312.530 40.920 312.740 ;
        RECT 41.640 312.530 44.760 312.740 ;
        RECT 45.480 312.530 48.600 312.740 ;
        RECT 49.320 312.530 52.440 312.740 ;
        RECT 53.160 312.530 56.280 312.740 ;
        RECT 57.000 312.530 60.120 312.740 ;
        RECT 60.840 312.530 63.960 312.740 ;
        RECT 64.680 312.530 67.800 312.740 ;
        RECT 68.520 312.530 71.640 312.740 ;
        RECT 72.360 312.530 75.480 312.740 ;
        RECT 76.200 312.530 79.320 312.740 ;
        RECT 80.040 312.530 83.160 312.740 ;
        RECT 83.880 312.530 87.000 312.740 ;
        RECT 87.720 312.530 90.840 312.740 ;
        RECT 91.560 312.530 94.680 312.740 ;
        RECT 95.400 312.530 98.520 312.740 ;
        RECT 99.240 312.530 102.360 312.740 ;
        RECT 103.080 312.530 106.200 312.740 ;
        RECT 106.920 312.530 110.040 312.740 ;
        RECT 110.760 312.530 113.880 312.740 ;
        RECT 114.600 312.530 117.720 312.740 ;
        RECT 118.440 312.530 121.560 312.740 ;
        RECT 122.280 312.530 125.400 312.740 ;
        RECT 126.120 312.530 129.240 312.740 ;
        RECT 129.960 312.530 133.080 312.740 ;
        RECT 133.800 312.530 136.920 312.740 ;
        RECT 137.640 312.530 140.760 312.740 ;
        RECT 141.480 312.530 144.600 312.740 ;
        RECT 145.320 312.530 148.440 312.740 ;
        RECT 149.160 312.530 152.280 312.740 ;
        RECT 153.000 312.530 156.120 312.740 ;
        RECT 156.840 312.530 159.960 312.740 ;
        RECT 160.680 312.530 163.800 312.740 ;
        RECT 164.520 312.530 167.640 312.740 ;
        RECT 168.360 312.530 171.480 312.740 ;
        RECT 172.200 312.530 175.320 312.740 ;
        RECT 176.040 312.530 179.160 312.740 ;
        RECT 179.880 312.530 183.000 312.740 ;
        RECT 183.720 312.530 186.840 312.740 ;
        RECT 187.560 312.530 190.680 312.740 ;
        RECT 191.400 312.530 1695.010 312.740 ;
        RECT 15.560 3.635 1695.010 312.530 ;
      LAYER Metal5 ;
        RECT 15.515 3.470 1695.055 310.270 ;
  END
END tt_um_tinymoa_ihp26a
END LIBRARY

