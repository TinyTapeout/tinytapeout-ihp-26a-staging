module tt_um_hoene_smart_led_digital (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire \all_input_selector.counter0[0] ;
 wire \all_input_selector.counter0[1] ;
 wire \all_input_selector.counter0[2] ;
 wire \all_input_selector.counter0[3] ;
 wire \all_input_selector.counter0[4] ;
 wire \all_input_selector.counter0[5] ;
 wire \all_input_selector.counter1[0] ;
 wire \all_input_selector.counter1[1] ;
 wire \all_input_selector.counter1[2] ;
 wire \all_input_selector.counter1[3] ;
 wire \all_input_selector.counter1[4] ;
 wire \all_input_selector.counter1[5] ;
 wire \all_input_selector.counter1[6] ;
 wire \all_input_selector.counter1[7] ;
 wire \all_input_selector.in0selected ;
 wire \all_input_selector.last_in0 ;
 wire \all_input_selector.last_in1 ;
 wire \all_input_selector.out ;
 wire \all_low_pass_filter.last0 ;
 wire \all_low_pass_filter.last1 ;
 wire \all_low_pass_filter.out ;
 wire dout_data;
 wire dout_enable;
 wire manchester_decoder_out_clk;
 wire manchester_decoder_out_data;
 wire manchester_decoder_out_error;
 wire \protocol_counters_bits[0] ;
 wire \protocol_counters_bits[1] ;
 wire \protocol_counters_bits[2] ;
 wire \protocol_counters_bits[3] ;
 wire \protocol_counters_bits[4] ;
 wire protocol_counters_out_clk;
 wire protocol_counters_test_mode_out;
 wire protocol_insync_out;
 wire protocol_insync_out_clk;
 wire protocol_parity_error;
 wire clknet_0_clk;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire \user_manchester_decoder.counter[0] ;
 wire \user_manchester_decoder.counter[1] ;
 wire \user_manchester_decoder.counter[2] ;
 wire \user_manchester_decoder.counter[3] ;
 wire \user_manchester_decoder.counter[4] ;
 wire \user_manchester_decoder.counter[5] ;
 wire \user_manchester_decoder.last_in ;
 wire \user_manchester_decoder.middle ;
 wire \user_manchester_encoder.counter[0] ;
 wire \user_manchester_encoder.counter[1] ;
 wire \user_manchester_encoder.counter[2] ;
 wire \user_manchester_encoder.counter[3] ;
 wire \user_manchester_encoder.counter[4] ;
 wire \user_manchester_encoder.middle ;
 wire \user_protocol_counters.led_counter[0] ;
 wire \user_protocol_counters.led_counter[10] ;
 wire \user_protocol_counters.led_counter[11] ;
 wire \user_protocol_counters.led_counter[1] ;
 wire \user_protocol_counters.led_counter[2] ;
 wire \user_protocol_counters.led_counter[3] ;
 wire \user_protocol_counters.led_counter[4] ;
 wire \user_protocol_counters.led_counter[5] ;
 wire \user_protocol_counters.led_counter[6] ;
 wire \user_protocol_counters.led_counter[7] ;
 wire \user_protocol_counters.led_counter[8] ;
 wire \user_protocol_counters.led_counter[9] ;
 wire \user_protocol_parity.parity ;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;

 sg13g2_inv_1 _296_ (.Y(_068_),
    .A(net154));
 sg13g2_inv_1 _297_ (.Y(_069_),
    .A(uio_out[4]));
 sg13g2_inv_1 _298_ (.Y(_070_),
    .A(net169));
 sg13g2_inv_1 _299_ (.Y(_071_),
    .A(net162));
 sg13g2_inv_1 _300_ (.Y(_072_),
    .A(net168));
 sg13g2_inv_1 _301_ (.Y(_073_),
    .A(net92));
 sg13g2_inv_1 _302_ (.Y(_074_),
    .A(net207));
 sg13g2_inv_1 _303_ (.Y(_075_),
    .A(net108));
 sg13g2_inv_1 _304_ (.Y(_076_),
    .A(net143));
 sg13g2_inv_1 _305_ (.Y(_077_),
    .A(net189));
 sg13g2_inv_1 _306_ (.Y(_078_),
    .A(net156));
 sg13g2_inv_1 _307_ (.Y(_079_),
    .A(net218));
 sg13g2_inv_1 _308_ (.Y(_080_),
    .A(net145));
 sg13g2_inv_1 _309_ (.Y(_081_),
    .A(net148));
 sg13g2_inv_1 _310_ (.Y(_082_),
    .A(net164));
 sg13g2_inv_1 _311_ (.Y(_083_),
    .A(net200));
 sg13g2_inv_4 _312_ (.A(net26),
    .Y(_084_));
 sg13g2_inv_1 _313_ (.Y(_085_),
    .A(net30));
 sg13g2_inv_1 _314_ (.Y(_086_),
    .A(net2));
 sg13g2_and2_1 _315_ (.A(net125),
    .B(net27),
    .X(_000_));
 sg13g2_or2_1 _316_ (.X(_087_),
    .B(net27),
    .A(net192));
 sg13g2_nor2_2 _317_ (.A(net216),
    .B(net28),
    .Y(_088_));
 sg13g2_and3_1 _318_ (.X(_029_),
    .A(net25),
    .B(_087_),
    .C(_088_));
 sg13g2_a21o_1 _319_ (.A2(_088_),
    .A1(net27),
    .B1(_029_),
    .X(_001_));
 sg13g2_o21ai_1 _320_ (.B1(_088_),
    .Y(_089_),
    .A1(net192),
    .A2(net25));
 sg13g2_inv_1 _321_ (.Y(_002_),
    .A(net193));
 sg13g2_nand3_1 _322_ (.B(\protocol_counters_bits[1] ),
    .C(\protocol_counters_bits[0] ),
    .A(net125),
    .Y(_090_));
 sg13g2_and4_1 _323_ (.A(net125),
    .B(net151),
    .C(\protocol_counters_bits[1] ),
    .D(\protocol_counters_bits[0] ),
    .X(_091_));
 sg13g2_nand3_1 _324_ (.B(\protocol_counters_bits[3] ),
    .C(_091_),
    .A(\protocol_counters_bits[4] ),
    .Y(_092_));
 sg13g2_inv_1 _325_ (.Y(_093_),
    .A(_092_));
 sg13g2_and3_1 _326_ (.X(_094_),
    .A(net164),
    .B(\user_protocol_counters.led_counter[1] ),
    .C(\user_protocol_counters.led_counter[0] ));
 sg13g2_nand4_1 _327_ (.B(\user_protocol_counters.led_counter[2] ),
    .C(\user_protocol_counters.led_counter[1] ),
    .A(net117),
    .Y(_095_),
    .D(\user_protocol_counters.led_counter[0] ));
 sg13g2_nand2_2 _328_ (.Y(_096_),
    .A(net136),
    .B(net106));
 sg13g2_nand2_1 _329_ (.Y(_097_),
    .A(net110),
    .B(\user_protocol_counters.led_counter[6] ));
 sg13g2_or3_1 _330_ (.A(_095_),
    .B(_096_),
    .C(_097_),
    .X(_098_));
 sg13g2_nand3_1 _331_ (.B(\user_protocol_counters.led_counter[9] ),
    .C(net141),
    .A(net148),
    .Y(_099_));
 sg13g2_nand4_1 _332_ (.B(\user_protocol_counters.led_counter[10] ),
    .C(\user_protocol_counters.led_counter[9] ),
    .A(\user_protocol_counters.led_counter[11] ),
    .Y(_100_),
    .D(\user_protocol_counters.led_counter[8] ));
 sg13g2_nor4_2 _333_ (.A(_095_),
    .B(_096_),
    .C(_097_),
    .Y(_101_),
    .D(_100_));
 sg13g2_nor2_1 _334_ (.A(_092_),
    .B(_101_),
    .Y(_102_));
 sg13g2_nor3_1 _335_ (.A(_083_),
    .B(_092_),
    .C(_101_),
    .Y(_103_));
 sg13g2_o21ai_1 _336_ (.B1(net26),
    .Y(_104_),
    .A1(net200),
    .A2(_102_));
 sg13g2_nor2_1 _337_ (.A(_103_),
    .B(_104_),
    .Y(_003_));
 sg13g2_nand2_1 _338_ (.Y(_105_),
    .A(net202),
    .B(_103_));
 sg13g2_o21ai_1 _339_ (.B1(net27),
    .Y(_106_),
    .A1(net202),
    .A2(_103_));
 sg13g2_nor2b_1 _340_ (.A(_106_),
    .B_N(_105_),
    .Y(_004_));
 sg13g2_a221oi_1 _341_ (.B2(_082_),
    .C1(_084_),
    .B1(_105_),
    .A1(_094_),
    .Y(_005_),
    .A2(_102_));
 sg13g2_a21oi_1 _342_ (.A1(_094_),
    .A2(_102_),
    .Y(_107_),
    .B1(net117));
 sg13g2_nor3_2 _343_ (.A(_092_),
    .B(_095_),
    .C(_101_),
    .Y(_108_));
 sg13g2_nor3_1 _344_ (.A(_084_),
    .B(net118),
    .C(_108_),
    .Y(_006_));
 sg13g2_o21ai_1 _345_ (.B1(net27),
    .Y(_109_),
    .A1(net106),
    .A2(_108_));
 sg13g2_a21oi_1 _346_ (.A1(net106),
    .A2(_108_),
    .Y(_007_),
    .B1(_109_));
 sg13g2_a21oi_1 _347_ (.A1(net106),
    .A2(_108_),
    .Y(_110_),
    .B1(net136));
 sg13g2_nor4_2 _348_ (.A(_092_),
    .B(_095_),
    .C(_096_),
    .Y(_111_),
    .D(_101_));
 sg13g2_nor3_1 _349_ (.A(_084_),
    .B(net137),
    .C(_111_),
    .Y(_008_));
 sg13g2_o21ai_1 _350_ (.B1(net26),
    .Y(_112_),
    .A1(net134),
    .A2(_111_));
 sg13g2_a21oi_1 _351_ (.A1(net134),
    .A2(_111_),
    .Y(_009_),
    .B1(_112_));
 sg13g2_a21oi_1 _352_ (.A1(\user_protocol_counters.led_counter[6] ),
    .A2(_111_),
    .Y(_113_),
    .B1(net110));
 sg13g2_nor3_2 _353_ (.A(_092_),
    .B(_098_),
    .C(_101_),
    .Y(_114_));
 sg13g2_nor3_1 _354_ (.A(_084_),
    .B(net111),
    .C(_114_),
    .Y(_010_));
 sg13g2_o21ai_1 _355_ (.B1(net26),
    .Y(_115_),
    .A1(net141),
    .A2(_114_));
 sg13g2_a21oi_1 _356_ (.A1(net141),
    .A2(_114_),
    .Y(_011_),
    .B1(_115_));
 sg13g2_a21o_1 _357_ (.A2(_114_),
    .A1(net141),
    .B1(net215),
    .X(_116_));
 sg13g2_nand3_1 _358_ (.B(net141),
    .C(_114_),
    .A(net215),
    .Y(_117_));
 sg13g2_and3_1 _359_ (.X(_012_),
    .A(net26),
    .B(_116_),
    .C(_117_));
 sg13g2_nor4_1 _360_ (.A(_092_),
    .B(_098_),
    .C(_099_),
    .D(_101_),
    .Y(_118_));
 sg13g2_nand2b_1 _361_ (.Y(_119_),
    .B(net26),
    .A_N(_118_));
 sg13g2_a21oi_1 _362_ (.A1(_081_),
    .A2(_117_),
    .Y(_013_),
    .B1(_119_));
 sg13g2_o21ai_1 _363_ (.B1(net26),
    .Y(_120_),
    .A1(net174),
    .A2(_118_));
 sg13g2_inv_1 _364_ (.Y(_014_),
    .A(net175));
 sg13g2_a21oi_1 _365_ (.A1(_093_),
    .A2(_101_),
    .Y(_121_),
    .B1(net99));
 sg13g2_nor2_1 _366_ (.A(_084_),
    .B(net100),
    .Y(_015_));
 sg13g2_o21ai_1 _367_ (.B1(protocol_insync_out),
    .Y(_122_),
    .A1(net125),
    .A2(\protocol_counters_bits[0] ));
 sg13g2_a21oi_1 _368_ (.A1(net125),
    .A2(\protocol_counters_bits[0] ),
    .Y(_016_),
    .B1(_122_));
 sg13g2_a21oi_1 _369_ (.A1(net125),
    .A2(\protocol_counters_bits[0] ),
    .Y(_123_),
    .B1(\protocol_counters_bits[1] ));
 sg13g2_nand2_1 _370_ (.Y(_124_),
    .A(net128),
    .B(_090_));
 sg13g2_nor2_1 _371_ (.A(_123_),
    .B(net129),
    .Y(_017_));
 sg13g2_nor2b_1 _372_ (.A(net151),
    .B_N(_090_),
    .Y(_125_));
 sg13g2_nor3_1 _373_ (.A(_084_),
    .B(_091_),
    .C(net152),
    .Y(_018_));
 sg13g2_o21ai_1 _374_ (.B1(net26),
    .Y(_126_),
    .A1(net115),
    .A2(_091_));
 sg13g2_a21oi_1 _375_ (.A1(net115),
    .A2(_091_),
    .Y(_019_),
    .B1(_126_));
 sg13g2_a21oi_1 _376_ (.A1(net115),
    .A2(_091_),
    .Y(_127_),
    .B1(net131));
 sg13g2_nor3_1 _377_ (.A(_084_),
    .B(_093_),
    .C(net132),
    .Y(_020_));
 sg13g2_xnor2_1 _378_ (.Y(_128_),
    .A(net91),
    .B(net139));
 sg13g2_xor2_1 _379_ (.B(net139),
    .A(net91),
    .X(_129_));
 sg13g2_nand2_2 _380_ (.Y(_130_),
    .A(net32),
    .B(_128_));
 sg13g2_nor2_1 _381_ (.A(net92),
    .B(_130_),
    .Y(_021_));
 sg13g2_a21o_1 _382_ (.A2(net92),
    .A1(net168),
    .B1(_130_),
    .X(_131_));
 sg13g2_a21oi_1 _383_ (.A1(_072_),
    .A2(_073_),
    .Y(_022_),
    .B1(_131_));
 sg13g2_a21oi_1 _384_ (.A1(net168),
    .A2(net92),
    .Y(_132_),
    .B1(net162));
 sg13g2_and3_1 _385_ (.X(_133_),
    .A(net162),
    .B(net168),
    .C(net92));
 sg13g2_nor3_1 _386_ (.A(_130_),
    .B(_132_),
    .C(_133_),
    .Y(_023_));
 sg13g2_and2_1 _387_ (.A(net171),
    .B(_133_),
    .X(_134_));
 sg13g2_nor2_1 _388_ (.A(net171),
    .B(_133_),
    .Y(_135_));
 sg13g2_nor3_1 _389_ (.A(_130_),
    .B(_134_),
    .C(_135_),
    .Y(_024_));
 sg13g2_nand2_1 _390_ (.Y(_136_),
    .A(net194),
    .B(_134_));
 sg13g2_xnor2_1 _391_ (.Y(_137_),
    .A(net194),
    .B(_134_));
 sg13g2_nor2_1 _392_ (.A(_130_),
    .B(_137_),
    .Y(_025_));
 sg13g2_xor2_1 _393_ (.B(_136_),
    .A(net198),
    .X(_138_));
 sg13g2_nor2_1 _394_ (.A(_130_),
    .B(_138_),
    .Y(_026_));
 sg13g2_nor3_1 _395_ (.A(net151),
    .B(\protocol_counters_bits[1] ),
    .C(\protocol_counters_bits[0] ),
    .Y(_139_));
 sg13g2_nand3_1 _396_ (.B(protocol_counters_out_clk),
    .C(_139_),
    .A(net102),
    .Y(_140_));
 sg13g2_nor3_1 _397_ (.A(net131),
    .B(net115),
    .C(_140_),
    .Y(_141_));
 sg13g2_o21ai_1 _398_ (.B1(net27),
    .Y(_142_),
    .A1(net166),
    .A2(_141_));
 sg13g2_inv_1 _399_ (.Y(_027_),
    .A(net167));
 sg13g2_o21ai_1 _400_ (.B1(net27),
    .Y(_143_),
    .A1(net102),
    .A2(protocol_counters_out_clk));
 sg13g2_a21oi_1 _401_ (.A1(net102),
    .A2(protocol_counters_out_clk),
    .Y(_028_),
    .B1(_143_));
 sg13g2_nor2_1 _402_ (.A(\user_manchester_encoder.counter[1] ),
    .B(\user_manchester_encoder.counter[0] ),
    .Y(_144_));
 sg13g2_nor3_1 _403_ (.A(net185),
    .B(\user_manchester_encoder.counter[1] ),
    .C(\user_manchester_encoder.counter[0] ),
    .Y(_145_));
 sg13g2_nor4_1 _404_ (.A(net159),
    .B(\user_manchester_encoder.counter[2] ),
    .C(\user_manchester_encoder.counter[1] ),
    .D(\user_manchester_encoder.counter[0] ),
    .Y(_146_));
 sg13g2_nand2_1 _405_ (.Y(_147_),
    .A(_080_),
    .B(_146_));
 sg13g2_nor3_1 _406_ (.A(manchester_decoder_out_error),
    .B(net179),
    .C(net28),
    .Y(_148_));
 sg13g2_a22oi_1 _407_ (.Y(_030_),
    .B1(_147_),
    .B2(net180),
    .A2(_088_),
    .A1(net25));
 sg13g2_a21oi_2 _408_ (.B1(net25),
    .Y(_149_),
    .A2(_146_),
    .A1(_080_));
 sg13g2_inv_1 _409_ (.Y(_150_),
    .A(_149_));
 sg13g2_nand2_1 _410_ (.Y(_151_),
    .A(net203),
    .B(_149_));
 sg13g2_nand2b_1 _411_ (.Y(_152_),
    .B(net179),
    .A_N(manchester_decoder_out_clk));
 sg13g2_o21ai_1 _412_ (.B1(_088_),
    .Y(_153_),
    .A1(_147_),
    .A2(_152_));
 sg13g2_o21ai_1 _413_ (.B1(net204),
    .Y(_154_),
    .A1(net199),
    .A2(_149_));
 sg13g2_nor2_1 _414_ (.A(_153_),
    .B(net205),
    .Y(_031_));
 sg13g2_and2_1 _415_ (.A(\user_manchester_encoder.counter[1] ),
    .B(\user_manchester_encoder.counter[0] ),
    .X(_155_));
 sg13g2_nor2_1 _416_ (.A(net195),
    .B(_149_),
    .Y(_156_));
 sg13g2_nor3_1 _417_ (.A(net25),
    .B(_144_),
    .C(_155_),
    .Y(_157_));
 sg13g2_nor3_1 _418_ (.A(_153_),
    .B(net196),
    .C(_157_),
    .Y(_032_));
 sg13g2_nor2b_1 _419_ (.A(_144_),
    .B_N(net185),
    .Y(_158_));
 sg13g2_nor3_1 _420_ (.A(net25),
    .B(net186),
    .C(_158_),
    .Y(_159_));
 sg13g2_nor2_1 _421_ (.A(net169),
    .B(_149_),
    .Y(_160_));
 sg13g2_nor3_1 _422_ (.A(_153_),
    .B(net187),
    .C(_160_),
    .Y(_033_));
 sg13g2_nand2b_1 _423_ (.Y(_161_),
    .B(net159),
    .A_N(_145_));
 sg13g2_nor2_1 _424_ (.A(net25),
    .B(_146_),
    .Y(_162_));
 sg13g2_a221oi_1 _425_ (.B2(_162_),
    .C1(_153_),
    .B1(net160),
    .A1(_069_),
    .Y(_034_),
    .A2(_150_));
 sg13g2_a22oi_1 _426_ (.Y(_163_),
    .B1(_162_),
    .B2(net145),
    .A2(_150_),
    .A1(uio_out[5]));
 sg13g2_nor2_1 _427_ (.A(_153_),
    .B(net146),
    .Y(_035_));
 sg13g2_nand2b_1 _428_ (.Y(_164_),
    .B(_152_),
    .A_N(_149_));
 sg13g2_nor2_1 _429_ (.A(dout_data),
    .B(net25),
    .Y(_165_));
 sg13g2_a21oi_1 _430_ (.A1(manchester_decoder_out_clk),
    .A2(manchester_decoder_out_data),
    .Y(_166_),
    .B1(_165_));
 sg13g2_xnor2_1 _431_ (.Y(_167_),
    .A(_164_),
    .B(_166_));
 sg13g2_and2_1 _432_ (.A(_088_),
    .B(_167_),
    .X(_036_));
 sg13g2_and2_1 _433_ (.A(net210),
    .B(net177),
    .X(_168_));
 sg13g2_nand4_1 _434_ (.B(\all_input_selector.counter1[2] ),
    .C(\all_input_selector.counter1[1] ),
    .A(net120),
    .Y(_169_),
    .D(\all_input_selector.counter1[0] ));
 sg13g2_or2_1 _435_ (.X(_170_),
    .B(_169_),
    .A(_078_));
 sg13g2_nand3_1 _436_ (.B(\all_input_selector.counter1[6] ),
    .C(\all_input_selector.counter1[5] ),
    .A(net104),
    .Y(_171_));
 sg13g2_nor3_2 _437_ (.A(_078_),
    .B(_169_),
    .C(_171_),
    .Y(_172_));
 sg13g2_nand2b_2 _438_ (.Y(_173_),
    .B(net2),
    .A_N(\all_input_selector.last_in1 ));
 sg13g2_o21ai_1 _439_ (.B1(_079_),
    .Y(_174_),
    .A1(_172_),
    .A2(_173_));
 sg13g2_nor3_2 _440_ (.A(_079_),
    .B(_172_),
    .C(_173_),
    .Y(_175_));
 sg13g2_nand2_1 _441_ (.Y(_176_),
    .A(net31),
    .B(net219));
 sg13g2_nor2_1 _442_ (.A(_175_),
    .B(_176_),
    .Y(_037_));
 sg13g2_xnor2_1 _443_ (.Y(_177_),
    .A(net177),
    .B(_175_));
 sg13g2_nor2_1 _444_ (.A(net28),
    .B(net178),
    .Y(_038_));
 sg13g2_a21o_1 _445_ (.A2(_175_),
    .A1(net177),
    .B1(net210),
    .X(_178_));
 sg13g2_nand2_1 _446_ (.Y(_179_),
    .A(_168_),
    .B(_175_));
 sg13g2_and3_1 _447_ (.X(_039_),
    .A(net31),
    .B(net211),
    .C(_179_));
 sg13g2_a21oi_1 _448_ (.A1(_168_),
    .A2(_175_),
    .Y(_180_),
    .B1(net120));
 sg13g2_nor3_1 _449_ (.A(_169_),
    .B(_172_),
    .C(_173_),
    .Y(_181_));
 sg13g2_nor3_1 _450_ (.A(net28),
    .B(net121),
    .C(_181_),
    .Y(_040_));
 sg13g2_nor2_1 _451_ (.A(net156),
    .B(_181_),
    .Y(_182_));
 sg13g2_nor3_1 _452_ (.A(_170_),
    .B(_172_),
    .C(_173_),
    .Y(_183_));
 sg13g2_nor3_1 _453_ (.A(net28),
    .B(net157),
    .C(_183_),
    .Y(_041_));
 sg13g2_nor4_2 _454_ (.A(_077_),
    .B(_170_),
    .C(_172_),
    .Y(_184_),
    .D(_173_));
 sg13g2_o21ai_1 _455_ (.B1(net30),
    .Y(_185_),
    .A1(net189),
    .A2(_183_));
 sg13g2_nor2_1 _456_ (.A(_184_),
    .B(net190),
    .Y(_042_));
 sg13g2_o21ai_1 _457_ (.B1(net30),
    .Y(_186_),
    .A1(net123),
    .A2(_184_));
 sg13g2_a21oi_1 _458_ (.A1(net123),
    .A2(_184_),
    .Y(_043_),
    .B1(_186_));
 sg13g2_a21oi_1 _459_ (.A1(\all_input_selector.counter1[6] ),
    .A2(_184_),
    .Y(_187_),
    .B1(net104));
 sg13g2_nor2_1 _460_ (.A(net29),
    .B(net105),
    .Y(_044_));
 sg13g2_nand3_1 _461_ (.B(\all_input_selector.counter0[1] ),
    .C(net113),
    .A(net143),
    .Y(_188_));
 sg13g2_and4_1 _462_ (.A(net97),
    .B(net143),
    .C(\all_input_selector.counter0[1] ),
    .D(net113),
    .X(_189_));
 sg13g2_inv_1 _463_ (.Y(_190_),
    .A(_189_));
 sg13g2_and3_2 _464_ (.X(_191_),
    .A(net108),
    .B(net182),
    .C(_189_));
 sg13g2_nand2b_2 _465_ (.Y(_192_),
    .B(net1),
    .A_N(\all_input_selector.last_in0 ));
 sg13g2_nor3_2 _466_ (.A(_172_),
    .B(_191_),
    .C(_192_),
    .Y(_193_));
 sg13g2_o21ai_1 _467_ (.B1(net30),
    .Y(_194_),
    .A1(net113),
    .A2(_193_));
 sg13g2_a21oi_1 _468_ (.A1(net113),
    .A2(_193_),
    .Y(_045_),
    .B1(_194_));
 sg13g2_a21o_1 _469_ (.A2(_193_),
    .A1(net113),
    .B1(net213),
    .X(_195_));
 sg13g2_nand3_1 _470_ (.B(net113),
    .C(_193_),
    .A(net213),
    .Y(_196_));
 sg13g2_and3_1 _471_ (.X(_046_),
    .A(net30),
    .B(net214),
    .C(_196_));
 sg13g2_nor4_1 _472_ (.A(_172_),
    .B(_188_),
    .C(_191_),
    .D(_192_),
    .Y(_197_));
 sg13g2_nand2b_1 _473_ (.Y(_198_),
    .B(net30),
    .A_N(_197_));
 sg13g2_a21oi_1 _474_ (.A1(_076_),
    .A2(_196_),
    .Y(_047_),
    .B1(_198_));
 sg13g2_o21ai_1 _475_ (.B1(net30),
    .Y(_199_),
    .A1(net97),
    .A2(_197_));
 sg13g2_a21oi_1 _476_ (.A1(net97),
    .A2(_197_),
    .Y(_048_),
    .B1(_199_));
 sg13g2_nor3_1 _477_ (.A(_172_),
    .B(_190_),
    .C(_192_),
    .Y(_200_));
 sg13g2_o21ai_1 _478_ (.B1(net31),
    .Y(_201_),
    .A1(net182),
    .A2(_200_));
 sg13g2_nand3_1 _479_ (.B(_189_),
    .C(_193_),
    .A(net182),
    .Y(_202_));
 sg13g2_nor2b_1 _480_ (.A(net183),
    .B_N(_202_),
    .Y(_049_));
 sg13g2_a21oi_1 _481_ (.A1(_075_),
    .A2(_202_),
    .Y(_050_),
    .B1(net29));
 sg13g2_xnor2_1 _482_ (.Y(_203_),
    .A(net3),
    .B(_191_));
 sg13g2_nor2_1 _483_ (.A(net1),
    .B(_203_),
    .Y(_204_));
 sg13g2_nor2_1 _484_ (.A(net29),
    .B(_203_),
    .Y(_052_));
 sg13g2_nor2_1 _485_ (.A(net29),
    .B(_086_),
    .Y(_056_));
 sg13g2_a21oi_1 _486_ (.A1(_086_),
    .A2(_203_),
    .Y(_205_),
    .B1(net29));
 sg13g2_nor2b_1 _487_ (.A(_204_),
    .B_N(_205_),
    .Y(_051_));
 sg13g2_and2_1 _488_ (.A(net31),
    .B(net1),
    .X(_053_));
 sg13g2_and2_1 _489_ (.A(net30),
    .B(net127),
    .X(_054_));
 sg13g2_a21oi_1 _490_ (.A1(\all_low_pass_filter.last0 ),
    .A2(\all_input_selector.out ),
    .Y(_206_),
    .B1(net94));
 sg13g2_and2_1 _491_ (.A(net32),
    .B(net150),
    .X(_067_));
 sg13g2_nor2_1 _492_ (.A(_054_),
    .B(_067_),
    .Y(_207_));
 sg13g2_nor2_1 _493_ (.A(net95),
    .B(_207_),
    .Y(_055_));
 sg13g2_or3_1 _494_ (.A(\user_manchester_decoder.counter[3] ),
    .B(\user_manchester_decoder.counter[2] ),
    .C(\user_manchester_decoder.counter[1] ),
    .X(_208_));
 sg13g2_a21o_2 _495_ (.A2(_208_),
    .A1(net194),
    .B1(net198),
    .X(_209_));
 sg13g2_or2_1 _496_ (.X(_210_),
    .B(\user_manchester_decoder.counter[3] ),
    .A(\user_manchester_decoder.counter[4] ));
 sg13g2_o21ai_1 _497_ (.B1(net222),
    .Y(_211_),
    .A1(\user_manchester_decoder.counter[2] ),
    .A2(_210_));
 sg13g2_and3_1 _498_ (.X(_212_),
    .A(_129_),
    .B(_209_),
    .C(_211_));
 sg13g2_nand3_1 _499_ (.B(_209_),
    .C(_211_),
    .A(_129_),
    .Y(_213_));
 sg13g2_a21oi_1 _500_ (.A1(net162),
    .A2(net168),
    .Y(_214_),
    .B1(_210_));
 sg13g2_or3_1 _501_ (.A(net216),
    .B(_209_),
    .C(_214_),
    .X(_215_));
 sg13g2_nor4_1 _502_ (.A(net216),
    .B(_128_),
    .C(_209_),
    .D(_214_),
    .Y(_216_));
 sg13g2_or2_1 _503_ (.X(_217_),
    .B(_216_),
    .A(net24));
 sg13g2_nor3_1 _504_ (.A(net207),
    .B(net24),
    .C(_216_),
    .Y(_218_));
 sg13g2_nor4_1 _505_ (.A(_074_),
    .B(_128_),
    .C(_209_),
    .D(_215_),
    .Y(_219_));
 sg13g2_nor3_1 _506_ (.A(net28),
    .B(net208),
    .C(_219_),
    .Y(_057_));
 sg13g2_a21o_1 _507_ (.A2(net223),
    .A1(_209_),
    .B1(_074_),
    .X(_220_));
 sg13g2_and3_1 _508_ (.X(_058_),
    .A(net32),
    .B(_217_),
    .C(_220_));
 sg13g2_o21ai_1 _509_ (.B1(net32),
    .Y(_221_),
    .A1(net176),
    .A2(net23));
 sg13g2_a21oi_1 _510_ (.A1(_073_),
    .A2(net23),
    .Y(_059_),
    .B1(_221_));
 sg13g2_o21ai_1 _511_ (.B1(net32),
    .Y(_222_),
    .A1(net199),
    .A2(net23));
 sg13g2_a21oi_1 _512_ (.A1(_072_),
    .A2(net23),
    .Y(_060_),
    .B1(_222_));
 sg13g2_o21ai_1 _513_ (.B1(net32),
    .Y(_223_),
    .A1(uio_out[2]),
    .A2(net23));
 sg13g2_a21oi_1 _514_ (.A1(_071_),
    .A2(net24),
    .Y(_061_),
    .B1(_223_));
 sg13g2_a21oi_1 _515_ (.A1(\user_manchester_decoder.counter[3] ),
    .A2(net23),
    .Y(_224_),
    .B1(net28));
 sg13g2_o21ai_1 _516_ (.B1(_224_),
    .Y(_062_),
    .A1(_070_),
    .A2(net23));
 sg13g2_a21o_1 _517_ (.A2(net23),
    .A1(\user_manchester_decoder.counter[4] ),
    .B1(net28),
    .X(_225_));
 sg13g2_a21o_1 _518_ (.A2(_213_),
    .A1(net172),
    .B1(_225_),
    .X(_063_));
 sg13g2_a21oi_1 _519_ (.A1(_068_),
    .A2(_213_),
    .Y(_064_),
    .B1(_225_));
 sg13g2_o21ai_1 _520_ (.B1(_215_),
    .Y(_226_),
    .A1(net216),
    .A2(_129_));
 sg13g2_o21ai_1 _521_ (.B1(net32),
    .Y(_065_),
    .A1(net24),
    .A2(_226_));
 sg13g2_and4_1 _522_ (.A(net139),
    .B(net32),
    .C(_217_),
    .D(_220_),
    .X(_066_));
 sg13g2_dfrbpq_1 _523_ (.RESET_B(net78),
    .D(_000_),
    .Q(protocol_counters_out_clk),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _524_ (.RESET_B(net33),
    .D(_001_),
    .Q(protocol_insync_out),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _525_ (.RESET_B(net21),
    .D(_002_),
    .Q(dout_enable),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _526_ (.RESET_B(net19),
    .D(net201),
    .Q(\user_protocol_counters.led_counter[0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _527_ (.RESET_B(net17),
    .D(_004_),
    .Q(\user_protocol_counters.led_counter[1] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _528_ (.RESET_B(net15),
    .D(net165),
    .Q(\user_protocol_counters.led_counter[2] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _529_ (.RESET_B(net13),
    .D(net119),
    .Q(\user_protocol_counters.led_counter[3] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _530_ (.RESET_B(net11),
    .D(net107),
    .Q(\user_protocol_counters.led_counter[4] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _531_ (.RESET_B(net88),
    .D(net138),
    .Q(\user_protocol_counters.led_counter[5] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _532_ (.RESET_B(net86),
    .D(net135),
    .Q(\user_protocol_counters.led_counter[6] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _533_ (.RESET_B(net84),
    .D(net112),
    .Q(\user_protocol_counters.led_counter[7] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _534_ (.RESET_B(net82),
    .D(net142),
    .Q(\user_protocol_counters.led_counter[8] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _535_ (.RESET_B(net80),
    .D(_012_),
    .Q(\user_protocol_counters.led_counter[9] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _536_ (.RESET_B(net77),
    .D(net149),
    .Q(\user_protocol_counters.led_counter[10] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _537_ (.RESET_B(net75),
    .D(_014_),
    .Q(\user_protocol_counters.led_counter[11] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _538_ (.RESET_B(net73),
    .D(net101),
    .Q(protocol_counters_test_mode_out),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _539_ (.RESET_B(net71),
    .D(net126),
    .Q(\protocol_counters_bits[0] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _540_ (.RESET_B(net69),
    .D(net130),
    .Q(\protocol_counters_bits[1] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _541_ (.RESET_B(net67),
    .D(net153),
    .Q(\protocol_counters_bits[2] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _542_ (.RESET_B(net65),
    .D(net116),
    .Q(\protocol_counters_bits[3] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _543_ (.RESET_B(net63),
    .D(net133),
    .Q(\protocol_counters_bits[4] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _544_ (.RESET_B(net61),
    .D(net93),
    .Q(\user_manchester_decoder.counter[0] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _545_ (.RESET_B(net60),
    .D(_022_),
    .Q(\user_manchester_decoder.counter[1] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _546_ (.RESET_B(net59),
    .D(_023_),
    .Q(\user_manchester_decoder.counter[2] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _547_ (.RESET_B(net58),
    .D(_024_),
    .Q(\user_manchester_decoder.counter[3] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _548_ (.RESET_B(net57),
    .D(_025_),
    .Q(\user_manchester_decoder.counter[4] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _549_ (.RESET_B(net56),
    .D(_026_),
    .Q(\user_manchester_decoder.counter[5] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _550_ (.RESET_B(net55),
    .D(_027_),
    .Q(protocol_parity_error),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _551_ (.RESET_B(net53),
    .D(net103),
    .Q(\user_protocol_parity.parity ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _552_ (.RESET_B(net51),
    .D(_029_),
    .Q(protocol_insync_out_clk),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _553_ (.RESET_B(net50),
    .D(net181),
    .Q(\user_manchester_encoder.middle ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _554_ (.RESET_B(net48),
    .D(net206),
    .Q(\user_manchester_encoder.counter[0] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _555_ (.RESET_B(net46),
    .D(net197),
    .Q(\user_manchester_encoder.counter[1] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _556_ (.RESET_B(net44),
    .D(net188),
    .Q(\user_manchester_encoder.counter[2] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _557_ (.RESET_B(net42),
    .D(net161),
    .Q(\user_manchester_encoder.counter[3] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _558_ (.RESET_B(net40),
    .D(net147),
    .Q(\user_manchester_encoder.counter[4] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _559_ (.RESET_B(net38),
    .D(net217),
    .Q(dout_data),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_1 _560_ (.RESET_B(net36),
    .D(net220),
    .Q(\all_input_selector.counter1[0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _561_ (.RESET_B(net34),
    .D(_038_),
    .Q(\all_input_selector.counter1[1] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _562_ (.RESET_B(net20),
    .D(net212),
    .Q(\all_input_selector.counter1[2] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _563_ (.RESET_B(net16),
    .D(net122),
    .Q(\all_input_selector.counter1[3] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _564_ (.RESET_B(net12),
    .D(net158),
    .Q(\all_input_selector.counter1[4] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _565_ (.RESET_B(net87),
    .D(net191),
    .Q(\all_input_selector.counter1[5] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _566_ (.RESET_B(net83),
    .D(net124),
    .Q(\all_input_selector.counter1[6] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _567_ (.RESET_B(net79),
    .D(_044_),
    .Q(\all_input_selector.counter1[7] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _568_ (.RESET_B(net74),
    .D(net114),
    .Q(\all_input_selector.counter0[0] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _569_ (.RESET_B(net70),
    .D(_046_),
    .Q(\all_input_selector.counter0[1] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _570_ (.RESET_B(net66),
    .D(net144),
    .Q(\all_input_selector.counter0[2] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _571_ (.RESET_B(net62),
    .D(net98),
    .Q(\all_input_selector.counter0[3] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _572_ (.RESET_B(net52),
    .D(net184),
    .Q(\all_input_selector.counter0[4] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _573_ (.RESET_B(net47),
    .D(net109),
    .Q(\all_input_selector.counter0[5] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _574_ (.RESET_B(net43),
    .D(_051_),
    .Q(\all_input_selector.out ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _575_ (.RESET_B(net41),
    .D(_052_),
    .Q(\all_input_selector.in0selected ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _576_ (.RESET_B(net39),
    .D(_053_),
    .Q(\all_input_selector.last_in0 ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _577_ (.RESET_B(net37),
    .D(_054_),
    .Q(\all_low_pass_filter.last1 ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _578_ (.RESET_B(net35),
    .D(net96),
    .Q(\all_low_pass_filter.out ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _579_ (.RESET_B(net49),
    .D(_056_),
    .Q(\all_input_selector.last_in1 ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _580_ (.RESET_B(net22),
    .D(net91),
    .Q(\user_manchester_decoder.last_in ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _581_ (.RESET_B(net18),
    .D(net209),
    .Q(\user_manchester_decoder.middle ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _582_ (.RESET_B(net89),
    .D(_058_),
    .Q(manchester_decoder_out_clk),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _583_ (.RESET_B(net85),
    .D(_059_),
    .Q(uio_out[0]),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _584_ (.RESET_B(net76),
    .D(_060_),
    .Q(uio_out[1]),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _585_ (.RESET_B(net68),
    .D(net163),
    .Q(uio_out[2]),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _586_ (.RESET_B(net54),
    .D(net170),
    .Q(uio_out[3]),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _587_ (.RESET_B(net45),
    .D(net173),
    .Q(uio_out[4]),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _588_ (.RESET_B(net81),
    .D(net155),
    .Q(uio_out[5]),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _589_ (.RESET_B(net64),
    .D(_065_),
    .Q(manchester_decoder_out_error),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _590_ (.RESET_B(net14),
    .D(net140),
    .Q(manchester_decoder_out_data),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_1 _591_ (.RESET_B(net72),
    .D(_067_),
    .Q(\all_low_pass_filter.last0 ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_tiehi _564__12 (.L_HI(net12));
 sg13g2_tiehi _529__13 (.L_HI(net13));
 sg13g2_tiehi _590__14 (.L_HI(net14));
 sg13g2_tiehi _528__15 (.L_HI(net15));
 sg13g2_tiehi _563__16 (.L_HI(net16));
 sg13g2_tiehi _527__17 (.L_HI(net17));
 sg13g2_tiehi _581__18 (.L_HI(net18));
 sg13g2_tiehi _526__19 (.L_HI(net19));
 sg13g2_tiehi _562__20 (.L_HI(net20));
 sg13g2_tiehi _525__21 (.L_HI(net21));
 sg13g2_tiehi _580__22 (.L_HI(net22));
 sg13g2_tiehi _524__23 (.L_HI(net33));
 sg13g2_tiehi _561__24 (.L_HI(net34));
 sg13g2_tiehi _578__25 (.L_HI(net35));
 sg13g2_tiehi _560__26 (.L_HI(net36));
 sg13g2_tiehi _577__27 (.L_HI(net37));
 sg13g2_tiehi _559__28 (.L_HI(net38));
 sg13g2_tiehi _576__29 (.L_HI(net39));
 sg13g2_tiehi _558__30 (.L_HI(net40));
 sg13g2_tiehi _575__31 (.L_HI(net41));
 sg13g2_tiehi _557__32 (.L_HI(net42));
 sg13g2_tiehi _574__33 (.L_HI(net43));
 sg13g2_tiehi _556__34 (.L_HI(net44));
 sg13g2_tiehi _587__35 (.L_HI(net45));
 sg13g2_tiehi _555__36 (.L_HI(net46));
 sg13g2_tiehi _573__37 (.L_HI(net47));
 sg13g2_tiehi _554__38 (.L_HI(net48));
 sg13g2_tiehi _579__39 (.L_HI(net49));
 sg13g2_tiehi _553__40 (.L_HI(net50));
 sg13g2_tiehi _552__41 (.L_HI(net51));
 sg13g2_tiehi _572__42 (.L_HI(net52));
 sg13g2_tiehi _551__43 (.L_HI(net53));
 sg13g2_tiehi _586__44 (.L_HI(net54));
 sg13g2_tiehi _550__45 (.L_HI(net55));
 sg13g2_tiehi _549__46 (.L_HI(net56));
 sg13g2_tiehi _548__47 (.L_HI(net57));
 sg13g2_tiehi _547__48 (.L_HI(net58));
 sg13g2_tiehi _546__49 (.L_HI(net59));
 sg13g2_tiehi _545__50 (.L_HI(net60));
 sg13g2_tiehi _544__51 (.L_HI(net61));
 sg13g2_tiehi _571__52 (.L_HI(net62));
 sg13g2_tiehi _543__53 (.L_HI(net63));
 sg13g2_tiehi _589__54 (.L_HI(net64));
 sg13g2_tiehi _542__55 (.L_HI(net65));
 sg13g2_tiehi _570__56 (.L_HI(net66));
 sg13g2_tiehi _541__57 (.L_HI(net67));
 sg13g2_tiehi _585__58 (.L_HI(net68));
 sg13g2_tiehi _540__59 (.L_HI(net69));
 sg13g2_tiehi _569__60 (.L_HI(net70));
 sg13g2_tiehi _539__61 (.L_HI(net71));
 sg13g2_tiehi _591__62 (.L_HI(net72));
 sg13g2_tiehi _538__63 (.L_HI(net73));
 sg13g2_tiehi _568__64 (.L_HI(net74));
 sg13g2_tiehi _537__65 (.L_HI(net75));
 sg13g2_tiehi _584__66 (.L_HI(net76));
 sg13g2_tiehi _536__67 (.L_HI(net77));
 sg13g2_tiehi _523__68 (.L_HI(net78));
 sg13g2_tiehi _567__69 (.L_HI(net79));
 sg13g2_tiehi _535__70 (.L_HI(net80));
 sg13g2_tiehi _588__71 (.L_HI(net81));
 sg13g2_tiehi _534__72 (.L_HI(net82));
 sg13g2_tiehi _566__73 (.L_HI(net83));
 sg13g2_tiehi _533__74 (.L_HI(net84));
 sg13g2_tiehi _583__75 (.L_HI(net85));
 sg13g2_tiehi _532__76 (.L_HI(net86));
 sg13g2_tiehi _565__77 (.L_HI(net87));
 sg13g2_tiehi _531__78 (.L_HI(net88));
 sg13g2_tiehi _582__79 (.L_HI(net89));
 sg13g2_tiehi tt_um_hoene_smart_led_digital_80 (.L_HI(net90));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_hoene_smart_led_digital_5 (.L_LO(net5));
 sg13g2_tielo tt_um_hoene_smart_led_digital_6 (.L_LO(net6));
 sg13g2_tielo tt_um_hoene_smart_led_digital_7 (.L_LO(net7));
 sg13g2_tielo tt_um_hoene_smart_led_digital_8 (.L_LO(net8));
 sg13g2_tielo tt_um_hoene_smart_led_digital_9 (.L_LO(net9));
 sg13g2_tielo tt_um_hoene_smart_led_digital_10 (.L_LO(net10));
 sg13g2_tiehi _530__11 (.L_HI(net11));
 sg13g2_buf_1 _669_ (.A(dout_enable),
    .X(uio_oe[7]));
 sg13g2_buf_1 _670_ (.A(dout_data),
    .X(uio_out[7]));
 sg13g2_buf_1 _671_ (.A(\all_input_selector.out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _672_ (.A(\all_input_selector.in0selected ),
    .X(uo_out[1]));
 sg13g2_buf_1 _673_ (.A(\all_low_pass_filter.out ),
    .X(uo_out[2]));
 sg13g2_buf_1 _674_ (.A(manchester_decoder_out_data),
    .X(uo_out[3]));
 sg13g2_buf_1 _675_ (.A(manchester_decoder_out_clk),
    .X(uo_out[4]));
 sg13g2_buf_1 _676_ (.A(manchester_decoder_out_error),
    .X(uo_out[5]));
 sg13g2_buf_1 _677_ (.A(protocol_counters_test_mode_out),
    .X(uo_out[6]));
 sg13g2_buf_1 _678_ (.A(protocol_parity_error),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout23 (.A(net24),
    .X(net23));
 sg13g2_buf_1 fanout24 (.A(_212_),
    .X(net24));
 sg13g2_buf_8 fanout25 (.A(net221),
    .X(net25));
 sg13g2_buf_8 fanout26 (.A(net27),
    .X(net26));
 sg13g2_buf_8 fanout27 (.A(net128),
    .X(net27));
 sg13g2_buf_8 fanout28 (.A(_085_),
    .X(net28));
 sg13g2_buf_1 fanout29 (.A(_085_),
    .X(net29));
 sg13g2_buf_8 fanout30 (.A(rst_n),
    .X(net30));
 sg13g2_buf_1 fanout31 (.A(rst_n),
    .X(net31));
 sg13g2_buf_8 fanout32 (.A(rst_n),
    .X(net32));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_tielo tt_um_hoene_smart_led_digital_4 (.L_LO(net4));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\all_low_pass_filter.out ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold2 (.A(\user_manchester_decoder.counter[0] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold3 (.A(_021_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold4 (.A(\all_low_pass_filter.last1 ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold5 (.A(_206_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold6 (.A(_055_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold7 (.A(\all_input_selector.counter0[3] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold8 (.A(_048_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold9 (.A(protocol_counters_test_mode_out),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold10 (.A(_121_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold11 (.A(_015_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold12 (.A(\user_protocol_parity.parity ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold13 (.A(_028_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold14 (.A(\all_input_selector.counter1[7] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold15 (.A(_187_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold16 (.A(\user_protocol_counters.led_counter[4] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold17 (.A(_007_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold18 (.A(\all_input_selector.counter0[5] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold19 (.A(_050_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold20 (.A(\user_protocol_counters.led_counter[7] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold21 (.A(_113_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold22 (.A(_010_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold23 (.A(\all_input_selector.counter0[0] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold24 (.A(_045_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold25 (.A(\protocol_counters_bits[3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold26 (.A(_019_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold27 (.A(\user_protocol_counters.led_counter[3] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold28 (.A(_107_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold29 (.A(_006_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold30 (.A(\all_input_selector.counter1[3] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold31 (.A(_180_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold32 (.A(_040_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold33 (.A(\all_input_selector.counter1[6] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold34 (.A(_043_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold35 (.A(protocol_insync_out_clk),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold36 (.A(_016_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold37 (.A(\all_low_pass_filter.last0 ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold38 (.A(protocol_insync_out),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold39 (.A(_124_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold40 (.A(_017_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold41 (.A(\protocol_counters_bits[4] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold42 (.A(_127_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold43 (.A(_020_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold44 (.A(\user_protocol_counters.led_counter[6] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold45 (.A(_009_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold46 (.A(\user_protocol_counters.led_counter[5] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold47 (.A(_110_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold48 (.A(_008_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold49 (.A(\user_manchester_decoder.last_in ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold50 (.A(_066_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold51 (.A(\user_protocol_counters.led_counter[8] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold52 (.A(_011_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold53 (.A(\all_input_selector.counter0[2] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold54 (.A(_047_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold55 (.A(\user_manchester_encoder.counter[4] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold56 (.A(_163_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold57 (.A(_035_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold58 (.A(\user_protocol_counters.led_counter[10] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold59 (.A(_013_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold60 (.A(\all_input_selector.out ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold61 (.A(\protocol_counters_bits[2] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold62 (.A(_125_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold63 (.A(_018_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold64 (.A(uio_out[5]),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold65 (.A(_064_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold66 (.A(\all_input_selector.counter1[4] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold67 (.A(_182_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold68 (.A(_041_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold69 (.A(\user_manchester_encoder.counter[3] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold70 (.A(_161_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold71 (.A(_034_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold72 (.A(\user_manchester_decoder.counter[2] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold73 (.A(_061_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold74 (.A(\user_protocol_counters.led_counter[2] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold75 (.A(_005_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold76 (.A(protocol_parity_error),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold77 (.A(_142_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold78 (.A(\user_manchester_decoder.counter[1] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold79 (.A(uio_out[3]),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold80 (.A(_062_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold81 (.A(\user_manchester_decoder.counter[3] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold82 (.A(uio_out[4]),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold83 (.A(_063_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold84 (.A(\user_protocol_counters.led_counter[11] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold85 (.A(_120_),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold86 (.A(uio_out[0]),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold87 (.A(\all_input_selector.counter1[1] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold88 (.A(_177_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold89 (.A(\user_manchester_encoder.middle ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold90 (.A(_148_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold91 (.A(_030_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold92 (.A(\all_input_selector.counter0[4] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold93 (.A(_201_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold94 (.A(_049_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold95 (.A(\user_manchester_encoder.counter[2] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold96 (.A(_145_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold97 (.A(_159_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold98 (.A(_033_),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold99 (.A(\all_input_selector.counter1[5] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold100 (.A(_185_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold101 (.A(_042_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold102 (.A(dout_enable),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold103 (.A(_089_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold104 (.A(\user_manchester_decoder.counter[4] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold105 (.A(uio_out[2]),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold106 (.A(_156_),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold107 (.A(_032_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold108 (.A(\user_manchester_decoder.counter[5] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold109 (.A(uio_out[1]),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold110 (.A(\user_protocol_counters.led_counter[0] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold111 (.A(_003_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold112 (.A(\user_protocol_counters.led_counter[1] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold113 (.A(\user_manchester_encoder.counter[0] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold114 (.A(_151_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold115 (.A(_154_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold116 (.A(_031_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold117 (.A(\user_manchester_decoder.middle ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold118 (.A(_218_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold119 (.A(_057_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold120 (.A(\all_input_selector.counter1[2] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold121 (.A(_178_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold122 (.A(_039_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold123 (.A(\all_input_selector.counter0[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold124 (.A(_195_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold125 (.A(\user_protocol_counters.led_counter[9] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold126 (.A(manchester_decoder_out_error),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold127 (.A(_036_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold128 (.A(\all_input_selector.counter1[0] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold129 (.A(_174_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold130 (.A(_037_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold131 (.A(manchester_decoder_out_clk),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold132 (.A(\user_manchester_decoder.counter[5] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold133 (.A(_211_),
    .X(net223));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_fill_1 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_47 ();
 sg13g2_decap_8 FILLER_14_54 ();
 sg13g2_decap_8 FILLER_14_61 ();
 sg13g2_decap_8 FILLER_14_68 ();
 sg13g2_decap_8 FILLER_14_75 ();
 sg13g2_decap_8 FILLER_14_82 ();
 sg13g2_decap_8 FILLER_14_89 ();
 sg13g2_decap_8 FILLER_14_96 ();
 sg13g2_decap_8 FILLER_14_103 ();
 sg13g2_decap_8 FILLER_14_110 ();
 sg13g2_decap_8 FILLER_14_117 ();
 sg13g2_decap_8 FILLER_14_124 ();
 sg13g2_decap_8 FILLER_14_131 ();
 sg13g2_decap_8 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_152 ();
 sg13g2_decap_8 FILLER_14_159 ();
 sg13g2_decap_8 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_173 ();
 sg13g2_decap_8 FILLER_14_180 ();
 sg13g2_decap_8 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_8 FILLER_14_215 ();
 sg13g2_decap_8 FILLER_14_222 ();
 sg13g2_decap_8 FILLER_14_229 ();
 sg13g2_decap_8 FILLER_14_236 ();
 sg13g2_decap_8 FILLER_14_243 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_decap_8 FILLER_14_257 ();
 sg13g2_decap_8 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_271 ();
 sg13g2_decap_8 FILLER_14_278 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_64 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_8 FILLER_15_78 ();
 sg13g2_decap_8 FILLER_15_85 ();
 sg13g2_decap_8 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_decap_8 FILLER_15_113 ();
 sg13g2_decap_8 FILLER_15_120 ();
 sg13g2_decap_8 FILLER_15_127 ();
 sg13g2_decap_8 FILLER_15_134 ();
 sg13g2_decap_8 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_148 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_169 ();
 sg13g2_decap_8 FILLER_15_176 ();
 sg13g2_decap_8 FILLER_15_183 ();
 sg13g2_decap_8 FILLER_15_190 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_260 ();
 sg13g2_decap_8 FILLER_15_267 ();
 sg13g2_decap_8 FILLER_15_274 ();
 sg13g2_decap_8 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_288 ();
 sg13g2_decap_8 FILLER_15_295 ();
 sg13g2_decap_8 FILLER_15_302 ();
 sg13g2_decap_8 FILLER_15_309 ();
 sg13g2_decap_8 FILLER_15_316 ();
 sg13g2_decap_8 FILLER_15_323 ();
 sg13g2_decap_8 FILLER_15_330 ();
 sg13g2_decap_8 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_344 ();
 sg13g2_decap_8 FILLER_15_351 ();
 sg13g2_decap_8 FILLER_15_358 ();
 sg13g2_decap_8 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_379 ();
 sg13g2_decap_8 FILLER_15_386 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_4 ();
 sg13g2_fill_2 FILLER_16_33 ();
 sg13g2_fill_1 FILLER_16_35 ();
 sg13g2_fill_2 FILLER_16_41 ();
 sg13g2_fill_2 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_65 ();
 sg13g2_fill_1 FILLER_16_72 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_40 ();
 sg13g2_fill_2 FILLER_17_50 ();
 sg13g2_decap_8 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_8 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_decap_8 FILLER_17_137 ();
 sg13g2_decap_8 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_151 ();
 sg13g2_decap_8 FILLER_17_158 ();
 sg13g2_decap_8 FILLER_17_165 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_fill_2 FILLER_18_35 ();
 sg13g2_decap_4 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_66 ();
 sg13g2_decap_8 FILLER_18_89 ();
 sg13g2_fill_1 FILLER_18_96 ();
 sg13g2_decap_4 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_118 ();
 sg13g2_decap_8 FILLER_18_125 ();
 sg13g2_decap_8 FILLER_18_132 ();
 sg13g2_decap_8 FILLER_18_139 ();
 sg13g2_decap_8 FILLER_18_146 ();
 sg13g2_decap_8 FILLER_18_153 ();
 sg13g2_decap_8 FILLER_18_160 ();
 sg13g2_decap_8 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_174 ();
 sg13g2_decap_8 FILLER_18_181 ();
 sg13g2_decap_8 FILLER_18_188 ();
 sg13g2_decap_8 FILLER_18_195 ();
 sg13g2_decap_8 FILLER_18_202 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_decap_8 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_237 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_11 ();
 sg13g2_decap_4 FILLER_19_17 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_66 ();
 sg13g2_fill_2 FILLER_19_107 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_decap_8 FILLER_19_150 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_decap_8 FILLER_19_164 ();
 sg13g2_decap_8 FILLER_19_171 ();
 sg13g2_decap_8 FILLER_19_178 ();
 sg13g2_decap_8 FILLER_19_185 ();
 sg13g2_decap_8 FILLER_19_192 ();
 sg13g2_decap_8 FILLER_19_199 ();
 sg13g2_decap_8 FILLER_19_206 ();
 sg13g2_decap_8 FILLER_19_213 ();
 sg13g2_decap_8 FILLER_19_220 ();
 sg13g2_decap_8 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_234 ();
 sg13g2_decap_8 FILLER_19_241 ();
 sg13g2_decap_8 FILLER_19_248 ();
 sg13g2_decap_8 FILLER_19_255 ();
 sg13g2_decap_8 FILLER_19_262 ();
 sg13g2_decap_8 FILLER_19_269 ();
 sg13g2_decap_8 FILLER_19_276 ();
 sg13g2_decap_8 FILLER_19_283 ();
 sg13g2_decap_8 FILLER_19_290 ();
 sg13g2_decap_8 FILLER_19_297 ();
 sg13g2_decap_8 FILLER_19_304 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_332 ();
 sg13g2_decap_8 FILLER_19_339 ();
 sg13g2_decap_8 FILLER_19_346 ();
 sg13g2_decap_8 FILLER_19_353 ();
 sg13g2_decap_8 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_367 ();
 sg13g2_decap_8 FILLER_19_374 ();
 sg13g2_decap_8 FILLER_19_381 ();
 sg13g2_decap_8 FILLER_19_388 ();
 sg13g2_decap_8 FILLER_19_395 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_4 ();
 sg13g2_fill_1 FILLER_20_33 ();
 sg13g2_fill_2 FILLER_20_47 ();
 sg13g2_fill_1 FILLER_20_61 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_148 ();
 sg13g2_decap_8 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_162 ();
 sg13g2_decap_8 FILLER_20_169 ();
 sg13g2_decap_8 FILLER_20_176 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_197 ();
 sg13g2_decap_8 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_218 ();
 sg13g2_decap_8 FILLER_20_225 ();
 sg13g2_decap_8 FILLER_20_232 ();
 sg13g2_decap_8 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_decap_8 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_20_337 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_decap_4 FILLER_21_26 ();
 sg13g2_fill_2 FILLER_21_61 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_2 FILLER_21_101 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_40 ();
 sg13g2_fill_1 FILLER_22_68 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_13 ();
 sg13g2_fill_1 FILLER_23_20 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_fill_1 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_fill_1 FILLER_24_121 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_4 FILLER_24_147 ();
 sg13g2_fill_2 FILLER_24_151 ();
 sg13g2_fill_2 FILLER_24_181 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_fill_1 FILLER_24_212 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_fill_2 FILLER_24_226 ();
 sg13g2_fill_1 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_8 FILLER_24_289 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_decap_8 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_373 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_139 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_184 ();
 sg13g2_decap_4 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_25_203 ();
 sg13g2_decap_4 FILLER_25_213 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_fill_2 FILLER_25_326 ();
 sg13g2_fill_1 FILLER_25_328 ();
 sg13g2_decap_4 FILLER_25_333 ();
 sg13g2_decap_4 FILLER_25_346 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_fill_1 FILLER_26_95 ();
 sg13g2_fill_2 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_134 ();
 sg13g2_fill_2 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_226 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_fill_2 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_2 FILLER_26_287 ();
 sg13g2_fill_1 FILLER_26_289 ();
 sg13g2_fill_2 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_decap_4 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_373 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_90 ();
 sg13g2_decap_8 FILLER_27_122 ();
 sg13g2_decap_8 FILLER_27_129 ();
 sg13g2_decap_4 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_144 ();
 sg13g2_fill_2 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_251 ();
 sg13g2_fill_2 FILLER_27_258 ();
 sg13g2_fill_1 FILLER_27_260 ();
 sg13g2_decap_4 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_332 ();
 sg13g2_decap_4 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_34 ();
 sg13g2_fill_2 FILLER_28_54 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_decap_4 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_decap_4 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_319 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_decap_8 FILLER_29_103 ();
 sg13g2_decap_8 FILLER_29_110 ();
 sg13g2_decap_4 FILLER_29_117 ();
 sg13g2_fill_2 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_206 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_2 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_316 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_decap_8 FILLER_29_398 ();
 sg13g2_decap_4 FILLER_29_405 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_4 FILLER_30_21 ();
 sg13g2_fill_2 FILLER_30_25 ();
 sg13g2_fill_2 FILLER_30_58 ();
 sg13g2_decap_8 FILLER_30_92 ();
 sg13g2_decap_8 FILLER_30_99 ();
 sg13g2_decap_8 FILLER_30_106 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_fill_2 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_248 ();
 sg13g2_decap_8 FILLER_30_255 ();
 sg13g2_fill_2 FILLER_30_262 ();
 sg13g2_decap_4 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_310 ();
 sg13g2_decap_4 FILLER_30_321 ();
 sg13g2_fill_2 FILLER_30_358 ();
 sg13g2_decap_8 FILLER_30_390 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_fill_1 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_80 ();
 sg13g2_decap_4 FILLER_31_113 ();
 sg13g2_fill_1 FILLER_31_117 ();
 sg13g2_decap_4 FILLER_31_122 ();
 sg13g2_fill_2 FILLER_31_126 ();
 sg13g2_fill_1 FILLER_31_155 ();
 sg13g2_decap_8 FILLER_31_174 ();
 sg13g2_decap_4 FILLER_31_181 ();
 sg13g2_fill_1 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_decap_4 FILLER_31_259 ();
 sg13g2_fill_1 FILLER_31_263 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_decap_8 FILLER_31_379 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_decap_8 FILLER_31_393 ();
 sg13g2_decap_8 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_42 ();
 sg13g2_fill_1 FILLER_32_96 ();
 sg13g2_fill_2 FILLER_32_173 ();
 sg13g2_fill_1 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_decap_4 FILLER_32_218 ();
 sg13g2_decap_4 FILLER_32_240 ();
 sg13g2_decap_8 FILLER_32_248 ();
 sg13g2_decap_8 FILLER_32_255 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_fill_1 FILLER_32_286 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_decap_8 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_313 ();
 sg13g2_decap_8 FILLER_32_318 ();
 sg13g2_decap_8 FILLER_32_325 ();
 sg13g2_decap_4 FILLER_32_332 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_53 ();
 sg13g2_fill_1 FILLER_33_62 ();
 sg13g2_decap_4 FILLER_33_96 ();
 sg13g2_fill_1 FILLER_33_100 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_decap_4 FILLER_33_234 ();
 sg13g2_fill_1 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_fill_2 FILLER_33_362 ();
 sg13g2_fill_2 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_60 ();
 sg13g2_decap_4 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_105 ();
 sg13g2_fill_1 FILLER_34_143 ();
 sg13g2_fill_2 FILLER_34_181 ();
 sg13g2_fill_1 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_decap_8 FILLER_34_245 ();
 sg13g2_fill_2 FILLER_34_269 ();
 sg13g2_decap_4 FILLER_34_284 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_decap_4 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_312 ();
 sg13g2_fill_1 FILLER_34_327 ();
 sg13g2_fill_2 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_4 FILLER_35_74 ();
 sg13g2_fill_2 FILLER_35_78 ();
 sg13g2_fill_2 FILLER_35_85 ();
 sg13g2_fill_1 FILLER_35_87 ();
 sg13g2_fill_2 FILLER_35_97 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_180 ();
 sg13g2_fill_1 FILLER_35_182 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_fill_1 FILLER_35_248 ();
 sg13g2_fill_2 FILLER_35_362 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_383 ();
 sg13g2_decap_8 FILLER_35_390 ();
 sg13g2_decap_8 FILLER_35_397 ();
 sg13g2_decap_4 FILLER_35_404 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_4 FILLER_36_98 ();
 sg13g2_fill_2 FILLER_36_102 ();
 sg13g2_fill_2 FILLER_36_126 ();
 sg13g2_fill_1 FILLER_36_168 ();
 sg13g2_fill_1 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_4 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_297 ();
 sg13g2_fill_1 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_4 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_fill_2 FILLER_37_138 ();
 sg13g2_fill_2 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_219 ();
 sg13g2_decap_4 FILLER_37_230 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_fill_1 FILLER_38_63 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_240 ();
 sg13g2_decap_4 FILLER_38_245 ();
 sg13g2_fill_2 FILLER_38_289 ();
 sg13g2_fill_1 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_296 ();
 sg13g2_decap_8 FILLER_38_303 ();
 sg13g2_decap_4 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_314 ();
 sg13g2_fill_1 FILLER_38_320 ();
 sg13g2_fill_1 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net90;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_out[6] = net10;
endmodule
