module tt_um_themightyduckofdoom_bitserial_collatz_checker (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire \bit_counter_q[0] ;
 wire \bit_counter_q[1] ;
 wire \bit_counter_q[2] ;
 wire \bit_counter_q[3] ;
 wire \bit_counter_q[4] ;
 wire \bit_counter_q[5] ;
 wire \bit_counter_q[6] ;
 wire \bit_counter_q[7] ;
 wire \bit_counter_q[8] ;
 wire \bit_counter_q[9] ;
 wire carry_q;
 wire finished_q;
 wire \i_main_reg.data_d[0] ;
 wire \i_main_reg.data_d[100] ;
 wire \i_main_reg.data_d[101] ;
 wire \i_main_reg.data_d[102] ;
 wire \i_main_reg.data_d[103] ;
 wire \i_main_reg.data_d[104] ;
 wire \i_main_reg.data_d[105] ;
 wire \i_main_reg.data_d[106] ;
 wire \i_main_reg.data_d[107] ;
 wire \i_main_reg.data_d[108] ;
 wire \i_main_reg.data_d[109] ;
 wire \i_main_reg.data_d[10] ;
 wire \i_main_reg.data_d[110] ;
 wire \i_main_reg.data_d[111] ;
 wire \i_main_reg.data_d[112] ;
 wire \i_main_reg.data_d[113] ;
 wire \i_main_reg.data_d[114] ;
 wire \i_main_reg.data_d[115] ;
 wire \i_main_reg.data_d[116] ;
 wire \i_main_reg.data_d[117] ;
 wire \i_main_reg.data_d[118] ;
 wire \i_main_reg.data_d[119] ;
 wire \i_main_reg.data_d[11] ;
 wire \i_main_reg.data_d[120] ;
 wire \i_main_reg.data_d[121] ;
 wire \i_main_reg.data_d[122] ;
 wire \i_main_reg.data_d[123] ;
 wire \i_main_reg.data_d[124] ;
 wire \i_main_reg.data_d[125] ;
 wire \i_main_reg.data_d[126] ;
 wire \i_main_reg.data_d[127] ;
 wire \i_main_reg.data_d[128] ;
 wire \i_main_reg.data_d[129] ;
 wire \i_main_reg.data_d[12] ;
 wire \i_main_reg.data_d[130] ;
 wire \i_main_reg.data_d[131] ;
 wire \i_main_reg.data_d[132] ;
 wire \i_main_reg.data_d[133] ;
 wire \i_main_reg.data_d[134] ;
 wire \i_main_reg.data_d[135] ;
 wire \i_main_reg.data_d[136] ;
 wire \i_main_reg.data_d[137] ;
 wire \i_main_reg.data_d[138] ;
 wire \i_main_reg.data_d[139] ;
 wire \i_main_reg.data_d[13] ;
 wire \i_main_reg.data_d[140] ;
 wire \i_main_reg.data_d[141] ;
 wire \i_main_reg.data_d[142] ;
 wire \i_main_reg.data_d[143] ;
 wire \i_main_reg.data_d[144] ;
 wire \i_main_reg.data_d[145] ;
 wire \i_main_reg.data_d[146] ;
 wire \i_main_reg.data_d[147] ;
 wire \i_main_reg.data_d[148] ;
 wire \i_main_reg.data_d[149] ;
 wire \i_main_reg.data_d[14] ;
 wire \i_main_reg.data_d[150] ;
 wire \i_main_reg.data_d[151] ;
 wire \i_main_reg.data_d[152] ;
 wire \i_main_reg.data_d[153] ;
 wire \i_main_reg.data_d[154] ;
 wire \i_main_reg.data_d[155] ;
 wire \i_main_reg.data_d[156] ;
 wire \i_main_reg.data_d[157] ;
 wire \i_main_reg.data_d[158] ;
 wire \i_main_reg.data_d[159] ;
 wire \i_main_reg.data_d[15] ;
 wire \i_main_reg.data_d[160] ;
 wire \i_main_reg.data_d[161] ;
 wire \i_main_reg.data_d[162] ;
 wire \i_main_reg.data_d[163] ;
 wire \i_main_reg.data_d[164] ;
 wire \i_main_reg.data_d[165] ;
 wire \i_main_reg.data_d[166] ;
 wire \i_main_reg.data_d[167] ;
 wire \i_main_reg.data_d[168] ;
 wire \i_main_reg.data_d[169] ;
 wire \i_main_reg.data_d[16] ;
 wire \i_main_reg.data_d[170] ;
 wire \i_main_reg.data_d[171] ;
 wire \i_main_reg.data_d[172] ;
 wire \i_main_reg.data_d[173] ;
 wire \i_main_reg.data_d[174] ;
 wire \i_main_reg.data_d[175] ;
 wire \i_main_reg.data_d[176] ;
 wire \i_main_reg.data_d[177] ;
 wire \i_main_reg.data_d[178] ;
 wire \i_main_reg.data_d[179] ;
 wire \i_main_reg.data_d[17] ;
 wire \i_main_reg.data_d[180] ;
 wire \i_main_reg.data_d[181] ;
 wire \i_main_reg.data_d[182] ;
 wire \i_main_reg.data_d[183] ;
 wire \i_main_reg.data_d[184] ;
 wire \i_main_reg.data_d[185] ;
 wire \i_main_reg.data_d[186] ;
 wire \i_main_reg.data_d[187] ;
 wire \i_main_reg.data_d[188] ;
 wire \i_main_reg.data_d[189] ;
 wire \i_main_reg.data_d[18] ;
 wire \i_main_reg.data_d[190] ;
 wire \i_main_reg.data_d[191] ;
 wire \i_main_reg.data_d[192] ;
 wire \i_main_reg.data_d[193] ;
 wire \i_main_reg.data_d[194] ;
 wire \i_main_reg.data_d[195] ;
 wire \i_main_reg.data_d[196] ;
 wire \i_main_reg.data_d[197] ;
 wire \i_main_reg.data_d[198] ;
 wire \i_main_reg.data_d[199] ;
 wire \i_main_reg.data_d[19] ;
 wire \i_main_reg.data_d[1] ;
 wire \i_main_reg.data_d[200] ;
 wire \i_main_reg.data_d[201] ;
 wire \i_main_reg.data_d[202] ;
 wire \i_main_reg.data_d[203] ;
 wire \i_main_reg.data_d[204] ;
 wire \i_main_reg.data_d[205] ;
 wire \i_main_reg.data_d[206] ;
 wire \i_main_reg.data_d[207] ;
 wire \i_main_reg.data_d[208] ;
 wire \i_main_reg.data_d[209] ;
 wire \i_main_reg.data_d[20] ;
 wire \i_main_reg.data_d[210] ;
 wire \i_main_reg.data_d[211] ;
 wire \i_main_reg.data_d[212] ;
 wire \i_main_reg.data_d[213] ;
 wire \i_main_reg.data_d[214] ;
 wire \i_main_reg.data_d[215] ;
 wire \i_main_reg.data_d[216] ;
 wire \i_main_reg.data_d[217] ;
 wire \i_main_reg.data_d[218] ;
 wire \i_main_reg.data_d[219] ;
 wire \i_main_reg.data_d[21] ;
 wire \i_main_reg.data_d[220] ;
 wire \i_main_reg.data_d[221] ;
 wire \i_main_reg.data_d[222] ;
 wire \i_main_reg.data_d[223] ;
 wire \i_main_reg.data_d[224] ;
 wire \i_main_reg.data_d[225] ;
 wire \i_main_reg.data_d[226] ;
 wire \i_main_reg.data_d[227] ;
 wire \i_main_reg.data_d[228] ;
 wire \i_main_reg.data_d[229] ;
 wire \i_main_reg.data_d[22] ;
 wire \i_main_reg.data_d[230] ;
 wire \i_main_reg.data_d[231] ;
 wire \i_main_reg.data_d[232] ;
 wire \i_main_reg.data_d[233] ;
 wire \i_main_reg.data_d[234] ;
 wire \i_main_reg.data_d[235] ;
 wire \i_main_reg.data_d[236] ;
 wire \i_main_reg.data_d[237] ;
 wire \i_main_reg.data_d[238] ;
 wire \i_main_reg.data_d[239] ;
 wire \i_main_reg.data_d[23] ;
 wire \i_main_reg.data_d[240] ;
 wire \i_main_reg.data_d[241] ;
 wire \i_main_reg.data_d[242] ;
 wire \i_main_reg.data_d[243] ;
 wire \i_main_reg.data_d[244] ;
 wire \i_main_reg.data_d[245] ;
 wire \i_main_reg.data_d[246] ;
 wire \i_main_reg.data_d[247] ;
 wire \i_main_reg.data_d[248] ;
 wire \i_main_reg.data_d[249] ;
 wire \i_main_reg.data_d[24] ;
 wire \i_main_reg.data_d[250] ;
 wire \i_main_reg.data_d[251] ;
 wire \i_main_reg.data_d[252] ;
 wire \i_main_reg.data_d[253] ;
 wire \i_main_reg.data_d[254] ;
 wire \i_main_reg.data_d[255] ;
 wire \i_main_reg.data_d[256] ;
 wire \i_main_reg.data_d[257] ;
 wire \i_main_reg.data_d[258] ;
 wire \i_main_reg.data_d[259] ;
 wire \i_main_reg.data_d[25] ;
 wire \i_main_reg.data_d[260] ;
 wire \i_main_reg.data_d[261] ;
 wire \i_main_reg.data_d[262] ;
 wire \i_main_reg.data_d[263] ;
 wire \i_main_reg.data_d[264] ;
 wire \i_main_reg.data_d[265] ;
 wire \i_main_reg.data_d[266] ;
 wire \i_main_reg.data_d[267] ;
 wire \i_main_reg.data_d[268] ;
 wire \i_main_reg.data_d[269] ;
 wire \i_main_reg.data_d[26] ;
 wire \i_main_reg.data_d[270] ;
 wire \i_main_reg.data_d[271] ;
 wire \i_main_reg.data_d[272] ;
 wire \i_main_reg.data_d[273] ;
 wire \i_main_reg.data_d[274] ;
 wire \i_main_reg.data_d[275] ;
 wire \i_main_reg.data_d[276] ;
 wire \i_main_reg.data_d[277] ;
 wire \i_main_reg.data_d[278] ;
 wire \i_main_reg.data_d[279] ;
 wire \i_main_reg.data_d[27] ;
 wire \i_main_reg.data_d[280] ;
 wire \i_main_reg.data_d[281] ;
 wire \i_main_reg.data_d[282] ;
 wire \i_main_reg.data_d[283] ;
 wire \i_main_reg.data_d[284] ;
 wire \i_main_reg.data_d[285] ;
 wire \i_main_reg.data_d[286] ;
 wire \i_main_reg.data_d[287] ;
 wire \i_main_reg.data_d[288] ;
 wire \i_main_reg.data_d[289] ;
 wire \i_main_reg.data_d[28] ;
 wire \i_main_reg.data_d[290] ;
 wire \i_main_reg.data_d[291] ;
 wire \i_main_reg.data_d[292] ;
 wire \i_main_reg.data_d[293] ;
 wire \i_main_reg.data_d[294] ;
 wire \i_main_reg.data_d[295] ;
 wire \i_main_reg.data_d[296] ;
 wire \i_main_reg.data_d[297] ;
 wire \i_main_reg.data_d[298] ;
 wire \i_main_reg.data_d[299] ;
 wire \i_main_reg.data_d[29] ;
 wire \i_main_reg.data_d[2] ;
 wire \i_main_reg.data_d[300] ;
 wire \i_main_reg.data_d[301] ;
 wire \i_main_reg.data_d[302] ;
 wire \i_main_reg.data_d[303] ;
 wire \i_main_reg.data_d[304] ;
 wire \i_main_reg.data_d[305] ;
 wire \i_main_reg.data_d[306] ;
 wire \i_main_reg.data_d[307] ;
 wire \i_main_reg.data_d[308] ;
 wire \i_main_reg.data_d[309] ;
 wire \i_main_reg.data_d[30] ;
 wire \i_main_reg.data_d[310] ;
 wire \i_main_reg.data_d[311] ;
 wire \i_main_reg.data_d[312] ;
 wire \i_main_reg.data_d[313] ;
 wire \i_main_reg.data_d[314] ;
 wire \i_main_reg.data_d[315] ;
 wire \i_main_reg.data_d[316] ;
 wire \i_main_reg.data_d[317] ;
 wire \i_main_reg.data_d[318] ;
 wire \i_main_reg.data_d[319] ;
 wire \i_main_reg.data_d[31] ;
 wire \i_main_reg.data_d[320] ;
 wire \i_main_reg.data_d[321] ;
 wire \i_main_reg.data_d[322] ;
 wire \i_main_reg.data_d[323] ;
 wire \i_main_reg.data_d[324] ;
 wire \i_main_reg.data_d[325] ;
 wire \i_main_reg.data_d[326] ;
 wire \i_main_reg.data_d[327] ;
 wire \i_main_reg.data_d[328] ;
 wire \i_main_reg.data_d[329] ;
 wire \i_main_reg.data_d[32] ;
 wire \i_main_reg.data_d[330] ;
 wire \i_main_reg.data_d[331] ;
 wire \i_main_reg.data_d[332] ;
 wire \i_main_reg.data_d[333] ;
 wire \i_main_reg.data_d[334] ;
 wire \i_main_reg.data_d[335] ;
 wire \i_main_reg.data_d[336] ;
 wire \i_main_reg.data_d[337] ;
 wire \i_main_reg.data_d[338] ;
 wire \i_main_reg.data_d[339] ;
 wire \i_main_reg.data_d[33] ;
 wire \i_main_reg.data_d[340] ;
 wire \i_main_reg.data_d[341] ;
 wire \i_main_reg.data_d[342] ;
 wire \i_main_reg.data_d[343] ;
 wire \i_main_reg.data_d[344] ;
 wire \i_main_reg.data_d[345] ;
 wire \i_main_reg.data_d[346] ;
 wire \i_main_reg.data_d[347] ;
 wire \i_main_reg.data_d[348] ;
 wire \i_main_reg.data_d[349] ;
 wire \i_main_reg.data_d[34] ;
 wire \i_main_reg.data_d[350] ;
 wire \i_main_reg.data_d[351] ;
 wire \i_main_reg.data_d[352] ;
 wire \i_main_reg.data_d[353] ;
 wire \i_main_reg.data_d[354] ;
 wire \i_main_reg.data_d[355] ;
 wire \i_main_reg.data_d[356] ;
 wire \i_main_reg.data_d[357] ;
 wire \i_main_reg.data_d[358] ;
 wire \i_main_reg.data_d[359] ;
 wire \i_main_reg.data_d[35] ;
 wire \i_main_reg.data_d[360] ;
 wire \i_main_reg.data_d[361] ;
 wire \i_main_reg.data_d[362] ;
 wire \i_main_reg.data_d[363] ;
 wire \i_main_reg.data_d[364] ;
 wire \i_main_reg.data_d[365] ;
 wire \i_main_reg.data_d[366] ;
 wire \i_main_reg.data_d[367] ;
 wire \i_main_reg.data_d[368] ;
 wire \i_main_reg.data_d[369] ;
 wire \i_main_reg.data_d[36] ;
 wire \i_main_reg.data_d[370] ;
 wire \i_main_reg.data_d[371] ;
 wire \i_main_reg.data_d[372] ;
 wire \i_main_reg.data_d[373] ;
 wire \i_main_reg.data_d[374] ;
 wire \i_main_reg.data_d[375] ;
 wire \i_main_reg.data_d[376] ;
 wire \i_main_reg.data_d[377] ;
 wire \i_main_reg.data_d[378] ;
 wire \i_main_reg.data_d[379] ;
 wire \i_main_reg.data_d[37] ;
 wire \i_main_reg.data_d[380] ;
 wire \i_main_reg.data_d[381] ;
 wire \i_main_reg.data_d[382] ;
 wire \i_main_reg.data_d[38] ;
 wire \i_main_reg.data_d[39] ;
 wire \i_main_reg.data_d[3] ;
 wire \i_main_reg.data_d[40] ;
 wire \i_main_reg.data_d[41] ;
 wire \i_main_reg.data_d[42] ;
 wire \i_main_reg.data_d[43] ;
 wire \i_main_reg.data_d[44] ;
 wire \i_main_reg.data_d[45] ;
 wire \i_main_reg.data_d[46] ;
 wire \i_main_reg.data_d[47] ;
 wire \i_main_reg.data_d[48] ;
 wire \i_main_reg.data_d[49] ;
 wire \i_main_reg.data_d[4] ;
 wire \i_main_reg.data_d[50] ;
 wire \i_main_reg.data_d[51] ;
 wire \i_main_reg.data_d[52] ;
 wire \i_main_reg.data_d[53] ;
 wire \i_main_reg.data_d[54] ;
 wire \i_main_reg.data_d[55] ;
 wire \i_main_reg.data_d[56] ;
 wire \i_main_reg.data_d[57] ;
 wire \i_main_reg.data_d[58] ;
 wire \i_main_reg.data_d[59] ;
 wire \i_main_reg.data_d[5] ;
 wire \i_main_reg.data_d[60] ;
 wire \i_main_reg.data_d[61] ;
 wire \i_main_reg.data_d[62] ;
 wire \i_main_reg.data_d[63] ;
 wire \i_main_reg.data_d[64] ;
 wire \i_main_reg.data_d[65] ;
 wire \i_main_reg.data_d[66] ;
 wire \i_main_reg.data_d[67] ;
 wire \i_main_reg.data_d[68] ;
 wire \i_main_reg.data_d[69] ;
 wire \i_main_reg.data_d[6] ;
 wire \i_main_reg.data_d[70] ;
 wire \i_main_reg.data_d[71] ;
 wire \i_main_reg.data_d[72] ;
 wire \i_main_reg.data_d[73] ;
 wire \i_main_reg.data_d[74] ;
 wire \i_main_reg.data_d[75] ;
 wire \i_main_reg.data_d[76] ;
 wire \i_main_reg.data_d[77] ;
 wire \i_main_reg.data_d[78] ;
 wire \i_main_reg.data_d[79] ;
 wire \i_main_reg.data_d[7] ;
 wire \i_main_reg.data_d[80] ;
 wire \i_main_reg.data_d[81] ;
 wire \i_main_reg.data_d[82] ;
 wire \i_main_reg.data_d[83] ;
 wire \i_main_reg.data_d[84] ;
 wire \i_main_reg.data_d[85] ;
 wire \i_main_reg.data_d[86] ;
 wire \i_main_reg.data_d[87] ;
 wire \i_main_reg.data_d[88] ;
 wire \i_main_reg.data_d[89] ;
 wire \i_main_reg.data_d[8] ;
 wire \i_main_reg.data_d[90] ;
 wire \i_main_reg.data_d[91] ;
 wire \i_main_reg.data_d[92] ;
 wire \i_main_reg.data_d[93] ;
 wire \i_main_reg.data_d[94] ;
 wire \i_main_reg.data_d[95] ;
 wire \i_main_reg.data_d[96] ;
 wire \i_main_reg.data_d[97] ;
 wire \i_main_reg.data_d[98] ;
 wire \i_main_reg.data_d[99] ;
 wire \i_main_reg.data_d[9] ;
 wire \i_main_reg.data_o ;
 wire \i_step_counter.data_d[0] ;
 wire \i_step_counter.data_d[10] ;
 wire \i_step_counter.data_d[11] ;
 wire \i_step_counter.data_d[12] ;
 wire \i_step_counter.data_d[13] ;
 wire \i_step_counter.data_d[14] ;
 wire \i_step_counter.data_d[1] ;
 wire \i_step_counter.data_d[2] ;
 wire \i_step_counter.data_d[3] ;
 wire \i_step_counter.data_d[4] ;
 wire \i_step_counter.data_d[5] ;
 wire \i_step_counter.data_d[6] ;
 wire \i_step_counter.data_d[7] ;
 wire \i_step_counter.data_d[8] ;
 wire \i_step_counter.data_d[9] ;
 wire \i_step_counter.data_o ;
 wire \one_count_q[0] ;
 wire \one_count_q[1] ;
 wire overflow_q;
 wire previous_bit_q;
 wire \state_q[0] ;
 wire \state_q[1] ;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire clknet_leaf_0_clk;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;

 sg13g2_inv_1 _0555_ (.Y(_0432_),
    .A(net774));
 sg13g2_inv_1 _0556_ (.Y(_0433_),
    .A(net715));
 sg13g2_inv_1 _0557_ (.Y(_0434_),
    .A(\i_step_counter.data_d[0] ));
 sg13g2_inv_1 _0558_ (.Y(_0435_),
    .A(net709));
 sg13g2_inv_1 _0559_ (.Y(_0436_),
    .A(\i_step_counter.data_d[1] ));
 sg13g2_inv_1 _0560_ (.Y(_0437_),
    .A(net34));
 sg13g2_inv_1 _0561_ (.Y(_0438_),
    .A(\i_step_counter.data_d[12] ));
 sg13g2_inv_1 _0562_ (.Y(_0439_),
    .A(net755));
 sg13g2_nor2b_2 _0563_ (.A(\state_q[0] ),
    .B_N(\state_q[1] ),
    .Y(_0440_));
 sg13g2_nand2b_1 _0564_ (.Y(_0441_),
    .B(\state_q[1] ),
    .A_N(\state_q[0] ));
 sg13g2_a21oi_2 _0565_ (.B1(net33),
    .Y(_0442_),
    .A2(\bit_counter_q[7] ),
    .A1(\bit_counter_q[8] ));
 sg13g2_a21o_2 _0566_ (.A2(\bit_counter_q[7] ),
    .A1(\bit_counter_q[8] ),
    .B1(net33),
    .X(_0443_));
 sg13g2_nor2b_1 _0567_ (.A(net378),
    .B_N(net31),
    .Y(_0444_));
 sg13g2_nor2_1 _0568_ (.A(net753),
    .B(net31),
    .Y(_0445_));
 sg13g2_nor2b_1 _0569_ (.A(net753),
    .B_N(net378),
    .Y(_0446_));
 sg13g2_nor4_1 _0570_ (.A(net376),
    .B(_0442_),
    .C(_0445_),
    .D(_0446_),
    .Y(_0447_));
 sg13g2_nor2_1 _0571_ (.A(\state_q[0] ),
    .B(\state_q[1] ),
    .Y(_0448_));
 sg13g2_and2_1 _0572_ (.A(net3),
    .B(_0448_),
    .X(_0449_));
 sg13g2_o21ai_1 _0573_ (.B1(_0448_),
    .Y(_0450_),
    .A1(net4),
    .A2(net3));
 sg13g2_nor2b_2 _0574_ (.A(net375),
    .B_N(_0450_),
    .Y(_0451_));
 sg13g2_nand2b_1 _0575_ (.Y(_0452_),
    .B(_0450_),
    .A_N(net374));
 sg13g2_nor2_1 _0576_ (.A(net709),
    .B(net371),
    .Y(_0453_));
 sg13g2_a22oi_1 _0577_ (.Y(_0454_),
    .B1(net372),
    .B2(\i_step_counter.data_d[0] ),
    .A2(_0440_),
    .A1(_0435_));
 sg13g2_a21oi_1 _0578_ (.A1(_0452_),
    .A2(_0454_),
    .Y(_0000_),
    .B1(_0453_));
 sg13g2_nand2_1 _0579_ (.Y(_0455_),
    .A(net764),
    .B(net373));
 sg13g2_nor2_1 _0580_ (.A(_0434_),
    .B(_0435_),
    .Y(_0456_));
 sg13g2_o21ai_1 _0581_ (.B1(net371),
    .Y(_0457_),
    .A1(net376),
    .A2(_0456_));
 sg13g2_o21ai_1 _0582_ (.B1(_0457_),
    .Y(_0458_),
    .A1(\i_step_counter.data_d[0] ),
    .A2(net709));
 sg13g2_a22oi_1 _0583_ (.Y(_0001_),
    .B1(_0455_),
    .B2(_0458_),
    .A2(_0451_),
    .A1(_0434_));
 sg13g2_nand2_1 _0584_ (.Y(_0459_),
    .A(net725),
    .B(net373));
 sg13g2_or2_1 _0585_ (.X(_0460_),
    .B(_0456_),
    .A(\i_step_counter.data_d[1] ));
 sg13g2_nor2_1 _0586_ (.A(\i_step_counter.data_d[1] ),
    .B(net376),
    .Y(_0461_));
 sg13g2_o21ai_1 _0587_ (.B1(_0460_),
    .Y(_0462_),
    .A1(_0457_),
    .A2(_0461_));
 sg13g2_a22oi_1 _0588_ (.Y(_0002_),
    .B1(_0459_),
    .B2(_0462_),
    .A2(_0451_),
    .A1(_0436_));
 sg13g2_nand4_1 _0589_ (.B(net709),
    .C(net764),
    .A(net769),
    .Y(_0463_),
    .D(net725));
 sg13g2_nand4_1 _0590_ (.B(\i_step_counter.data_d[2] ),
    .C(net375),
    .A(\i_step_counter.data_d[1] ),
    .Y(_0464_),
    .D(_0456_));
 sg13g2_a21o_1 _0591_ (.A2(_0456_),
    .A1(net764),
    .B1(net725),
    .X(_0465_));
 sg13g2_nand3_1 _0592_ (.B(_0463_),
    .C(_0465_),
    .A(net375),
    .Y(_0466_));
 sg13g2_a22oi_1 _0593_ (.Y(_0467_),
    .B1(_0451_),
    .B2(net725),
    .A2(net373),
    .A1(net34));
 sg13g2_nand2_1 _0594_ (.Y(_0003_),
    .A(_0466_),
    .B(_0467_));
 sg13g2_nor2_1 _0595_ (.A(_0437_),
    .B(_0463_),
    .Y(_0468_));
 sg13g2_o21ai_1 _0596_ (.B1(net371),
    .Y(_0469_),
    .A1(net376),
    .A2(_0468_));
 sg13g2_a22oi_1 _0597_ (.Y(_0470_),
    .B1(_0469_),
    .B2(net34),
    .A2(net373),
    .A1(\i_step_counter.data_d[4] ));
 sg13g2_o21ai_1 _0598_ (.B1(_0470_),
    .Y(_0004_),
    .A1(net34),
    .A2(_0464_));
 sg13g2_nand3b_1 _0599_ (.B(net374),
    .C(_0468_),
    .Y(_0471_),
    .A_N(net771));
 sg13g2_a22oi_1 _0600_ (.Y(_0472_),
    .B1(_0469_),
    .B2(net771),
    .A2(net373),
    .A1(\i_step_counter.data_d[5] ));
 sg13g2_nand2_1 _0601_ (.Y(_0005_),
    .A(_0471_),
    .B(net772));
 sg13g2_nand2_1 _0602_ (.Y(_0473_),
    .A(net41),
    .B(net373));
 sg13g2_and3_1 _0603_ (.X(_0474_),
    .A(net771),
    .B(net773),
    .C(_0468_));
 sg13g2_o21ai_1 _0604_ (.B1(net371),
    .Y(_0475_),
    .A1(net376),
    .A2(_0474_));
 sg13g2_and3_1 _0605_ (.X(_0476_),
    .A(\i_step_counter.data_d[4] ),
    .B(net371),
    .C(_0468_));
 sg13g2_o21ai_1 _0606_ (.B1(_0475_),
    .Y(_0477_),
    .A1(\i_step_counter.data_d[5] ),
    .A2(_0476_));
 sg13g2_nand2_1 _0607_ (.Y(_0006_),
    .A(_0473_),
    .B(_0477_));
 sg13g2_nand3b_1 _0608_ (.B(net374),
    .C(_0474_),
    .Y(_0478_),
    .A_N(net41));
 sg13g2_a22oi_1 _0609_ (.Y(_0479_),
    .B1(_0475_),
    .B2(net41),
    .A2(net372),
    .A1(net770));
 sg13g2_nand2_1 _0610_ (.Y(_0007_),
    .A(_0478_),
    .B(_0479_));
 sg13g2_nand4_1 _0611_ (.B(net771),
    .C(net773),
    .A(net34),
    .Y(_0480_),
    .D(net41));
 sg13g2_nor2_2 _0612_ (.A(_0463_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_and2_1 _0613_ (.A(net770),
    .B(_0481_),
    .X(_0482_));
 sg13g2_o21ai_1 _0614_ (.B1(net371),
    .Y(_0483_),
    .A1(net376),
    .A2(_0482_));
 sg13g2_nand3b_1 _0615_ (.B(net374),
    .C(_0481_),
    .Y(_0484_),
    .A_N(net770));
 sg13g2_a22oi_1 _0616_ (.Y(_0485_),
    .B1(_0483_),
    .B2(net770),
    .A2(net372),
    .A1(net766));
 sg13g2_nand2_1 _0617_ (.Y(_0008_),
    .A(_0484_),
    .B(_0485_));
 sg13g2_a22oi_1 _0618_ (.Y(_0486_),
    .B1(_0483_),
    .B2(net766),
    .A2(net372),
    .A1(net740));
 sg13g2_nand3b_1 _0619_ (.B(net374),
    .C(_0482_),
    .Y(_0487_),
    .A_N(net766));
 sg13g2_nand2_1 _0620_ (.Y(_0009_),
    .A(_0486_),
    .B(_0487_));
 sg13g2_and4_1 _0621_ (.A(\i_step_counter.data_d[7] ),
    .B(net766),
    .C(net740),
    .D(_0481_),
    .X(_0488_));
 sg13g2_o21ai_1 _0622_ (.B1(net371),
    .Y(_0489_),
    .A1(net376),
    .A2(_0488_));
 sg13g2_a22oi_1 _0623_ (.Y(_0490_),
    .B1(_0489_),
    .B2(net740),
    .A2(net372),
    .A1(\i_step_counter.data_d[10] ));
 sg13g2_nand4_1 _0624_ (.B(net766),
    .C(net374),
    .A(\i_step_counter.data_d[7] ),
    .Y(_0491_),
    .D(_0481_));
 sg13g2_o21ai_1 _0625_ (.B1(_0490_),
    .Y(_0010_),
    .A1(_0488_),
    .A2(net767));
 sg13g2_nand2b_1 _0626_ (.Y(_0492_),
    .B(net740),
    .A_N(\i_step_counter.data_d[10] ));
 sg13g2_a22oi_1 _0627_ (.Y(_0493_),
    .B1(_0489_),
    .B2(\i_step_counter.data_d[10] ),
    .A2(net372),
    .A1(net719));
 sg13g2_o21ai_1 _0628_ (.B1(_0493_),
    .Y(_0011_),
    .A1(_0491_),
    .A2(net741));
 sg13g2_and4_1 _0629_ (.A(net770),
    .B(net766),
    .C(net740),
    .D(\i_step_counter.data_d[10] ),
    .X(_0494_));
 sg13g2_and2_1 _0630_ (.A(\i_step_counter.data_d[11] ),
    .B(_0494_),
    .X(_0495_));
 sg13g2_and2_1 _0631_ (.A(_0481_),
    .B(_0495_),
    .X(_0496_));
 sg13g2_and2_1 _0632_ (.A(_0481_),
    .B(_0494_),
    .X(_0497_));
 sg13g2_o21ai_1 _0633_ (.B1(net371),
    .Y(_0498_),
    .A1(net376),
    .A2(_0496_));
 sg13g2_nand3b_1 _0634_ (.B(net374),
    .C(_0497_),
    .Y(_0499_),
    .A_N(net719));
 sg13g2_a22oi_1 _0635_ (.Y(_0500_),
    .B1(_0498_),
    .B2(net719),
    .A2(net372),
    .A1(net775));
 sg13g2_nand2_1 _0636_ (.Y(_0012_),
    .A(_0499_),
    .B(_0500_));
 sg13g2_nand4_1 _0637_ (.B(_0438_),
    .C(net374),
    .A(net719),
    .Y(_0501_),
    .D(_0497_));
 sg13g2_a22oi_1 _0638_ (.Y(_0502_),
    .B1(_0498_),
    .B2(\i_step_counter.data_d[12] ),
    .A2(net372),
    .A1(\i_step_counter.data_d[13] ));
 sg13g2_nand2_1 _0639_ (.Y(_0013_),
    .A(net720),
    .B(_0502_));
 sg13g2_nand4_1 _0640_ (.B(\i_step_counter.data_d[13] ),
    .C(_0481_),
    .A(\i_step_counter.data_d[12] ),
    .Y(_0503_),
    .D(_0495_));
 sg13g2_and3_1 _0641_ (.X(_0504_),
    .A(net719),
    .B(\i_step_counter.data_d[12] ),
    .C(_0497_));
 sg13g2_nand2_1 _0642_ (.Y(_0505_),
    .A(\i_step_counter.data_d[13] ),
    .B(_0504_));
 sg13g2_and2_1 _0643_ (.A(_0440_),
    .B(_0503_),
    .X(_0506_));
 sg13g2_o21ai_1 _0644_ (.B1(_0506_),
    .Y(_0507_),
    .A1(net755),
    .A2(_0504_));
 sg13g2_a21oi_1 _0645_ (.A1(net182),
    .A2(net373),
    .Y(_0508_),
    .B1(_0451_));
 sg13g2_a22oi_1 _0646_ (.Y(_0014_),
    .B1(_0507_),
    .B2(_0508_),
    .A2(_0451_),
    .A1(_0439_));
 sg13g2_o21ai_1 _0647_ (.B1(net182),
    .Y(_0509_),
    .A1(_0451_),
    .A2(_0506_));
 sg13g2_nand2b_1 _0648_ (.Y(_0510_),
    .B(net375),
    .A_N(net182));
 sg13g2_o21ai_1 _0649_ (.B1(net183),
    .Y(_0015_),
    .A1(_0505_),
    .A2(_0510_));
 sg13g2_nor4_2 _0650_ (.A(\one_count_q[1] ),
    .B(net377),
    .C(_0442_),
    .Y(_0511_),
    .D(_0444_));
 sg13g2_nor2_1 _0651_ (.A(net36),
    .B(_0511_),
    .Y(_0512_));
 sg13g2_a21oi_1 _0652_ (.A1(net4),
    .A2(_0448_),
    .Y(_0016_),
    .B1(net37));
 sg13g2_nor2_1 _0653_ (.A(net377),
    .B(_0443_),
    .Y(_0513_));
 sg13g2_nor3_2 _0654_ (.A(net777),
    .B(net774),
    .C(net4),
    .Y(_0514_));
 sg13g2_or2_1 _0655_ (.X(_0515_),
    .B(_0514_),
    .A(_0511_));
 sg13g2_nor4_1 _0656_ (.A(\state_q[0] ),
    .B(_0503_),
    .C(_0513_),
    .D(_0515_),
    .Y(_0516_));
 sg13g2_a21oi_1 _0657_ (.A1(\i_step_counter.data_d[14] ),
    .A2(_0516_),
    .Y(_0517_),
    .B1(net25));
 sg13g2_a21oi_1 _0658_ (.A1(net4),
    .A2(_0448_),
    .Y(_0017_),
    .B1(net26));
 sg13g2_nor3_1 _0659_ (.A(net379),
    .B(net377),
    .C(_0445_),
    .Y(_0518_));
 sg13g2_inv_1 _0660_ (.Y(_0519_),
    .A(_0518_));
 sg13g2_nand2b_2 _0661_ (.Y(_0520_),
    .B(net761),
    .A_N(\state_q[1] ));
 sg13g2_nor2_2 _0662_ (.A(_0443_),
    .B(_0520_),
    .Y(_0521_));
 sg13g2_o21ai_1 _0663_ (.B1(_0519_),
    .Y(_0522_),
    .A1(net375),
    .A2(_0521_));
 sg13g2_inv_1 _0664_ (.Y(_0030_),
    .A(_0522_));
 sg13g2_a21oi_1 _0665_ (.A1(net378),
    .A2(previous_bit_q),
    .Y(_0523_),
    .B1(_0520_));
 sg13g2_or2_1 _0666_ (.X(_0524_),
    .B(previous_bit_q),
    .A(net378));
 sg13g2_o21ai_1 _0667_ (.B1(net264),
    .Y(_0525_),
    .A1(_0522_),
    .A2(_0524_));
 sg13g2_o21ai_1 _0668_ (.B1(net265),
    .Y(_0018_),
    .A1(_0522_),
    .A2(_0523_));
 sg13g2_a22oi_1 _0669_ (.Y(_0526_),
    .B1(_0522_),
    .B2(net758),
    .A2(_0521_),
    .A1(net378));
 sg13g2_inv_1 _0670_ (.Y(_0019_),
    .A(net759));
 sg13g2_and2_1 _0671_ (.A(net777),
    .B(net778),
    .X(_0527_));
 sg13g2_nor2_2 _0672_ (.A(_0515_),
    .B(_0527_),
    .Y(_0528_));
 sg13g2_a21oi_2 _0673_ (.B1(_0443_),
    .Y(_0529_),
    .A2(_0520_),
    .A1(net377));
 sg13g2_inv_1 _0674_ (.Y(_0530_),
    .A(_0529_));
 sg13g2_nor3_2 _0675_ (.A(_0515_),
    .B(_0527_),
    .C(_0529_),
    .Y(_0531_));
 sg13g2_xnor2_1 _0676_ (.Y(_0532_),
    .A(net760),
    .B(_0528_));
 sg13g2_nor2_1 _0677_ (.A(_0531_),
    .B(_0532_),
    .Y(_0020_));
 sg13g2_a21oi_1 _0678_ (.A1(\bit_counter_q[0] ),
    .A2(_0528_),
    .Y(_0533_),
    .B1(net47));
 sg13g2_nand2_1 _0679_ (.Y(_0534_),
    .A(net760),
    .B(net47));
 sg13g2_nor4_2 _0680_ (.A(_0511_),
    .B(_0514_),
    .C(_0527_),
    .Y(_0535_),
    .D(_0534_));
 sg13g2_nor3_1 _0681_ (.A(_0531_),
    .B(net48),
    .C(_0535_),
    .Y(_0021_));
 sg13g2_nor2_1 _0682_ (.A(net763),
    .B(_0535_),
    .Y(_0536_));
 sg13g2_and2_1 _0683_ (.A(net763),
    .B(_0535_),
    .X(_0537_));
 sg13g2_nor3_1 _0684_ (.A(_0531_),
    .B(_0536_),
    .C(_0537_),
    .Y(_0022_));
 sg13g2_nor2_1 _0685_ (.A(net89),
    .B(_0537_),
    .Y(_0538_));
 sg13g2_and2_1 _0686_ (.A(\bit_counter_q[2] ),
    .B(net89),
    .X(_0539_));
 sg13g2_a221oi_1 _0687_ (.B2(_0539_),
    .C1(net90),
    .B1(_0535_),
    .A1(_0528_),
    .Y(_0023_),
    .A2(_0530_));
 sg13g2_a21oi_1 _0688_ (.A1(_0535_),
    .A2(_0539_),
    .Y(_0540_),
    .B1(net28));
 sg13g2_nand4_1 _0689_ (.B(\bit_counter_q[1] ),
    .C(net28),
    .A(\bit_counter_q[0] ),
    .Y(_0541_),
    .D(_0539_));
 sg13g2_nor4_1 _0690_ (.A(_0511_),
    .B(_0514_),
    .C(_0527_),
    .D(_0541_),
    .Y(_0542_));
 sg13g2_nor3_1 _0691_ (.A(_0531_),
    .B(net29),
    .C(_0542_),
    .Y(_0024_));
 sg13g2_nor2_1 _0692_ (.A(net43),
    .B(_0542_),
    .Y(_0543_));
 sg13g2_and2_1 _0693_ (.A(net43),
    .B(_0542_),
    .X(_0544_));
 sg13g2_nor3_1 _0694_ (.A(_0531_),
    .B(net44),
    .C(_0544_),
    .Y(_0025_));
 sg13g2_nor2_1 _0695_ (.A(net749),
    .B(_0544_),
    .Y(_0545_));
 sg13g2_a21oi_1 _0696_ (.A1(net749),
    .A2(_0544_),
    .Y(_0546_),
    .B1(_0531_));
 sg13g2_nor2b_1 _0697_ (.A(net750),
    .B_N(_0546_),
    .Y(_0026_));
 sg13g2_a21oi_1 _0698_ (.A1(\bit_counter_q[6] ),
    .A2(_0544_),
    .Y(_0547_),
    .B1(net745));
 sg13g2_and3_1 _0699_ (.X(_0548_),
    .A(net745),
    .B(\bit_counter_q[6] ),
    .C(_0544_));
 sg13g2_nand3_1 _0700_ (.B(\bit_counter_q[6] ),
    .C(_0544_),
    .A(\bit_counter_q[7] ),
    .Y(_0549_));
 sg13g2_nor3_1 _0701_ (.A(_0531_),
    .B(net746),
    .C(_0548_),
    .Y(_0027_));
 sg13g2_a21oi_1 _0702_ (.A1(_0433_),
    .A2(_0549_),
    .Y(_0028_),
    .B1(_0531_));
 sg13g2_nor2b_1 _0703_ (.A(_0528_),
    .B_N(net33),
    .Y(_0029_));
 sg13g2_nor3_1 _0704_ (.A(_0432_),
    .B(_0518_),
    .C(_0529_),
    .Y(_0550_));
 sg13g2_nor3_1 _0705_ (.A(_0514_),
    .B(_0521_),
    .C(_0550_),
    .Y(_0031_));
 sg13g2_nor2_1 _0706_ (.A(net2),
    .B(_0529_),
    .Y(_0551_));
 sg13g2_nor3_2 _0707_ (.A(net2),
    .B(_0518_),
    .C(_0529_),
    .Y(_0552_));
 sg13g2_nand2_1 _0708_ (.Y(_0553_),
    .A(_0519_),
    .B(_0551_));
 sg13g2_a22oi_1 _0709_ (.Y(_0554_),
    .B1(_0553_),
    .B2(net39),
    .A2(_0551_),
    .A1(net378));
 sg13g2_inv_1 _0710_ (.Y(_0032_),
    .A(net40));
 sg13g2_mux2_1 _0711_ (.A0(net241),
    .A1(net39),
    .S(net368),
    .X(_0033_));
 sg13g2_mux2_1 _0712_ (.A0(\i_main_reg.data_d[2] ),
    .A1(net241),
    .S(net368),
    .X(_0034_));
 sg13g2_mux2_1 _0713_ (.A0(\i_main_reg.data_d[3] ),
    .A1(net300),
    .S(net368),
    .X(_0035_));
 sg13g2_mux2_1 _0714_ (.A0(net675),
    .A1(net683),
    .S(net368),
    .X(_0036_));
 sg13g2_mux2_1 _0715_ (.A0(\i_main_reg.data_d[5] ),
    .A1(net675),
    .S(net366),
    .X(_0037_));
 sg13g2_mux2_1 _0716_ (.A0(net697),
    .A1(net729),
    .S(net366),
    .X(_0038_));
 sg13g2_mux2_1 _0717_ (.A0(\i_main_reg.data_d[7] ),
    .A1(net697),
    .S(net366),
    .X(_0039_));
 sg13g2_mux2_1 _0718_ (.A0(net699),
    .A1(\i_main_reg.data_d[7] ),
    .S(net361),
    .X(_0040_));
 sg13g2_mux2_1 _0719_ (.A0(net734),
    .A1(net699),
    .S(net362),
    .X(_0041_));
 sg13g2_mux2_1 _0720_ (.A0(net476),
    .A1(\i_main_reg.data_d[9] ),
    .S(net362),
    .X(_0042_));
 sg13g2_mux2_1 _0721_ (.A0(net509),
    .A1(net476),
    .S(net362),
    .X(_0043_));
 sg13g2_mux2_1 _0722_ (.A0(net534),
    .A1(net509),
    .S(net362),
    .X(_0044_));
 sg13g2_mux2_1 _0723_ (.A0(net596),
    .A1(net534),
    .S(net364),
    .X(_0045_));
 sg13g2_mux2_1 _0724_ (.A0(net494),
    .A1(net596),
    .S(net364),
    .X(_0046_));
 sg13g2_mux2_1 _0725_ (.A0(\i_main_reg.data_d[15] ),
    .A1(net494),
    .S(net364),
    .X(_0047_));
 sg13g2_mux2_1 _0726_ (.A0(net582),
    .A1(\i_main_reg.data_d[15] ),
    .S(net364),
    .X(_0048_));
 sg13g2_mux2_1 _0727_ (.A0(net613),
    .A1(net582),
    .S(net364),
    .X(_0049_));
 sg13g2_mux2_1 _0728_ (.A0(net283),
    .A1(net613),
    .S(net360),
    .X(_0050_));
 sg13g2_mux2_1 _0729_ (.A0(\i_main_reg.data_d[19] ),
    .A1(net283),
    .S(net359),
    .X(_0051_));
 sg13g2_mux2_1 _0730_ (.A0(\i_main_reg.data_d[20] ),
    .A1(net587),
    .S(net360),
    .X(_0052_));
 sg13g2_mux2_1 _0731_ (.A0(net50),
    .A1(\i_main_reg.data_d[20] ),
    .S(net360),
    .X(_0053_));
 sg13g2_mux2_1 _0732_ (.A0(net237),
    .A1(net50),
    .S(net360),
    .X(_0054_));
 sg13g2_mux2_1 _0733_ (.A0(\i_main_reg.data_d[23] ),
    .A1(net237),
    .S(net335),
    .X(_0055_));
 sg13g2_mux2_1 _0734_ (.A0(\i_main_reg.data_d[24] ),
    .A1(net504),
    .S(net334),
    .X(_0056_));
 sg13g2_mux2_1 _0735_ (.A0(net104),
    .A1(\i_main_reg.data_d[24] ),
    .S(net334),
    .X(_0057_));
 sg13g2_mux2_1 _0736_ (.A0(net230),
    .A1(net104),
    .S(net359),
    .X(_0058_));
 sg13g2_mux2_1 _0737_ (.A0(net113),
    .A1(net230),
    .S(net359),
    .X(_0059_));
 sg13g2_mux2_1 _0738_ (.A0(\i_main_reg.data_d[28] ),
    .A1(net113),
    .S(net359),
    .X(_0060_));
 sg13g2_mux2_1 _0739_ (.A0(net272),
    .A1(\i_main_reg.data_d[28] ),
    .S(net359),
    .X(_0061_));
 sg13g2_mux2_1 _0740_ (.A0(net151),
    .A1(\i_main_reg.data_d[29] ),
    .S(net359),
    .X(_0062_));
 sg13g2_mux2_1 _0741_ (.A0(net175),
    .A1(net151),
    .S(net359),
    .X(_0063_));
 sg13g2_mux2_1 _0742_ (.A0(net631),
    .A1(net175),
    .S(net359),
    .X(_0064_));
 sg13g2_mux2_1 _0743_ (.A0(\i_main_reg.data_d[33] ),
    .A1(net631),
    .S(net361),
    .X(_0065_));
 sg13g2_mux2_1 _0744_ (.A0(net454),
    .A1(net692),
    .S(net361),
    .X(_0066_));
 sg13g2_mux2_1 _0745_ (.A0(\i_main_reg.data_d[35] ),
    .A1(net454),
    .S(net361),
    .X(_0067_));
 sg13g2_mux2_1 _0746_ (.A0(net606),
    .A1(net693),
    .S(net361),
    .X(_0068_));
 sg13g2_mux2_1 _0747_ (.A0(net577),
    .A1(net606),
    .S(net361),
    .X(_0069_));
 sg13g2_mux2_1 _0748_ (.A0(\i_main_reg.data_d[38] ),
    .A1(net577),
    .S(net361),
    .X(_0070_));
 sg13g2_mux2_1 _0749_ (.A0(\i_main_reg.data_d[39] ),
    .A1(net694),
    .S(net361),
    .X(_0071_));
 sg13g2_mux2_1 _0750_ (.A0(net609),
    .A1(net739),
    .S(net369),
    .X(_0072_));
 sg13g2_mux2_1 _0751_ (.A0(net254),
    .A1(net609),
    .S(net369),
    .X(_0073_));
 sg13g2_mux2_1 _0752_ (.A0(\i_main_reg.data_d[42] ),
    .A1(net254),
    .S(net369),
    .X(_0074_));
 sg13g2_mux2_1 _0753_ (.A0(\i_main_reg.data_d[43] ),
    .A1(net490),
    .S(net354),
    .X(_0075_));
 sg13g2_mux2_1 _0754_ (.A0(net302),
    .A1(net555),
    .S(net354),
    .X(_0076_));
 sg13g2_mux2_1 _0755_ (.A0(\i_main_reg.data_d[45] ),
    .A1(net302),
    .S(net356),
    .X(_0077_));
 sg13g2_mux2_1 _0756_ (.A0(net489),
    .A1(net584),
    .S(net356),
    .X(_0078_));
 sg13g2_mux2_1 _0757_ (.A0(net102),
    .A1(net489),
    .S(net356),
    .X(_0079_));
 sg13g2_mux2_1 _0758_ (.A0(\i_main_reg.data_d[48] ),
    .A1(net102),
    .S(net356),
    .X(_0080_));
 sg13g2_mux2_1 _0759_ (.A0(net527),
    .A1(net674),
    .S(net356),
    .X(_0081_));
 sg13g2_mux2_1 _0760_ (.A0(\i_main_reg.data_d[50] ),
    .A1(net527),
    .S(net356),
    .X(_0082_));
 sg13g2_mux2_1 _0761_ (.A0(\i_main_reg.data_d[51] ),
    .A1(net562),
    .S(net357),
    .X(_0083_));
 sg13g2_mux2_1 _0762_ (.A0(net643),
    .A1(net706),
    .S(net357),
    .X(_0084_));
 sg13g2_mux2_1 _0763_ (.A0(net499),
    .A1(net643),
    .S(net357),
    .X(_0085_));
 sg13g2_mux2_1 _0764_ (.A0(net485),
    .A1(net499),
    .S(net354),
    .X(_0086_));
 sg13g2_mux2_1 _0765_ (.A0(\i_main_reg.data_d[55] ),
    .A1(net485),
    .S(net347),
    .X(_0087_));
 sg13g2_mux2_1 _0766_ (.A0(\i_main_reg.data_d[56] ),
    .A1(net518),
    .S(net347),
    .X(_0088_));
 sg13g2_mux2_1 _0767_ (.A0(net127),
    .A1(net540),
    .S(net348),
    .X(_0089_));
 sg13g2_mux2_1 _0768_ (.A0(\i_main_reg.data_d[58] ),
    .A1(net127),
    .S(net348),
    .X(_0090_));
 sg13g2_mux2_1 _0769_ (.A0(net173),
    .A1(\i_main_reg.data_d[58] ),
    .S(net347),
    .X(_0091_));
 sg13g2_mux2_1 _0770_ (.A0(net218),
    .A1(net173),
    .S(net347),
    .X(_0092_));
 sg13g2_mux2_1 _0771_ (.A0(net155),
    .A1(net218),
    .S(net346),
    .X(_0093_));
 sg13g2_mux2_1 _0772_ (.A0(\i_main_reg.data_d[62] ),
    .A1(net155),
    .S(net346),
    .X(_0094_));
 sg13g2_mux2_1 _0773_ (.A0(net96),
    .A1(net227),
    .S(net346),
    .X(_0095_));
 sg13g2_mux2_1 _0774_ (.A0(\i_main_reg.data_d[64] ),
    .A1(net96),
    .S(net345),
    .X(_0096_));
 sg13g2_mux2_1 _0775_ (.A0(net135),
    .A1(net157),
    .S(net345),
    .X(_0097_));
 sg13g2_mux2_1 _0776_ (.A0(\i_main_reg.data_d[66] ),
    .A1(net135),
    .S(net346),
    .X(_0098_));
 sg13g2_mux2_1 _0777_ (.A0(net66),
    .A1(net481),
    .S(net319),
    .X(_0099_));
 sg13g2_mux2_1 _0778_ (.A0(\i_main_reg.data_d[68] ),
    .A1(net66),
    .S(net319),
    .X(_0100_));
 sg13g2_mux2_1 _0779_ (.A0(net557),
    .A1(net566),
    .S(net320),
    .X(_0101_));
 sg13g2_mux2_1 _0780_ (.A0(net110),
    .A1(net557),
    .S(net320),
    .X(_0102_));
 sg13g2_mux2_1 _0781_ (.A0(\i_main_reg.data_d[71] ),
    .A1(net110),
    .S(net319),
    .X(_0103_));
 sg13g2_mux2_1 _0782_ (.A0(net665),
    .A1(\i_main_reg.data_d[71] ),
    .S(net320),
    .X(_0104_));
 sg13g2_mux2_1 _0783_ (.A0(net522),
    .A1(\i_main_reg.data_d[72] ),
    .S(net319),
    .X(_0105_));
 sg13g2_mux2_1 _0784_ (.A0(net507),
    .A1(net522),
    .S(net319),
    .X(_0106_));
 sg13g2_mux2_1 _0785_ (.A0(net214),
    .A1(net507),
    .S(net317),
    .X(_0107_));
 sg13g2_mux2_1 _0786_ (.A0(\i_main_reg.data_d[76] ),
    .A1(net214),
    .S(net317),
    .X(_0108_));
 sg13g2_mux2_1 _0787_ (.A0(net543),
    .A1(net561),
    .S(net317),
    .X(_0109_));
 sg13g2_mux2_1 _0788_ (.A0(\i_main_reg.data_d[78] ),
    .A1(net543),
    .S(net317),
    .X(_0110_));
 sg13g2_mux2_1 _0789_ (.A0(net690),
    .A1(\i_main_reg.data_d[78] ),
    .S(net309),
    .X(_0111_));
 sg13g2_mux2_1 _0790_ (.A0(net667),
    .A1(\i_main_reg.data_d[79] ),
    .S(net309),
    .X(_0112_));
 sg13g2_mux2_1 _0791_ (.A0(net223),
    .A1(\i_main_reg.data_d[80] ),
    .S(net309),
    .X(_0113_));
 sg13g2_mux2_1 _0792_ (.A0(net471),
    .A1(net223),
    .S(net309),
    .X(_0114_));
 sg13g2_mux2_1 _0793_ (.A0(\i_main_reg.data_d[83] ),
    .A1(net471),
    .S(net309),
    .X(_0115_));
 sg13g2_mux2_1 _0794_ (.A0(net617),
    .A1(\i_main_reg.data_d[83] ),
    .S(net307),
    .X(_0116_));
 sg13g2_mux2_1 _0795_ (.A0(net233),
    .A1(net617),
    .S(net304),
    .X(_0117_));
 sg13g2_mux2_1 _0796_ (.A0(\i_main_reg.data_d[86] ),
    .A1(net233),
    .S(net304),
    .X(_0118_));
 sg13g2_mux2_1 _0797_ (.A0(net500),
    .A1(net724),
    .S(net304),
    .X(_0119_));
 sg13g2_mux2_1 _0798_ (.A0(net158),
    .A1(net500),
    .S(net304),
    .X(_0120_));
 sg13g2_mux2_1 _0799_ (.A0(\i_main_reg.data_d[89] ),
    .A1(net158),
    .S(net306),
    .X(_0121_));
 sg13g2_mux2_1 _0800_ (.A0(\i_main_reg.data_d[90] ),
    .A1(net629),
    .S(net306),
    .X(_0122_));
 sg13g2_mux2_1 _0801_ (.A0(net743),
    .A1(\i_main_reg.data_d[90] ),
    .S(net306),
    .X(_0123_));
 sg13g2_mux2_1 _0802_ (.A0(net704),
    .A1(\i_main_reg.data_d[91] ),
    .S(net306),
    .X(_0124_));
 sg13g2_mux2_1 _0803_ (.A0(net645),
    .A1(net704),
    .S(net313),
    .X(_0125_));
 sg13g2_mux2_1 _0804_ (.A0(net614),
    .A1(net645),
    .S(net313),
    .X(_0126_));
 sg13g2_mux2_1 _0805_ (.A0(net598),
    .A1(net614),
    .S(net313),
    .X(_0127_));
 sg13g2_mux2_1 _0806_ (.A0(\i_main_reg.data_d[96] ),
    .A1(net598),
    .S(net313),
    .X(_0128_));
 sg13g2_mux2_1 _0807_ (.A0(\i_main_reg.data_d[97] ),
    .A1(net707),
    .S(net313),
    .X(_0129_));
 sg13g2_mux2_1 _0808_ (.A0(net730),
    .A1(\i_main_reg.data_d[97] ),
    .S(net315),
    .X(_0130_));
 sg13g2_mux2_1 _0809_ (.A0(net600),
    .A1(\i_main_reg.data_d[98] ),
    .S(net315),
    .X(_0131_));
 sg13g2_mux2_1 _0810_ (.A0(net545),
    .A1(\i_main_reg.data_d[99] ),
    .S(net315),
    .X(_0132_));
 sg13g2_mux2_1 _0811_ (.A0(net501),
    .A1(\i_main_reg.data_d[100] ),
    .S(net315),
    .X(_0133_));
 sg13g2_mux2_1 _0812_ (.A0(net590),
    .A1(net501),
    .S(net315),
    .X(_0134_));
 sg13g2_mux2_1 _0813_ (.A0(net144),
    .A1(net590),
    .S(net314),
    .X(_0135_));
 sg13g2_mux2_1 _0814_ (.A0(net100),
    .A1(net144),
    .S(net319),
    .X(_0136_));
 sg13g2_mux2_1 _0815_ (.A0(\i_main_reg.data_d[105] ),
    .A1(net100),
    .S(net319),
    .X(_0137_));
 sg13g2_mux2_1 _0816_ (.A0(net117),
    .A1(\i_main_reg.data_d[105] ),
    .S(net319),
    .X(_0138_));
 sg13g2_mux2_1 _0817_ (.A0(net243),
    .A1(net117),
    .S(net345),
    .X(_0139_));
 sg13g2_mux2_1 _0818_ (.A0(net210),
    .A1(\i_main_reg.data_d[107] ),
    .S(net345),
    .X(_0140_));
 sg13g2_mux2_1 _0819_ (.A0(net149),
    .A1(net210),
    .S(net345),
    .X(_0141_));
 sg13g2_mux2_1 _0820_ (.A0(\i_main_reg.data_d[110] ),
    .A1(net149),
    .S(net345),
    .X(_0142_));
 sg13g2_mux2_1 _0821_ (.A0(net129),
    .A1(\i_main_reg.data_d[110] ),
    .S(net345),
    .X(_0143_));
 sg13g2_mux2_1 _0822_ (.A0(net535),
    .A1(net129),
    .S(net345),
    .X(_0144_));
 sg13g2_mux2_1 _0823_ (.A0(net235),
    .A1(net535),
    .S(net347),
    .X(_0145_));
 sg13g2_mux2_1 _0824_ (.A0(\i_main_reg.data_d[114] ),
    .A1(net235),
    .S(net347),
    .X(_0146_));
 sg13g2_mux2_1 _0825_ (.A0(net569),
    .A1(net593),
    .S(net347),
    .X(_0147_));
 sg13g2_mux2_1 _0826_ (.A0(net457),
    .A1(net569),
    .S(net347),
    .X(_0148_));
 sg13g2_mux2_1 _0827_ (.A0(net267),
    .A1(net457),
    .S(net354),
    .X(_0149_));
 sg13g2_mux2_1 _0828_ (.A0(\i_main_reg.data_d[118] ),
    .A1(net267),
    .S(net354),
    .X(_0150_));
 sg13g2_mux2_1 _0829_ (.A0(net684),
    .A1(\i_main_reg.data_d[118] ),
    .S(net354),
    .X(_0151_));
 sg13g2_mux2_1 _0830_ (.A0(net192),
    .A1(\i_main_reg.data_d[119] ),
    .S(net354),
    .X(_0152_));
 sg13g2_mux2_1 _0831_ (.A0(net168),
    .A1(net192),
    .S(net354),
    .X(_0153_));
 sg13g2_mux2_1 _0832_ (.A0(\i_main_reg.data_d[122] ),
    .A1(net168),
    .S(net355),
    .X(_0154_));
 sg13g2_mux2_1 _0833_ (.A0(\i_main_reg.data_d[123] ),
    .A1(net530),
    .S(net355),
    .X(_0155_));
 sg13g2_mux2_1 _0834_ (.A0(\i_main_reg.data_d[124] ),
    .A1(net607),
    .S(net355),
    .X(_0156_));
 sg13g2_mux2_1 _0835_ (.A0(net663),
    .A1(\i_main_reg.data_d[124] ),
    .S(net355),
    .X(_0157_));
 sg13g2_mux2_1 _0836_ (.A0(net654),
    .A1(net663),
    .S(net355),
    .X(_0158_));
 sg13g2_mux2_1 _0837_ (.A0(\i_main_reg.data_d[127] ),
    .A1(net654),
    .S(net355),
    .X(_0159_));
 sg13g2_mux2_1 _0838_ (.A0(net657),
    .A1(\i_main_reg.data_d[127] ),
    .S(net355),
    .X(_0160_));
 sg13g2_mux2_1 _0839_ (.A0(net276),
    .A1(\i_main_reg.data_d[128] ),
    .S(net356),
    .X(_0161_));
 sg13g2_mux2_1 _0840_ (.A0(net506),
    .A1(net276),
    .S(net355),
    .X(_0162_));
 sg13g2_mux2_1 _0841_ (.A0(net291),
    .A1(net506),
    .S(net352),
    .X(_0163_));
 sg13g2_mux2_1 _0842_ (.A0(\i_main_reg.data_d[132] ),
    .A1(net291),
    .S(net352),
    .X(_0164_));
 sg13g2_mux2_1 _0843_ (.A0(net611),
    .A1(\i_main_reg.data_d[132] ),
    .S(net352),
    .X(_0165_));
 sg13g2_mux2_1 _0844_ (.A0(net289),
    .A1(\i_main_reg.data_d[133] ),
    .S(net352),
    .X(_0166_));
 sg13g2_mux2_1 _0845_ (.A0(net508),
    .A1(net289),
    .S(net353),
    .X(_0167_));
 sg13g2_mux2_1 _0846_ (.A0(net74),
    .A1(net508),
    .S(net352),
    .X(_0168_));
 sg13g2_mux2_1 _0847_ (.A0(\i_main_reg.data_d[137] ),
    .A1(net74),
    .S(net351),
    .X(_0169_));
 sg13g2_mux2_1 _0848_ (.A0(net138),
    .A1(\i_main_reg.data_d[137] ),
    .S(net351),
    .X(_0170_));
 sg13g2_mux2_1 _0849_ (.A0(net458),
    .A1(net138),
    .S(net353),
    .X(_0171_));
 sg13g2_mux2_1 _0850_ (.A0(\i_main_reg.data_d[140] ),
    .A1(net458),
    .S(net351),
    .X(_0172_));
 sg13g2_mux2_1 _0851_ (.A0(\i_main_reg.data_d[141] ),
    .A1(net727),
    .S(net352),
    .X(_0173_));
 sg13g2_mux2_1 _0852_ (.A0(\i_main_reg.data_d[142] ),
    .A1(net732),
    .S(net352),
    .X(_0174_));
 sg13g2_mux2_1 _0853_ (.A0(net640),
    .A1(\i_main_reg.data_d[142] ),
    .S(net352),
    .X(_0175_));
 sg13g2_mux2_1 _0854_ (.A0(net748),
    .A1(net640),
    .S(net350),
    .X(_0176_));
 sg13g2_mux2_1 _0855_ (.A0(net752),
    .A1(net748),
    .S(net350),
    .X(_0177_));
 sg13g2_mux2_1 _0856_ (.A0(net133),
    .A1(\i_main_reg.data_d[145] ),
    .S(net350),
    .X(_0178_));
 sg13g2_mux2_1 _0857_ (.A0(net76),
    .A1(\i_main_reg.data_d[146] ),
    .S(net350),
    .X(_0179_));
 sg13g2_mux2_1 _0858_ (.A0(net279),
    .A1(net76),
    .S(net350),
    .X(_0180_));
 sg13g2_mux2_1 _0859_ (.A0(\i_main_reg.data_d[149] ),
    .A1(net279),
    .S(net350),
    .X(_0181_));
 sg13g2_mux2_1 _0860_ (.A0(net496),
    .A1(net547),
    .S(net343),
    .X(_0182_));
 sg13g2_mux2_1 _0861_ (.A0(\i_main_reg.data_d[151] ),
    .A1(net496),
    .S(net343),
    .X(_0183_));
 sg13g2_mux2_1 _0862_ (.A0(\i_main_reg.data_d[152] ),
    .A1(net679),
    .S(net343),
    .X(_0184_));
 sg13g2_mux2_1 _0863_ (.A0(net646),
    .A1(\i_main_reg.data_d[152] ),
    .S(net343),
    .X(_0185_));
 sg13g2_mux2_1 _0864_ (.A0(net686),
    .A1(net646),
    .S(net343),
    .X(_0186_));
 sg13g2_mux2_1 _0865_ (.A0(net659),
    .A1(net686),
    .S(net341),
    .X(_0187_));
 sg13g2_mux2_1 _0866_ (.A0(net249),
    .A1(net659),
    .S(net344),
    .X(_0188_));
 sg13g2_mux2_1 _0867_ (.A0(\i_main_reg.data_d[157] ),
    .A1(net249),
    .S(net344),
    .X(_0189_));
 sg13g2_mux2_1 _0868_ (.A0(net247),
    .A1(net521),
    .S(net344),
    .X(_0190_));
 sg13g2_mux2_1 _0869_ (.A0(\i_main_reg.data_d[159] ),
    .A1(net247),
    .S(net343),
    .X(_0191_));
 sg13g2_mux2_1 _0870_ (.A0(\i_main_reg.data_d[160] ),
    .A1(net672),
    .S(net343),
    .X(_0192_));
 sg13g2_mux2_1 _0871_ (.A0(net196),
    .A1(\i_main_reg.data_d[160] ),
    .S(net342),
    .X(_0193_));
 sg13g2_mux2_1 _0872_ (.A0(net468),
    .A1(net196),
    .S(net342),
    .X(_0194_));
 sg13g2_mux2_1 _0873_ (.A0(net594),
    .A1(net468),
    .S(net342),
    .X(_0195_));
 sg13g2_mux2_1 _0874_ (.A0(net70),
    .A1(\i_main_reg.data_d[163] ),
    .S(net342),
    .X(_0196_));
 sg13g2_mux2_1 _0875_ (.A0(net532),
    .A1(net70),
    .S(net342),
    .X(_0197_));
 sg13g2_mux2_1 _0876_ (.A0(net484),
    .A1(net532),
    .S(net349),
    .X(_0198_));
 sg13g2_mux2_1 _0877_ (.A0(net205),
    .A1(net484),
    .S(net349),
    .X(_0199_));
 sg13g2_mux2_1 _0878_ (.A0(net171),
    .A1(net205),
    .S(net349),
    .X(_0200_));
 sg13g2_mux2_1 _0879_ (.A0(\i_main_reg.data_d[169] ),
    .A1(net171),
    .S(net350),
    .X(_0201_));
 sg13g2_mux2_1 _0880_ (.A0(\i_main_reg.data_d[170] ),
    .A1(net541),
    .S(net349),
    .X(_0202_));
 sg13g2_mux2_1 _0881_ (.A0(net464),
    .A1(\i_main_reg.data_d[170] ),
    .S(net351),
    .X(_0203_));
 sg13g2_mux2_1 _0882_ (.A0(net269),
    .A1(\i_main_reg.data_d[171] ),
    .S(net351),
    .X(_0204_));
 sg13g2_mux2_1 _0883_ (.A0(net131),
    .A1(net269),
    .S(net351),
    .X(_0205_));
 sg13g2_mux2_1 _0884_ (.A0(\i_main_reg.data_d[174] ),
    .A1(net131),
    .S(net351),
    .X(_0206_));
 sg13g2_mux2_1 _0885_ (.A0(\i_main_reg.data_d[175] ),
    .A1(net637),
    .S(net351),
    .X(_0207_));
 sg13g2_mux2_1 _0886_ (.A0(net560),
    .A1(net678),
    .S(net349),
    .X(_0208_));
 sg13g2_mux2_1 _0887_ (.A0(net498),
    .A1(net560),
    .S(net349),
    .X(_0209_));
 sg13g2_mux2_1 _0888_ (.A0(net288),
    .A1(net498),
    .S(net349),
    .X(_0210_));
 sg13g2_mux2_1 _0889_ (.A0(net198),
    .A1(net288),
    .S(net349),
    .X(_0211_));
 sg13g2_mux2_1 _0890_ (.A0(\i_main_reg.data_d[180] ),
    .A1(net198),
    .S(net342),
    .X(_0212_));
 sg13g2_mux2_1 _0891_ (.A0(net252),
    .A1(\i_main_reg.data_d[180] ),
    .S(net342),
    .X(_0213_));
 sg13g2_mux2_1 _0892_ (.A0(net274),
    .A1(net252),
    .S(net342),
    .X(_0214_));
 sg13g2_mux2_1 _0893_ (.A0(net165),
    .A1(\i_main_reg.data_d[182] ),
    .S(net341),
    .X(_0215_));
 sg13g2_mux2_1 _0894_ (.A0(net576),
    .A1(net165),
    .S(net341),
    .X(_0216_));
 sg13g2_mux2_1 _0895_ (.A0(net119),
    .A1(\i_main_reg.data_d[184] ),
    .S(net341),
    .X(_0217_));
 sg13g2_mux2_1 _0896_ (.A0(net162),
    .A1(net119),
    .S(net341),
    .X(_0218_));
 sg13g2_mux2_1 _0897_ (.A0(net526),
    .A1(net162),
    .S(net341),
    .X(_0219_));
 sg13g2_mux2_1 _0898_ (.A0(net58),
    .A1(\i_main_reg.data_d[187] ),
    .S(net341),
    .X(_0220_));
 sg13g2_mux2_1 _0899_ (.A0(net160),
    .A1(net58),
    .S(net341),
    .X(_0221_));
 sg13g2_mux2_1 _0900_ (.A0(net121),
    .A1(net160),
    .S(net314),
    .X(_0222_));
 sg13g2_mux2_1 _0901_ (.A0(\i_main_reg.data_d[191] ),
    .A1(net121),
    .S(net314),
    .X(_0223_));
 sg13g2_mux2_1 _0902_ (.A0(\i_main_reg.data_d[192] ),
    .A1(net188),
    .S(net314),
    .X(_0224_));
 sg13g2_mux2_1 _0903_ (.A0(net45),
    .A1(\i_main_reg.data_d[192] ),
    .S(net314),
    .X(_0225_));
 sg13g2_mux2_1 _0904_ (.A0(net161),
    .A1(net45),
    .S(net314),
    .X(_0226_));
 sg13g2_mux2_1 _0905_ (.A0(net271),
    .A1(net161),
    .S(net314),
    .X(_0227_));
 sg13g2_mux2_1 _0906_ (.A0(net503),
    .A1(net271),
    .S(net314),
    .X(_0228_));
 sg13g2_mux2_1 _0907_ (.A0(net570),
    .A1(net503),
    .S(net312),
    .X(_0229_));
 sg13g2_mux2_1 _0908_ (.A0(net278),
    .A1(net570),
    .S(net312),
    .X(_0230_));
 sg13g2_mux2_1 _0909_ (.A0(net212),
    .A1(net278),
    .S(net312),
    .X(_0231_));
 sg13g2_mux2_1 _0910_ (.A0(\i_main_reg.data_d[200] ),
    .A1(net212),
    .S(net312),
    .X(_0232_));
 sg13g2_mux2_1 _0911_ (.A0(\i_main_reg.data_d[201] ),
    .A1(net514),
    .S(net312),
    .X(_0233_));
 sg13g2_mux2_1 _0912_ (.A0(net529),
    .A1(net653),
    .S(net312),
    .X(_0234_));
 sg13g2_mux2_1 _0913_ (.A0(net466),
    .A1(net529),
    .S(net305),
    .X(_0235_));
 sg13g2_mux2_1 _0914_ (.A0(\i_main_reg.data_d[204] ),
    .A1(net466),
    .S(net305),
    .X(_0236_));
 sg13g2_mux2_1 _0915_ (.A0(\i_main_reg.data_d[205] ),
    .A1(net469),
    .S(net305),
    .X(_0237_));
 sg13g2_mux2_1 _0916_ (.A0(net200),
    .A1(\i_main_reg.data_d[205] ),
    .S(net305),
    .X(_0238_));
 sg13g2_mux2_1 _0917_ (.A0(net258),
    .A1(net200),
    .S(net304),
    .X(_0239_));
 sg13g2_mux2_1 _0918_ (.A0(net552),
    .A1(net258),
    .S(net304),
    .X(_0240_));
 sg13g2_mux2_1 _0919_ (.A0(net626),
    .A1(net552),
    .S(net303),
    .X(_0241_));
 sg13g2_mux2_1 _0920_ (.A0(\i_main_reg.data_d[210] ),
    .A1(net626),
    .S(net303),
    .X(_0242_));
 sg13g2_mux2_1 _0921_ (.A0(net231),
    .A1(\i_main_reg.data_d[210] ),
    .S(net303),
    .X(_0243_));
 sg13g2_mux2_1 _0922_ (.A0(net635),
    .A1(net231),
    .S(net303),
    .X(_0244_));
 sg13g2_mux2_1 _0923_ (.A0(net86),
    .A1(\i_main_reg.data_d[212] ),
    .S(net303),
    .X(_0245_));
 sg13g2_mux2_1 _0924_ (.A0(net251),
    .A1(net86),
    .S(net303),
    .X(_0246_));
 sg13g2_mux2_1 _0925_ (.A0(net548),
    .A1(net251),
    .S(net304),
    .X(_0247_));
 sg13g2_mux2_1 _0926_ (.A0(net478),
    .A1(\i_main_reg.data_d[215] ),
    .S(net303),
    .X(_0248_));
 sg13g2_mux2_1 _0927_ (.A0(net176),
    .A1(net478),
    .S(net303),
    .X(_0249_));
 sg13g2_mux2_1 _0928_ (.A0(\i_main_reg.data_d[218] ),
    .A1(net176),
    .S(net305),
    .X(_0250_));
 sg13g2_mux2_1 _0929_ (.A0(net84),
    .A1(\i_main_reg.data_d[218] ),
    .S(net305),
    .X(_0251_));
 sg13g2_mux2_1 _0930_ (.A0(net112),
    .A1(net84),
    .S(net305),
    .X(_0252_));
 sg13g2_mux2_1 _0931_ (.A0(net263),
    .A1(net112),
    .S(net305),
    .X(_0253_));
 sg13g2_mux2_1 _0932_ (.A0(net194),
    .A1(net263),
    .S(net312),
    .X(_0254_));
 sg13g2_mux2_1 _0933_ (.A0(\i_main_reg.data_d[223] ),
    .A1(net194),
    .S(net312),
    .X(_0255_));
 sg13g2_mux2_1 _0934_ (.A0(net244),
    .A1(\i_main_reg.data_d[223] ),
    .S(net313),
    .X(_0256_));
 sg13g2_mux2_1 _0935_ (.A0(net460),
    .A1(net244),
    .S(net313),
    .X(_0257_));
 sg13g2_mux2_1 _0936_ (.A0(\i_main_reg.data_d[226] ),
    .A1(net460),
    .S(net313),
    .X(_0258_));
 sg13g2_mux2_1 _0937_ (.A0(net717),
    .A1(\i_main_reg.data_d[226] ),
    .S(net317),
    .X(_0259_));
 sg13g2_mux2_1 _0938_ (.A0(net696),
    .A1(net717),
    .S(net317),
    .X(_0260_));
 sg13g2_mux2_1 _0939_ (.A0(net636),
    .A1(net696),
    .S(net317),
    .X(_0261_));
 sg13g2_mux2_1 _0940_ (.A0(net551),
    .A1(net636),
    .S(net317),
    .X(_0262_));
 sg13g2_mux2_1 _0941_ (.A0(net145),
    .A1(net551),
    .S(net318),
    .X(_0263_));
 sg13g2_mux2_1 _0942_ (.A0(\i_main_reg.data_d[232] ),
    .A1(net145),
    .S(net318),
    .X(_0264_));
 sg13g2_mux2_1 _0943_ (.A0(net553),
    .A1(\i_main_reg.data_d[232] ),
    .S(net318),
    .X(_0265_));
 sg13g2_mux2_1 _0944_ (.A0(net677),
    .A1(net553),
    .S(net318),
    .X(_0266_));
 sg13g2_mux2_1 _0945_ (.A0(net669),
    .A1(net677),
    .S(net318),
    .X(_0267_));
 sg13g2_mux2_1 _0946_ (.A0(\i_main_reg.data_d[236] ),
    .A1(net669),
    .S(net333),
    .X(_0268_));
 sg13g2_mux2_1 _0947_ (.A0(net681),
    .A1(\i_main_reg.data_d[236] ),
    .S(net334),
    .X(_0269_));
 sg13g2_mux2_1 _0948_ (.A0(net203),
    .A1(\i_main_reg.data_d[237] ),
    .S(net334),
    .X(_0270_));
 sg13g2_mux2_1 _0949_ (.A0(net591),
    .A1(net203),
    .S(net334),
    .X(_0271_));
 sg13g2_mux2_1 _0950_ (.A0(\i_main_reg.data_d[240] ),
    .A1(net591),
    .S(net333),
    .X(_0272_));
 sg13g2_mux2_1 _0951_ (.A0(net572),
    .A1(net648),
    .S(net333),
    .X(_0273_));
 sg13g2_mux2_1 _0952_ (.A0(\i_main_reg.data_d[242] ),
    .A1(net572),
    .S(net333),
    .X(_0274_));
 sg13g2_mux2_1 _0953_ (.A0(net56),
    .A1(\i_main_reg.data_d[242] ),
    .S(net333),
    .X(_0275_));
 sg13g2_mux2_1 _0954_ (.A0(net88),
    .A1(net56),
    .S(net333),
    .X(_0276_));
 sg13g2_mux2_1 _0955_ (.A0(net143),
    .A1(net88),
    .S(net333),
    .X(_0277_));
 sg13g2_mux2_1 _0956_ (.A0(net558),
    .A1(net143),
    .S(net333),
    .X(_0278_));
 sg13g2_mux2_1 _0957_ (.A0(\i_main_reg.data_d[247] ),
    .A1(net558),
    .S(net324),
    .X(_0279_));
 sg13g2_mux2_1 _0958_ (.A0(net208),
    .A1(\i_main_reg.data_d[247] ),
    .S(net324),
    .X(_0280_));
 sg13g2_mux2_1 _0959_ (.A0(net261),
    .A1(net208),
    .S(net309),
    .X(_0281_));
 sg13g2_mux2_1 _0960_ (.A0(net688),
    .A1(net261),
    .S(net309),
    .X(_0282_));
 sg13g2_mux2_1 _0961_ (.A0(net652),
    .A1(net688),
    .S(net310),
    .X(_0283_));
 sg13g2_mux2_1 _0962_ (.A0(net536),
    .A1(net652),
    .S(net310),
    .X(_0284_));
 sg13g2_mux2_1 _0963_ (.A0(\i_main_reg.data_d[253] ),
    .A1(net536),
    .S(net309),
    .X(_0285_));
 sg13g2_mux2_1 _0964_ (.A0(net649),
    .A1(\i_main_reg.data_d[253] ),
    .S(net310),
    .X(_0286_));
 sg13g2_mux2_1 _0965_ (.A0(net206),
    .A1(\i_main_reg.data_d[254] ),
    .S(net308),
    .X(_0287_));
 sg13g2_mux2_1 _0966_ (.A0(net298),
    .A1(net206),
    .S(net308),
    .X(_0288_));
 sg13g2_mux2_1 _0967_ (.A0(net737),
    .A1(net298),
    .S(net307),
    .X(_0289_));
 sg13g2_mux2_1 _0968_ (.A0(net610),
    .A1(net737),
    .S(net307),
    .X(_0290_));
 sg13g2_mux2_1 _0969_ (.A0(net564),
    .A1(net610),
    .S(net307),
    .X(_0291_));
 sg13g2_mux2_1 _0970_ (.A0(\i_main_reg.data_d[260] ),
    .A1(net564),
    .S(net307),
    .X(_0292_));
 sg13g2_mux2_1 _0971_ (.A0(net239),
    .A1(net642),
    .S(net307),
    .X(_0293_));
 sg13g2_mux2_1 _0972_ (.A0(net106),
    .A1(net239),
    .S(net307),
    .X(_0294_));
 sg13g2_mux2_1 _0973_ (.A0(\i_main_reg.data_d[263] ),
    .A1(net106),
    .S(net307),
    .X(_0295_));
 sg13g2_mux2_1 _0974_ (.A0(net178),
    .A1(\i_main_reg.data_d[263] ),
    .S(net308),
    .X(_0296_));
 sg13g2_mux2_1 _0975_ (.A0(net581),
    .A1(net178),
    .S(net308),
    .X(_0297_));
 sg13g2_mux2_1 _0976_ (.A0(net671),
    .A1(net581),
    .S(net308),
    .X(_0298_));
 sg13g2_mux2_1 _0977_ (.A0(net615),
    .A1(\i_main_reg.data_d[266] ),
    .S(net308),
    .X(_0299_));
 sg13g2_mux2_1 _0978_ (.A0(net68),
    .A1(\i_main_reg.data_d[267] ),
    .S(net308),
    .X(_0300_));
 sg13g2_mux2_1 _0979_ (.A0(net473),
    .A1(net68),
    .S(net308),
    .X(_0301_));
 sg13g2_mux2_1 _0980_ (.A0(net281),
    .A1(\i_main_reg.data_d[269] ),
    .S(net321),
    .X(_0302_));
 sg13g2_mux2_1 _0981_ (.A0(net98),
    .A1(net281),
    .S(net321),
    .X(_0303_));
 sg13g2_mux2_1 _0982_ (.A0(\i_main_reg.data_d[272] ),
    .A1(net98),
    .S(net321),
    .X(_0304_));
 sg13g2_mux2_1 _0983_ (.A0(net82),
    .A1(net240),
    .S(net321),
    .X(_0305_));
 sg13g2_mux2_1 _0984_ (.A0(\i_main_reg.data_d[274] ),
    .A1(net82),
    .S(net321),
    .X(_0306_));
 sg13g2_mux2_1 _0985_ (.A0(\i_main_reg.data_d[275] ),
    .A1(net185),
    .S(net321),
    .X(_0307_));
 sg13g2_mux2_1 _0986_ (.A0(\i_main_reg.data_d[276] ),
    .A1(net524),
    .S(net321),
    .X(_0308_));
 sg13g2_mux2_1 _0987_ (.A0(net153),
    .A1(\i_main_reg.data_d[276] ),
    .S(net322),
    .X(_0309_));
 sg13g2_mux2_1 _0988_ (.A0(net549),
    .A1(net153),
    .S(net322),
    .X(_0310_));
 sg13g2_mux2_1 _0989_ (.A0(net482),
    .A1(\i_main_reg.data_d[278] ),
    .S(net322),
    .X(_0311_));
 sg13g2_mux2_1 _0990_ (.A0(net589),
    .A1(net482),
    .S(net323),
    .X(_0312_));
 sg13g2_mux2_1 _0991_ (.A0(net662),
    .A1(net589),
    .S(net323),
    .X(_0313_));
 sg13g2_mux2_1 _0992_ (.A0(net462),
    .A1(\i_main_reg.data_d[281] ),
    .S(net321),
    .X(_0314_));
 sg13g2_mux2_1 _0993_ (.A0(net221),
    .A1(net462),
    .S(net324),
    .X(_0315_));
 sg13g2_mux2_1 _0994_ (.A0(\i_main_reg.data_d[284] ),
    .A1(net221),
    .S(net324),
    .X(_0316_));
 sg13g2_mux2_1 _0995_ (.A0(net246),
    .A1(net299),
    .S(net324),
    .X(_0317_));
 sg13g2_mux2_1 _0996_ (.A0(net142),
    .A1(net246),
    .S(net324),
    .X(_0318_));
 sg13g2_mux2_1 _0997_ (.A0(net115),
    .A1(net142),
    .S(net325),
    .X(_0319_));
 sg13g2_mux2_1 _0998_ (.A0(\i_main_reg.data_d[288] ),
    .A1(net115),
    .S(net325),
    .X(_0320_));
 sg13g2_mux2_1 _0999_ (.A0(net60),
    .A1(\i_main_reg.data_d[288] ),
    .S(net325),
    .X(_0321_));
 sg13g2_mux2_1 _1000_ (.A0(net170),
    .A1(net60),
    .S(net325),
    .X(_0322_));
 sg13g2_mux2_1 _1001_ (.A0(net579),
    .A1(net170),
    .S(net324),
    .X(_0323_));
 sg13g2_mux2_1 _1002_ (.A0(net639),
    .A1(net579),
    .S(net324),
    .X(_0324_));
 sg13g2_mux2_1 _1003_ (.A0(net644),
    .A1(net639),
    .S(net330),
    .X(_0325_));
 sg13g2_mux2_1 _1004_ (.A0(net757),
    .A1(net644),
    .S(net330),
    .X(_0326_));
 sg13g2_mux2_1 _1005_ (.A0(net585),
    .A1(\i_main_reg.data_d[294] ),
    .S(net330),
    .X(_0327_));
 sg13g2_mux2_1 _1006_ (.A0(net722),
    .A1(net585),
    .S(net330),
    .X(_0328_));
 sg13g2_mux2_1 _1007_ (.A0(\i_main_reg.data_d[297] ),
    .A1(net722),
    .S(net330),
    .X(_0329_));
 sg13g2_mux2_1 _1008_ (.A0(net689),
    .A1(net738),
    .S(net322),
    .X(_0330_));
 sg13g2_mux2_1 _1009_ (.A0(net474),
    .A1(net689),
    .S(net323),
    .X(_0331_));
 sg13g2_mux2_1 _1010_ (.A0(\i_main_reg.data_d[300] ),
    .A1(net474),
    .S(net322),
    .X(_0332_));
 sg13g2_mux2_1 _1011_ (.A0(\i_main_reg.data_d[301] ),
    .A1(net735),
    .S(net322),
    .X(_0333_));
 sg13g2_mux2_1 _1012_ (.A0(net633),
    .A1(\i_main_reg.data_d[301] ),
    .S(net322),
    .X(_0334_));
 sg13g2_mux2_1 _1013_ (.A0(net687),
    .A1(net633),
    .S(net322),
    .X(_0335_));
 sg13g2_mux2_1 _1014_ (.A0(net125),
    .A1(\i_main_reg.data_d[303] ),
    .S(net328),
    .X(_0336_));
 sg13g2_mux2_1 _1015_ (.A0(net202),
    .A1(net125),
    .S(net328),
    .X(_0337_));
 sg13g2_mux2_1 _1016_ (.A0(net295),
    .A1(net202),
    .S(net328),
    .X(_0338_));
 sg13g2_mux2_1 _1017_ (.A0(net625),
    .A1(net295),
    .S(net328),
    .X(_0339_));
 sg13g2_mux2_1 _1018_ (.A0(net656),
    .A1(net625),
    .S(net328),
    .X(_0340_));
 sg13g2_mux2_1 _1019_ (.A0(net123),
    .A1(\i_main_reg.data_d[308] ),
    .S(net328),
    .X(_0341_));
 sg13g2_mux2_1 _1020_ (.A0(net533),
    .A1(net123),
    .S(net328),
    .X(_0342_));
 sg13g2_mux2_1 _1021_ (.A0(net574),
    .A1(net533),
    .S(net326),
    .X(_0343_));
 sg13g2_mux2_1 _1022_ (.A0(net567),
    .A1(\i_main_reg.data_d[311] ),
    .S(net326),
    .X(_0344_));
 sg13g2_mux2_1 _1023_ (.A0(net516),
    .A1(\i_main_reg.data_d[312] ),
    .S(net326),
    .X(_0345_));
 sg13g2_mux2_1 _1024_ (.A0(net556),
    .A1(net516),
    .S(net326),
    .X(_0346_));
 sg13g2_mux2_1 _1025_ (.A0(net661),
    .A1(net556),
    .S(net327),
    .X(_0347_));
 sg13g2_mux2_1 _1026_ (.A0(net602),
    .A1(\i_main_reg.data_d[315] ),
    .S(net326),
    .X(_0348_));
 sg13g2_mux2_1 _1027_ (.A0(net604),
    .A1(net602),
    .S(net326),
    .X(_0349_));
 sg13g2_mux2_1 _1028_ (.A0(\i_main_reg.data_d[318] ),
    .A1(net604),
    .S(net326),
    .X(_0350_));
 sg13g2_mux2_1 _1029_ (.A0(\i_main_reg.data_d[319] ),
    .A1(net713),
    .S(net326),
    .X(_0351_));
 sg13g2_mux2_1 _1030_ (.A0(net492),
    .A1(\i_main_reg.data_d[319] ),
    .S(net327),
    .X(_0352_));
 sg13g2_mux2_1 _1031_ (.A0(net651),
    .A1(net492),
    .S(net327),
    .X(_0353_));
 sg13g2_mux2_1 _1032_ (.A0(net512),
    .A1(net651),
    .S(net327),
    .X(_0354_));
 sg13g2_mux2_1 _1033_ (.A0(\i_main_reg.data_d[323] ),
    .A1(net512),
    .S(net327),
    .X(_0355_));
 sg13g2_mux2_1 _1034_ (.A0(net219),
    .A1(net580),
    .S(net329),
    .X(_0356_));
 sg13g2_mux2_1 _1035_ (.A0(\i_main_reg.data_d[325] ),
    .A1(net219),
    .S(net329),
    .X(_0357_));
 sg13g2_mux2_1 _1036_ (.A0(\i_main_reg.data_d[326] ),
    .A1(net619),
    .S(net329),
    .X(_0358_));
 sg13g2_mux2_1 _1037_ (.A0(net52),
    .A1(\i_main_reg.data_d[326] ),
    .S(net329),
    .X(_0359_));
 sg13g2_mux2_1 _1038_ (.A0(net181),
    .A1(net52),
    .S(net329),
    .X(_0360_));
 sg13g2_mux2_1 _1039_ (.A0(net94),
    .A1(net181),
    .S(net329),
    .X(_0361_));
 sg13g2_mux2_1 _1040_ (.A0(\i_main_reg.data_d[330] ),
    .A1(net94),
    .S(net329),
    .X(_0362_));
 sg13g2_mux2_1 _1041_ (.A0(\i_main_reg.data_d[331] ),
    .A1(net225),
    .S(net329),
    .X(_0363_));
 sg13g2_mux2_1 _1042_ (.A0(net54),
    .A1(\i_main_reg.data_d[331] ),
    .S(net330),
    .X(_0364_));
 sg13g2_mux2_1 _1043_ (.A0(net187),
    .A1(net54),
    .S(net330),
    .X(_0365_));
 sg13g2_mux2_1 _1044_ (.A0(net550),
    .A1(net187),
    .S(net331),
    .X(_0366_));
 sg13g2_mux2_1 _1045_ (.A0(net575),
    .A1(net550),
    .S(net331),
    .X(_0367_));
 sg13g2_mux2_1 _1046_ (.A0(net216),
    .A1(net575),
    .S(net337),
    .X(_0368_));
 sg13g2_mux2_1 _1047_ (.A0(\i_main_reg.data_d[337] ),
    .A1(net216),
    .S(net337),
    .X(_0369_));
 sg13g2_mux2_1 _1048_ (.A0(net64),
    .A1(\i_main_reg.data_d[337] ),
    .S(net337),
    .X(_0370_));
 sg13g2_mux2_1 _1049_ (.A0(net180),
    .A1(net64),
    .S(net337),
    .X(_0371_));
 sg13g2_mux2_1 _1050_ (.A0(net147),
    .A1(\i_main_reg.data_d[339] ),
    .S(net336),
    .X(_0372_));
 sg13g2_mux2_1 _1051_ (.A0(net167),
    .A1(net147),
    .S(net336),
    .X(_0373_));
 sg13g2_mux2_1 _1052_ (.A0(net510),
    .A1(net167),
    .S(net336),
    .X(_0374_));
 sg13g2_mux2_1 _1053_ (.A0(\i_main_reg.data_d[343] ),
    .A1(net510),
    .S(net337),
    .X(_0375_));
 sg13g2_mux2_1 _1054_ (.A0(net595),
    .A1(net660),
    .S(net339),
    .X(_0376_));
 sg13g2_mux2_1 _1055_ (.A0(net228),
    .A1(net595),
    .S(net339),
    .X(_0377_));
 sg13g2_mux2_1 _1056_ (.A0(\i_main_reg.data_d[346] ),
    .A1(net228),
    .S(net336),
    .X(_0378_));
 sg13g2_mux2_1 _1057_ (.A0(net597),
    .A1(net703),
    .S(net336),
    .X(_0379_));
 sg13g2_mux2_1 _1058_ (.A0(net108),
    .A1(net597),
    .S(net336),
    .X(_0380_));
 sg13g2_mux2_1 _1059_ (.A0(\i_main_reg.data_d[349] ),
    .A1(net108),
    .S(net336),
    .X(_0381_));
 sg13g2_mux2_1 _1060_ (.A0(net259),
    .A1(net287),
    .S(net336),
    .X(_0382_));
 sg13g2_mux2_1 _1061_ (.A0(\i_main_reg.data_d[351] ),
    .A1(net259),
    .S(net335),
    .X(_0383_));
 sg13g2_mux2_1 _1062_ (.A0(net72),
    .A1(\i_main_reg.data_d[351] ),
    .S(net334),
    .X(_0384_));
 sg13g2_mux2_1 _1063_ (.A0(net571),
    .A1(net72),
    .S(net334),
    .X(_0385_));
 sg13g2_mux2_1 _1064_ (.A0(net140),
    .A1(\i_main_reg.data_d[353] ),
    .S(net334),
    .X(_0386_));
 sg13g2_mux2_1 _1065_ (.A0(net296),
    .A1(net140),
    .S(net338),
    .X(_0387_));
 sg13g2_mux2_1 _1066_ (.A0(\i_main_reg.data_d[356] ),
    .A1(net296),
    .S(net338),
    .X(_0388_));
 sg13g2_mux2_1 _1067_ (.A0(net285),
    .A1(\i_main_reg.data_d[356] ),
    .S(net338),
    .X(_0389_));
 sg13g2_mux2_1 _1068_ (.A0(net78),
    .A1(net285),
    .S(net338),
    .X(_0390_));
 sg13g2_mux2_1 _1069_ (.A0(\i_main_reg.data_d[359] ),
    .A1(net78),
    .S(net338),
    .X(_0391_));
 sg13g2_mux2_1 _1070_ (.A0(\i_main_reg.data_d[360] ),
    .A1(net623),
    .S(net338),
    .X(_0392_));
 sg13g2_mux2_1 _1071_ (.A0(\i_main_reg.data_d[361] ),
    .A1(net711),
    .S(net338),
    .X(_0393_));
 sg13g2_mux2_1 _1072_ (.A0(net701),
    .A1(\i_main_reg.data_d[361] ),
    .S(net338),
    .X(_0394_));
 sg13g2_mux2_1 _1073_ (.A0(net621),
    .A1(\i_main_reg.data_d[362] ),
    .S(net365),
    .X(_0395_));
 sg13g2_mux2_1 _1074_ (.A0(net163),
    .A1(\i_main_reg.data_d[363] ),
    .S(net365),
    .X(_0396_));
 sg13g2_mux2_1 _1075_ (.A0(net275),
    .A1(net163),
    .S(net365),
    .X(_0397_));
 sg13g2_mux2_1 _1076_ (.A0(net262),
    .A1(net275),
    .S(net365),
    .X(_0398_));
 sg13g2_mux2_1 _1077_ (.A0(net256),
    .A1(net262),
    .S(net365),
    .X(_0399_));
 sg13g2_mux2_1 _1078_ (.A0(\i_main_reg.data_d[368] ),
    .A1(net256),
    .S(net364),
    .X(_0400_));
 sg13g2_mux2_1 _1079_ (.A0(net456),
    .A1(net480),
    .S(net364),
    .X(_0401_));
 sg13g2_mux2_1 _1080_ (.A0(net190),
    .A1(net456),
    .S(net364),
    .X(_0402_));
 sg13g2_mux2_1 _1081_ (.A0(\i_main_reg.data_d[371] ),
    .A1(net190),
    .S(net367),
    .X(_0403_));
 sg13g2_mux2_1 _1082_ (.A0(net628),
    .A1(net751),
    .S(net367),
    .X(_0404_));
 sg13g2_mux2_1 _1083_ (.A0(net520),
    .A1(net628),
    .S(net366),
    .X(_0405_));
 sg13g2_mux2_1 _1084_ (.A0(net293),
    .A1(net520),
    .S(net366),
    .X(_0406_));
 sg13g2_mux2_1 _1085_ (.A0(\i_main_reg.data_d[375] ),
    .A1(net293),
    .S(net366),
    .X(_0407_));
 sg13g2_mux2_1 _1086_ (.A0(\i_main_reg.data_d[376] ),
    .A1(net538),
    .S(net366),
    .X(_0408_));
 sg13g2_mux2_1 _1087_ (.A0(net487),
    .A1(\i_main_reg.data_d[376] ),
    .S(net366),
    .X(_0409_));
 sg13g2_mux2_1 _1088_ (.A0(net80),
    .A1(net487),
    .S(net368),
    .X(_0410_));
 sg13g2_mux2_1 _1089_ (.A0(\i_main_reg.data_d[379] ),
    .A1(net80),
    .S(net368),
    .X(_0411_));
 sg13g2_mux2_1 _1090_ (.A0(net62),
    .A1(\i_main_reg.data_d[379] ),
    .S(net368),
    .X(_0412_));
 sg13g2_mux2_1 _1091_ (.A0(net137),
    .A1(net62),
    .S(net368),
    .X(_0413_));
 sg13g2_mux2_1 _1092_ (.A0(net92),
    .A1(\i_main_reg.data_d[381] ),
    .S(net369),
    .X(_0414_));
 sg13g2_xor2_1 _1093_ (.B(previous_bit_q),
    .A(net378),
    .X(_0418_));
 sg13g2_xnor2_1 _1094_ (.Y(_0419_),
    .A(net264),
    .B(_0418_));
 sg13g2_o21ai_1 _1095_ (.B1(_0440_),
    .Y(_0420_),
    .A1(net378),
    .A2(_0443_));
 sg13g2_o21ai_1 _1096_ (.B1(_0420_),
    .Y(_0421_),
    .A1(_0520_),
    .A2(_0419_));
 sg13g2_and4_1 _1097_ (.A(net2),
    .B(net1),
    .C(_0519_),
    .D(_0530_),
    .X(_0422_));
 sg13g2_a221oi_1 _1098_ (.B2(_0529_),
    .C1(_0422_),
    .B1(net762),
    .A1(net92),
    .Y(_0423_),
    .A2(net369));
 sg13g2_inv_1 _1099_ (.Y(_0415_),
    .A(_0423_));
 sg13g2_nand2_1 _1100_ (.Y(_0424_),
    .A(net753),
    .B(net31));
 sg13g2_o21ai_1 _1101_ (.B1(_0440_),
    .Y(_0425_),
    .A1(net379),
    .A2(_0442_));
 sg13g2_a21oi_1 _1102_ (.A1(net379),
    .A2(_0424_),
    .Y(_0426_),
    .B1(_0425_));
 sg13g2_or4_1 _1103_ (.A(_0514_),
    .B(_0521_),
    .C(_0550_),
    .D(_0426_),
    .X(_0427_));
 sg13g2_nand2_1 _1104_ (.Y(_0428_),
    .A(net31),
    .B(_0427_));
 sg13g2_nand4_1 _1105_ (.B(_0513_),
    .C(_0031_),
    .A(net379),
    .Y(_0429_),
    .D(_0424_));
 sg13g2_o21ai_1 _1106_ (.B1(_0428_),
    .Y(_0416_),
    .A1(net31),
    .A2(_0429_));
 sg13g2_nand2_1 _1107_ (.Y(_0430_),
    .A(net753),
    .B(_0427_));
 sg13g2_nand2b_1 _1108_ (.Y(_0431_),
    .B(_0424_),
    .A_N(_0445_));
 sg13g2_o21ai_1 _1109_ (.B1(_0430_),
    .Y(_0417_),
    .A1(_0429_),
    .A2(_0431_));
 sg13g2_dfrbpq_2 _1110_ (.RESET_B(net445),
    .D(net710),
    .Q(\i_step_counter.data_o ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1111_ (.RESET_B(net445),
    .D(net765),
    .Q(\i_step_counter.data_d[0] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1112_ (.RESET_B(net445),
    .D(net726),
    .Q(\i_step_counter.data_d[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1113_ (.RESET_B(net445),
    .D(_0003_),
    .Q(\i_step_counter.data_d[2] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1114_ (.RESET_B(net445),
    .D(net35),
    .Q(\i_step_counter.data_d[3] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1115_ (.RESET_B(net445),
    .D(_0005_),
    .Q(\i_step_counter.data_d[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1116_ (.RESET_B(net445),
    .D(net42),
    .Q(\i_step_counter.data_d[5] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _1117_ (.RESET_B(net445),
    .D(_0007_),
    .Q(\i_step_counter.data_d[6] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _1118_ (.RESET_B(net447),
    .D(_0008_),
    .Q(\i_step_counter.data_d[7] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1119_ (.RESET_B(net447),
    .D(_0009_),
    .Q(\i_step_counter.data_d[8] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1120_ (.RESET_B(net447),
    .D(net768),
    .Q(\i_step_counter.data_d[9] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1121_ (.RESET_B(net447),
    .D(net742),
    .Q(\i_step_counter.data_d[10] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _1122_ (.RESET_B(net446),
    .D(net776),
    .Q(\i_step_counter.data_d[11] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1123_ (.RESET_B(net446),
    .D(net721),
    .Q(\i_step_counter.data_d[12] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1124_ (.RESET_B(net446),
    .D(net756),
    .Q(\i_step_counter.data_d[13] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1125_ (.RESET_B(net446),
    .D(net184),
    .Q(\i_step_counter.data_d[14] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1126_ (.RESET_B(net446),
    .D(net38),
    .Q(finished_q),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1127_ (.RESET_B(net446),
    .D(net27),
    .Q(overflow_q),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1128_ (.RESET_B(net449),
    .D(net266),
    .Q(carry_q),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1129_ (.RESET_B(net449),
    .D(_0019_),
    .Q(previous_bit_q),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _1130_ (.RESET_B(net448),
    .D(_0020_),
    .Q(\bit_counter_q[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1131_ (.RESET_B(net451),
    .D(net49),
    .Q(\bit_counter_q[1] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1132_ (.RESET_B(net448),
    .D(_0022_),
    .Q(\bit_counter_q[2] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1133_ (.RESET_B(net448),
    .D(net91),
    .Q(\bit_counter_q[3] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1134_ (.RESET_B(net451),
    .D(net30),
    .Q(\bit_counter_q[4] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1135_ (.RESET_B(net448),
    .D(_0025_),
    .Q(\bit_counter_q[5] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1136_ (.RESET_B(net448),
    .D(_0026_),
    .Q(\bit_counter_q[6] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_2 _1137_ (.RESET_B(net448),
    .D(net747),
    .Q(\bit_counter_q[7] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1138_ (.RESET_B(net448),
    .D(net716),
    .Q(\bit_counter_q[8] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _1139_ (.RESET_B(net449),
    .D(_0029_),
    .Q(\bit_counter_q[9] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1140_ (.RESET_B(net449),
    .D(_0030_),
    .Q(\state_q[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _1141_ (.RESET_B(net449),
    .D(_0031_),
    .Q(\state_q[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _1142_ (.RESET_B(net449),
    .D(_0032_),
    .Q(\i_main_reg.data_o ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1143_ (.RESET_B(net450),
    .D(_0033_),
    .Q(\i_main_reg.data_d[0] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1144_ (.RESET_B(net450),
    .D(net242),
    .Q(\i_main_reg.data_d[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1145_ (.RESET_B(net450),
    .D(net301),
    .Q(\i_main_reg.data_d[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1146_ (.RESET_B(net443),
    .D(_0036_),
    .Q(\i_main_reg.data_d[3] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1147_ (.RESET_B(net443),
    .D(net676),
    .Q(\i_main_reg.data_d[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1148_ (.RESET_B(net443),
    .D(_0038_),
    .Q(\i_main_reg.data_d[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1149_ (.RESET_B(net443),
    .D(net698),
    .Q(\i_main_reg.data_d[6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1150_ (.RESET_B(net440),
    .D(net700),
    .Q(\i_main_reg.data_d[7] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1151_ (.RESET_B(net440),
    .D(_0041_),
    .Q(\i_main_reg.data_d[8] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1152_ (.RESET_B(net440),
    .D(net477),
    .Q(\i_main_reg.data_d[9] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1153_ (.RESET_B(net438),
    .D(_0043_),
    .Q(\i_main_reg.data_d[10] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1154_ (.RESET_B(net438),
    .D(_0044_),
    .Q(\i_main_reg.data_d[11] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1155_ (.RESET_B(net441),
    .D(_0045_),
    .Q(\i_main_reg.data_d[12] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1156_ (.RESET_B(net441),
    .D(_0046_),
    .Q(\i_main_reg.data_d[13] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1157_ (.RESET_B(net441),
    .D(net495),
    .Q(\i_main_reg.data_d[14] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1158_ (.RESET_B(net441),
    .D(net583),
    .Q(\i_main_reg.data_d[15] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1159_ (.RESET_B(net441),
    .D(_0049_),
    .Q(\i_main_reg.data_d[16] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1160_ (.RESET_B(net440),
    .D(_0050_),
    .Q(\i_main_reg.data_d[17] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1161_ (.RESET_B(net440),
    .D(net284),
    .Q(\i_main_reg.data_d[18] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1162_ (.RESET_B(net440),
    .D(net588),
    .Q(\i_main_reg.data_d[19] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1163_ (.RESET_B(net414),
    .D(net51),
    .Q(\i_main_reg.data_d[20] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1164_ (.RESET_B(net414),
    .D(_0054_),
    .Q(\i_main_reg.data_d[21] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1165_ (.RESET_B(net413),
    .D(net238),
    .Q(\i_main_reg.data_d[22] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1166_ (.RESET_B(net413),
    .D(net505),
    .Q(\i_main_reg.data_d[23] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1167_ (.RESET_B(net413),
    .D(net105),
    .Q(\i_main_reg.data_d[24] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1168_ (.RESET_B(net413),
    .D(_0058_),
    .Q(\i_main_reg.data_d[25] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1169_ (.RESET_B(net413),
    .D(_0059_),
    .Q(\i_main_reg.data_d[26] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1170_ (.RESET_B(net438),
    .D(net114),
    .Q(\i_main_reg.data_d[27] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1171_ (.RESET_B(net438),
    .D(net273),
    .Q(\i_main_reg.data_d[28] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1172_ (.RESET_B(net438),
    .D(net152),
    .Q(\i_main_reg.data_d[29] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1173_ (.RESET_B(net438),
    .D(_0063_),
    .Q(\i_main_reg.data_d[30] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1174_ (.RESET_B(net438),
    .D(_0064_),
    .Q(\i_main_reg.data_d[31] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1175_ (.RESET_B(net438),
    .D(net632),
    .Q(\i_main_reg.data_d[32] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1176_ (.RESET_B(net439),
    .D(_0066_),
    .Q(\i_main_reg.data_d[33] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1177_ (.RESET_B(net439),
    .D(net455),
    .Q(\i_main_reg.data_d[34] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1178_ (.RESET_B(net439),
    .D(_0068_),
    .Q(\i_main_reg.data_d[35] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1179_ (.RESET_B(net439),
    .D(_0069_),
    .Q(\i_main_reg.data_d[36] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1180_ (.RESET_B(net439),
    .D(net578),
    .Q(\i_main_reg.data_d[37] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1181_ (.RESET_B(net439),
    .D(net695),
    .Q(\i_main_reg.data_d[38] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _1182_ (.RESET_B(net439),
    .D(_0072_),
    .Q(\i_main_reg.data_d[39] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1183_ (.RESET_B(net439),
    .D(_0073_),
    .Q(\i_main_reg.data_d[40] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _1184_ (.RESET_B(net447),
    .D(net255),
    .Q(\i_main_reg.data_d[41] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1185_ (.RESET_B(net447),
    .D(net491),
    .Q(\i_main_reg.data_d[42] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1186_ (.RESET_B(net434),
    .D(_0076_),
    .Q(\i_main_reg.data_d[43] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1187_ (.RESET_B(net434),
    .D(net453),
    .Q(\i_main_reg.data_d[44] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1188_ (.RESET_B(net434),
    .D(_0078_),
    .Q(\i_main_reg.data_d[45] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1189_ (.RESET_B(net437),
    .D(_0079_),
    .Q(\i_main_reg.data_d[46] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1190_ (.RESET_B(net437),
    .D(net103),
    .Q(\i_main_reg.data_d[47] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1191_ (.RESET_B(net437),
    .D(_0081_),
    .Q(\i_main_reg.data_d[48] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1192_ (.RESET_B(net435),
    .D(net528),
    .Q(\i_main_reg.data_d[49] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1193_ (.RESET_B(net435),
    .D(net563),
    .Q(\i_main_reg.data_d[50] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1194_ (.RESET_B(net435),
    .D(_0084_),
    .Q(\i_main_reg.data_d[51] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1195_ (.RESET_B(net435),
    .D(_0085_),
    .Q(\i_main_reg.data_d[52] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _1196_ (.RESET_B(net427),
    .D(_0086_),
    .Q(\i_main_reg.data_d[53] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1197_ (.RESET_B(net426),
    .D(net486),
    .Q(\i_main_reg.data_d[54] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1198_ (.RESET_B(net426),
    .D(net519),
    .Q(\i_main_reg.data_d[55] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1199_ (.RESET_B(net426),
    .D(_0089_),
    .Q(\i_main_reg.data_d[56] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1200_ (.RESET_B(net426),
    .D(net128),
    .Q(\i_main_reg.data_d[57] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1201_ (.RESET_B(net427),
    .D(net174),
    .Q(\i_main_reg.data_d[58] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1202_ (.RESET_B(net424),
    .D(_0092_),
    .Q(\i_main_reg.data_d[59] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1203_ (.RESET_B(net424),
    .D(_0093_),
    .Q(\i_main_reg.data_d[60] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1204_ (.RESET_B(net425),
    .D(net156),
    .Q(\i_main_reg.data_d[61] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1205_ (.RESET_B(net425),
    .D(_0095_),
    .Q(\i_main_reg.data_d[62] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _1206_ (.RESET_B(net425),
    .D(net97),
    .Q(\i_main_reg.data_d[63] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1207_ (.RESET_B(net425),
    .D(_0097_),
    .Q(\i_main_reg.data_d[64] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1208_ (.RESET_B(net425),
    .D(net136),
    .Q(\i_main_reg.data_d[65] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1209_ (.RESET_B(net397),
    .D(_0099_),
    .Q(\i_main_reg.data_d[66] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1210_ (.RESET_B(net397),
    .D(net67),
    .Q(\i_main_reg.data_d[67] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1211_ (.RESET_B(net398),
    .D(_0101_),
    .Q(\i_main_reg.data_d[68] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _1212_ (.RESET_B(net398),
    .D(_0102_),
    .Q(\i_main_reg.data_d[69] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1213_ (.RESET_B(net397),
    .D(net111),
    .Q(\i_main_reg.data_d[70] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1214_ (.RESET_B(net398),
    .D(net666),
    .Q(\i_main_reg.data_d[71] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1215_ (.RESET_B(net397),
    .D(net523),
    .Q(\i_main_reg.data_d[72] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1216_ (.RESET_B(net395),
    .D(_0106_),
    .Q(\i_main_reg.data_d[73] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1217_ (.RESET_B(net395),
    .D(_0107_),
    .Q(\i_main_reg.data_d[74] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1218_ (.RESET_B(net395),
    .D(net215),
    .Q(\i_main_reg.data_d[75] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1219_ (.RESET_B(net395),
    .D(_0109_),
    .Q(\i_main_reg.data_d[76] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1220_ (.RESET_B(net395),
    .D(net544),
    .Q(\i_main_reg.data_d[77] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1221_ (.RESET_B(net387),
    .D(net691),
    .Q(\i_main_reg.data_d[78] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1222_ (.RESET_B(net387),
    .D(net668),
    .Q(\i_main_reg.data_d[79] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1223_ (.RESET_B(net387),
    .D(net224),
    .Q(\i_main_reg.data_d[80] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1224_ (.RESET_B(net387),
    .D(_0114_),
    .Q(\i_main_reg.data_d[81] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1225_ (.RESET_B(net387),
    .D(net472),
    .Q(\i_main_reg.data_d[82] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1226_ (.RESET_B(net386),
    .D(net618),
    .Q(\i_main_reg.data_d[83] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1227_ (.RESET_B(net381),
    .D(_0117_),
    .Q(\i_main_reg.data_d[84] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1228_ (.RESET_B(net381),
    .D(net234),
    .Q(\i_main_reg.data_d[85] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1229_ (.RESET_B(net381),
    .D(_0119_),
    .Q(\i_main_reg.data_d[86] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1230_ (.RESET_B(net389),
    .D(_0120_),
    .Q(\i_main_reg.data_d[87] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1231_ (.RESET_B(net381),
    .D(net159),
    .Q(\i_main_reg.data_d[88] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1232_ (.RESET_B(net383),
    .D(net630),
    .Q(\i_main_reg.data_d[89] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1233_ (.RESET_B(net383),
    .D(net744),
    .Q(\i_main_reg.data_d[90] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1234_ (.RESET_B(net383),
    .D(net705),
    .Q(\i_main_reg.data_d[91] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1235_ (.RESET_B(net383),
    .D(_0125_),
    .Q(\i_main_reg.data_d[92] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1236_ (.RESET_B(net391),
    .D(_0126_),
    .Q(\i_main_reg.data_d[93] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1237_ (.RESET_B(net391),
    .D(_0127_),
    .Q(\i_main_reg.data_d[94] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1238_ (.RESET_B(net391),
    .D(net599),
    .Q(\i_main_reg.data_d[95] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1239_ (.RESET_B(net391),
    .D(net708),
    .Q(\i_main_reg.data_d[96] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1240_ (.RESET_B(net391),
    .D(net731),
    .Q(\i_main_reg.data_d[97] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1241_ (.RESET_B(net393),
    .D(net601),
    .Q(\i_main_reg.data_d[98] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1242_ (.RESET_B(net393),
    .D(net546),
    .Q(\i_main_reg.data_d[99] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1243_ (.RESET_B(net393),
    .D(net502),
    .Q(\i_main_reg.data_d[100] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1244_ (.RESET_B(net393),
    .D(_0134_),
    .Q(\i_main_reg.data_d[101] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1245_ (.RESET_B(net393),
    .D(_0135_),
    .Q(\i_main_reg.data_d[102] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1246_ (.RESET_B(net397),
    .D(_0136_),
    .Q(\i_main_reg.data_d[103] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1247_ (.RESET_B(net397),
    .D(net101),
    .Q(\i_main_reg.data_d[104] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1248_ (.RESET_B(net397),
    .D(net118),
    .Q(\i_main_reg.data_d[105] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1249_ (.RESET_B(net397),
    .D(_0139_),
    .Q(\i_main_reg.data_d[106] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1250_ (.RESET_B(net424),
    .D(net211),
    .Q(\i_main_reg.data_d[107] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1251_ (.RESET_B(net424),
    .D(_0141_),
    .Q(\i_main_reg.data_d[108] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1252_ (.RESET_B(net424),
    .D(net150),
    .Q(\i_main_reg.data_d[109] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _1253_ (.RESET_B(net424),
    .D(net130),
    .Q(\i_main_reg.data_d[110] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1254_ (.RESET_B(net424),
    .D(_0144_),
    .Q(\i_main_reg.data_d[111] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1255_ (.RESET_B(net424),
    .D(_0145_),
    .Q(\i_main_reg.data_d[112] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1256_ (.RESET_B(net426),
    .D(net236),
    .Q(\i_main_reg.data_d[113] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1257_ (.RESET_B(net426),
    .D(_0147_),
    .Q(\i_main_reg.data_d[114] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1258_ (.RESET_B(net426),
    .D(_0148_),
    .Q(\i_main_reg.data_d[115] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1259_ (.RESET_B(net426),
    .D(_0149_),
    .Q(\i_main_reg.data_d[116] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1260_ (.RESET_B(net434),
    .D(net268),
    .Q(\i_main_reg.data_d[117] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1261_ (.RESET_B(net434),
    .D(net685),
    .Q(\i_main_reg.data_d[118] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1262_ (.RESET_B(net434),
    .D(net193),
    .Q(\i_main_reg.data_d[119] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _1263_ (.RESET_B(net434),
    .D(_0153_),
    .Q(\i_main_reg.data_d[120] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1264_ (.RESET_B(net434),
    .D(net169),
    .Q(\i_main_reg.data_d[121] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1265_ (.RESET_B(net436),
    .D(net531),
    .Q(\i_main_reg.data_d[122] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1266_ (.RESET_B(net436),
    .D(net608),
    .Q(\i_main_reg.data_d[123] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1267_ (.RESET_B(net436),
    .D(net664),
    .Q(\i_main_reg.data_d[124] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1268_ (.RESET_B(net436),
    .D(_0158_),
    .Q(\i_main_reg.data_d[125] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1269_ (.RESET_B(net436),
    .D(net655),
    .Q(\i_main_reg.data_d[126] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1270_ (.RESET_B(net436),
    .D(net658),
    .Q(\i_main_reg.data_d[127] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1271_ (.RESET_B(net436),
    .D(net277),
    .Q(\i_main_reg.data_d[128] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_1 _1272_ (.RESET_B(net436),
    .D(_0162_),
    .Q(\i_main_reg.data_d[129] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1273_ (.RESET_B(net432),
    .D(_0163_),
    .Q(\i_main_reg.data_d[130] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1274_ (.RESET_B(net432),
    .D(net292),
    .Q(\i_main_reg.data_d[131] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1275_ (.RESET_B(net432),
    .D(net612),
    .Q(\i_main_reg.data_d[132] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1276_ (.RESET_B(net432),
    .D(net290),
    .Q(\i_main_reg.data_d[133] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1277_ (.RESET_B(net432),
    .D(_0167_),
    .Q(\i_main_reg.data_d[134] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _1278_ (.RESET_B(net431),
    .D(_0168_),
    .Q(\i_main_reg.data_d[135] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1279_ (.RESET_B(net431),
    .D(net75),
    .Q(\i_main_reg.data_d[136] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1280_ (.RESET_B(net431),
    .D(net139),
    .Q(\i_main_reg.data_d[137] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1281_ (.RESET_B(net431),
    .D(_0171_),
    .Q(\i_main_reg.data_d[138] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1282_ (.RESET_B(net431),
    .D(net459),
    .Q(\i_main_reg.data_d[139] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1283_ (.RESET_B(net431),
    .D(net728),
    .Q(\i_main_reg.data_d[140] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1284_ (.RESET_B(net432),
    .D(net733),
    .Q(\i_main_reg.data_d[141] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1285_ (.RESET_B(net430),
    .D(net641),
    .Q(\i_main_reg.data_d[142] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1286_ (.RESET_B(net430),
    .D(_0176_),
    .Q(\i_main_reg.data_d[143] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1287_ (.RESET_B(net430),
    .D(_0177_),
    .Q(\i_main_reg.data_d[144] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1288_ (.RESET_B(net430),
    .D(net134),
    .Q(\i_main_reg.data_d[145] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1289_ (.RESET_B(net430),
    .D(net77),
    .Q(\i_main_reg.data_d[146] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1290_ (.RESET_B(net433),
    .D(_0180_),
    .Q(\i_main_reg.data_d[147] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1291_ (.RESET_B(net423),
    .D(net280),
    .Q(\i_main_reg.data_d[148] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _1292_ (.RESET_B(net423),
    .D(_0182_),
    .Q(\i_main_reg.data_d[149] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1293_ (.RESET_B(net423),
    .D(net497),
    .Q(\i_main_reg.data_d[150] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _1294_ (.RESET_B(net423),
    .D(net680),
    .Q(\i_main_reg.data_d[151] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1295_ (.RESET_B(net423),
    .D(net647),
    .Q(\i_main_reg.data_d[152] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1296_ (.RESET_B(net420),
    .D(_0186_),
    .Q(\i_main_reg.data_d[153] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1297_ (.RESET_B(net421),
    .D(_0187_),
    .Q(\i_main_reg.data_d[154] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1298_ (.RESET_B(net420),
    .D(_0188_),
    .Q(\i_main_reg.data_d[155] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1299_ (.RESET_B(net421),
    .D(net250),
    .Q(\i_main_reg.data_d[156] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1300_ (.RESET_B(net421),
    .D(_0190_),
    .Q(\i_main_reg.data_d[157] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1301_ (.RESET_B(net421),
    .D(net248),
    .Q(\i_main_reg.data_d[158] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1302_ (.RESET_B(net421),
    .D(net673),
    .Q(\i_main_reg.data_d[159] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _1303_ (.RESET_B(net422),
    .D(net197),
    .Q(\i_main_reg.data_d[160] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1304_ (.RESET_B(net422),
    .D(_0194_),
    .Q(\i_main_reg.data_d[161] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1305_ (.RESET_B(net422),
    .D(_0195_),
    .Q(\i_main_reg.data_d[162] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1306_ (.RESET_B(net422),
    .D(net71),
    .Q(\i_main_reg.data_d[163] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1307_ (.RESET_B(net423),
    .D(_0197_),
    .Q(\i_main_reg.data_d[164] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1308_ (.RESET_B(net423),
    .D(_0198_),
    .Q(\i_main_reg.data_d[165] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1309_ (.RESET_B(net422),
    .D(_0199_),
    .Q(\i_main_reg.data_d[166] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1310_ (.RESET_B(net429),
    .D(_0200_),
    .Q(\i_main_reg.data_d[167] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1311_ (.RESET_B(net429),
    .D(net172),
    .Q(\i_main_reg.data_d[168] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1312_ (.RESET_B(net429),
    .D(net542),
    .Q(\i_main_reg.data_d[169] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1313_ (.RESET_B(net429),
    .D(net465),
    .Q(\i_main_reg.data_d[170] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1314_ (.RESET_B(net429),
    .D(net270),
    .Q(\i_main_reg.data_d[171] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1315_ (.RESET_B(net431),
    .D(_0205_),
    .Q(\i_main_reg.data_d[172] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1316_ (.RESET_B(net431),
    .D(net132),
    .Q(\i_main_reg.data_d[173] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1317_ (.RESET_B(net429),
    .D(net638),
    .Q(\i_main_reg.data_d[174] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _1318_ (.RESET_B(net430),
    .D(_0208_),
    .Q(\i_main_reg.data_d[175] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1319_ (.RESET_B(net430),
    .D(_0209_),
    .Q(\i_main_reg.data_d[176] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _1320_ (.RESET_B(net429),
    .D(_0210_),
    .Q(\i_main_reg.data_d[177] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1321_ (.RESET_B(net429),
    .D(_0211_),
    .Q(\i_main_reg.data_d[178] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1322_ (.RESET_B(net422),
    .D(net199),
    .Q(\i_main_reg.data_d[179] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _1323_ (.RESET_B(net422),
    .D(net253),
    .Q(\i_main_reg.data_d[180] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1324_ (.RESET_B(net422),
    .D(_0214_),
    .Q(\i_main_reg.data_d[181] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1325_ (.RESET_B(net420),
    .D(net166),
    .Q(\i_main_reg.data_d[182] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _1326_ (.RESET_B(net420),
    .D(_0216_),
    .Q(\i_main_reg.data_d[183] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1327_ (.RESET_B(net420),
    .D(net120),
    .Q(\i_main_reg.data_d[184] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1328_ (.RESET_B(net420),
    .D(_0218_),
    .Q(\i_main_reg.data_d[185] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1329_ (.RESET_B(net420),
    .D(_0219_),
    .Q(\i_main_reg.data_d[186] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1330_ (.RESET_B(net420),
    .D(net59),
    .Q(\i_main_reg.data_d[187] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1331_ (.RESET_B(net392),
    .D(_0221_),
    .Q(\i_main_reg.data_d[188] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1332_ (.RESET_B(net392),
    .D(_0222_),
    .Q(\i_main_reg.data_d[189] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _1333_ (.RESET_B(net392),
    .D(net122),
    .Q(\i_main_reg.data_d[190] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1334_ (.RESET_B(net392),
    .D(net189),
    .Q(\i_main_reg.data_d[191] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _1335_ (.RESET_B(net392),
    .D(net46),
    .Q(\i_main_reg.data_d[192] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1336_ (.RESET_B(net392),
    .D(_0226_),
    .Q(\i_main_reg.data_d[193] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1337_ (.RESET_B(net392),
    .D(_0227_),
    .Q(\i_main_reg.data_d[194] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1338_ (.RESET_B(net392),
    .D(_0228_),
    .Q(\i_main_reg.data_d[195] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _1339_ (.RESET_B(net390),
    .D(_0229_),
    .Q(\i_main_reg.data_d[196] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1340_ (.RESET_B(net390),
    .D(_0230_),
    .Q(\i_main_reg.data_d[197] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1341_ (.RESET_B(net390),
    .D(_0231_),
    .Q(\i_main_reg.data_d[198] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1342_ (.RESET_B(net390),
    .D(net213),
    .Q(\i_main_reg.data_d[199] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1343_ (.RESET_B(net390),
    .D(net515),
    .Q(\i_main_reg.data_d[200] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1344_ (.RESET_B(net390),
    .D(_0234_),
    .Q(\i_main_reg.data_d[201] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1345_ (.RESET_B(net382),
    .D(_0235_),
    .Q(\i_main_reg.data_d[202] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1346_ (.RESET_B(net383),
    .D(net467),
    .Q(\i_main_reg.data_d[203] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1347_ (.RESET_B(net382),
    .D(net470),
    .Q(\i_main_reg.data_d[204] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1348_ (.RESET_B(net382),
    .D(net201),
    .Q(\i_main_reg.data_d[205] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1349_ (.RESET_B(net381),
    .D(_0239_),
    .Q(\i_main_reg.data_d[206] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1350_ (.RESET_B(net381),
    .D(_0240_),
    .Q(\i_main_reg.data_d[207] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1351_ (.RESET_B(net380),
    .D(_0241_),
    .Q(\i_main_reg.data_d[208] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1352_ (.RESET_B(net380),
    .D(net627),
    .Q(\i_main_reg.data_d[209] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1353_ (.RESET_B(net380),
    .D(net232),
    .Q(\i_main_reg.data_d[210] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1354_ (.RESET_B(net380),
    .D(_0244_),
    .Q(\i_main_reg.data_d[211] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net380),
    .D(net87),
    .Q(\i_main_reg.data_d[212] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _1356_ (.RESET_B(net380),
    .D(_0246_),
    .Q(\i_main_reg.data_d[213] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net380),
    .D(_0247_),
    .Q(\i_main_reg.data_d[214] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1358_ (.RESET_B(net380),
    .D(net479),
    .Q(\i_main_reg.data_d[215] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1359_ (.RESET_B(net381),
    .D(_0249_),
    .Q(\i_main_reg.data_d[216] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _1360_ (.RESET_B(net382),
    .D(net177),
    .Q(\i_main_reg.data_d[217] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1361_ (.RESET_B(net382),
    .D(net85),
    .Q(\i_main_reg.data_d[218] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net382),
    .D(_0252_),
    .Q(\i_main_reg.data_d[219] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net382),
    .D(_0253_),
    .Q(\i_main_reg.data_d[220] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1364_ (.RESET_B(net382),
    .D(_0254_),
    .Q(\i_main_reg.data_d[221] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1365_ (.RESET_B(net390),
    .D(net195),
    .Q(\i_main_reg.data_d[222] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _1366_ (.RESET_B(net391),
    .D(net245),
    .Q(\i_main_reg.data_d[223] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1367_ (.RESET_B(net390),
    .D(_0257_),
    .Q(\i_main_reg.data_d[224] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _1368_ (.RESET_B(net391),
    .D(net461),
    .Q(\i_main_reg.data_d[225] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1369_ (.RESET_B(net395),
    .D(net718),
    .Q(\i_main_reg.data_d[226] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1370_ (.RESET_B(net395),
    .D(_0260_),
    .Q(\i_main_reg.data_d[227] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1371_ (.RESET_B(net395),
    .D(_0261_),
    .Q(\i_main_reg.data_d[228] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _1372_ (.RESET_B(net396),
    .D(_0262_),
    .Q(\i_main_reg.data_d[229] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1373_ (.RESET_B(net396),
    .D(_0263_),
    .Q(\i_main_reg.data_d[230] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1374_ (.RESET_B(net396),
    .D(net146),
    .Q(\i_main_reg.data_d[231] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1375_ (.RESET_B(net396),
    .D(net554),
    .Q(\i_main_reg.data_d[232] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1376_ (.RESET_B(net396),
    .D(_0266_),
    .Q(\i_main_reg.data_d[233] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _1377_ (.RESET_B(net396),
    .D(_0267_),
    .Q(\i_main_reg.data_d[234] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net411),
    .D(net670),
    .Q(\i_main_reg.data_d[235] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1379_ (.RESET_B(net411),
    .D(net682),
    .Q(\i_main_reg.data_d[236] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net411),
    .D(net204),
    .Q(\i_main_reg.data_d[237] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1381_ (.RESET_B(net411),
    .D(_0271_),
    .Q(\i_main_reg.data_d[238] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1382_ (.RESET_B(net412),
    .D(net592),
    .Q(\i_main_reg.data_d[239] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1383_ (.RESET_B(net412),
    .D(_0273_),
    .Q(\i_main_reg.data_d[240] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1384_ (.RESET_B(net411),
    .D(net573),
    .Q(\i_main_reg.data_d[241] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net411),
    .D(net57),
    .Q(\i_main_reg.data_d[242] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1386_ (.RESET_B(net411),
    .D(_0276_),
    .Q(\i_main_reg.data_d[243] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net411),
    .D(_0277_),
    .Q(\i_main_reg.data_d[244] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1388_ (.RESET_B(net402),
    .D(_0278_),
    .Q(\i_main_reg.data_d[245] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net402),
    .D(net559),
    .Q(\i_main_reg.data_d[246] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1390_ (.RESET_B(net402),
    .D(net209),
    .Q(\i_main_reg.data_d[247] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net387),
    .D(_0281_),
    .Q(\i_main_reg.data_d[248] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1392_ (.RESET_B(net388),
    .D(_0282_),
    .Q(\i_main_reg.data_d[249] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1393_ (.RESET_B(net387),
    .D(_0283_),
    .Q(\i_main_reg.data_d[250] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1394_ (.RESET_B(net387),
    .D(_0284_),
    .Q(\i_main_reg.data_d[251] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net388),
    .D(net537),
    .Q(\i_main_reg.data_d[252] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net385),
    .D(net650),
    .Q(\i_main_reg.data_d[253] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1397_ (.RESET_B(net385),
    .D(net207),
    .Q(\i_main_reg.data_d[254] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net386),
    .D(_0288_),
    .Q(\i_main_reg.data_d[255] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1399_ (.RESET_B(net384),
    .D(_0289_),
    .Q(\i_main_reg.data_d[256] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1400_ (.RESET_B(net384),
    .D(_0290_),
    .Q(\i_main_reg.data_d[257] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1401_ (.RESET_B(net384),
    .D(_0291_),
    .Q(\i_main_reg.data_d[258] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net384),
    .D(net565),
    .Q(\i_main_reg.data_d[259] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1403_ (.RESET_B(net384),
    .D(_0293_),
    .Q(\i_main_reg.data_d[260] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net384),
    .D(_0294_),
    .Q(\i_main_reg.data_d[261] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1405_ (.RESET_B(net384),
    .D(net107),
    .Q(\i_main_reg.data_d[262] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net384),
    .D(net179),
    .Q(\i_main_reg.data_d[263] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1407_ (.RESET_B(net385),
    .D(_0297_),
    .Q(\i_main_reg.data_d[264] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1408_ (.RESET_B(net385),
    .D(_0298_),
    .Q(\i_main_reg.data_d[265] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1409_ (.RESET_B(net385),
    .D(net616),
    .Q(\i_main_reg.data_d[266] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1410_ (.RESET_B(net385),
    .D(net69),
    .Q(\i_main_reg.data_d[267] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1411_ (.RESET_B(net385),
    .D(_0301_),
    .Q(\i_main_reg.data_d[268] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_1 _1412_ (.RESET_B(net385),
    .D(net282),
    .Q(\i_main_reg.data_d[269] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net399),
    .D(_0303_),
    .Q(\i_main_reg.data_d[270] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net399),
    .D(net99),
    .Q(\i_main_reg.data_d[271] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net399),
    .D(_0305_),
    .Q(\i_main_reg.data_d[272] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1416_ (.RESET_B(net399),
    .D(net83),
    .Q(\i_main_reg.data_d[273] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net399),
    .D(net186),
    .Q(\i_main_reg.data_d[274] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1418_ (.RESET_B(net399),
    .D(net525),
    .Q(\i_main_reg.data_d[275] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1419_ (.RESET_B(net400),
    .D(net154),
    .Q(\i_main_reg.data_d[276] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net400),
    .D(_0310_),
    .Q(\i_main_reg.data_d[277] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net400),
    .D(net483),
    .Q(\i_main_reg.data_d[278] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net399),
    .D(_0312_),
    .Q(\i_main_reg.data_d[279] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net401),
    .D(_0313_),
    .Q(\i_main_reg.data_d[280] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net399),
    .D(net463),
    .Q(\i_main_reg.data_d[281] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1425_ (.RESET_B(net402),
    .D(_0315_),
    .Q(\i_main_reg.data_d[282] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net402),
    .D(net222),
    .Q(\i_main_reg.data_d[283] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net402),
    .D(_0317_),
    .Q(\i_main_reg.data_d[284] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net402),
    .D(_0318_),
    .Q(\i_main_reg.data_d[285] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net403),
    .D(_0319_),
    .Q(\i_main_reg.data_d[286] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net403),
    .D(net116),
    .Q(\i_main_reg.data_d[287] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1431_ (.RESET_B(net403),
    .D(net61),
    .Q(\i_main_reg.data_d[288] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net403),
    .D(_0322_),
    .Q(\i_main_reg.data_d[289] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net403),
    .D(_0323_),
    .Q(\i_main_reg.data_d[290] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net402),
    .D(_0324_),
    .Q(\i_main_reg.data_d[291] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net407),
    .D(_0325_),
    .Q(\i_main_reg.data_d[292] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1436_ (.RESET_B(net409),
    .D(_0326_),
    .Q(\i_main_reg.data_d[293] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1437_ (.RESET_B(net407),
    .D(net586),
    .Q(\i_main_reg.data_d[294] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1438_ (.RESET_B(net407),
    .D(_0328_),
    .Q(\i_main_reg.data_d[295] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1439_ (.RESET_B(net407),
    .D(net723),
    .Q(\i_main_reg.data_d[296] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1440_ (.RESET_B(net401),
    .D(_0330_),
    .Q(\i_main_reg.data_d[297] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1441_ (.RESET_B(net401),
    .D(_0331_),
    .Q(\i_main_reg.data_d[298] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1442_ (.RESET_B(net400),
    .D(net475),
    .Q(\i_main_reg.data_d[299] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1443_ (.RESET_B(net400),
    .D(net736),
    .Q(\i_main_reg.data_d[300] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net400),
    .D(net634),
    .Q(\i_main_reg.data_d[301] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net400),
    .D(_0335_),
    .Q(\i_main_reg.data_d[302] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net400),
    .D(net126),
    .Q(\i_main_reg.data_d[303] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net406),
    .D(_0337_),
    .Q(\i_main_reg.data_d[304] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1448_ (.RESET_B(net406),
    .D(_0338_),
    .Q(\i_main_reg.data_d[305] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net406),
    .D(_0339_),
    .Q(\i_main_reg.data_d[306] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net406),
    .D(_0340_),
    .Q(\i_main_reg.data_d[307] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net406),
    .D(net124),
    .Q(\i_main_reg.data_d[308] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net406),
    .D(_0342_),
    .Q(\i_main_reg.data_d[309] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net406),
    .D(_0343_),
    .Q(\i_main_reg.data_d[310] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net404),
    .D(net568),
    .Q(\i_main_reg.data_d[311] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net404),
    .D(net517),
    .Q(\i_main_reg.data_d[312] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1456_ (.RESET_B(net404),
    .D(_0346_),
    .Q(\i_main_reg.data_d[313] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net404),
    .D(_0347_),
    .Q(\i_main_reg.data_d[314] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net405),
    .D(net603),
    .Q(\i_main_reg.data_d[315] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net404),
    .D(_0349_),
    .Q(\i_main_reg.data_d[316] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net404),
    .D(net605),
    .Q(\i_main_reg.data_d[317] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net404),
    .D(net714),
    .Q(\i_main_reg.data_d[318] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1462_ (.RESET_B(net404),
    .D(net493),
    .Q(\i_main_reg.data_d[319] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1463_ (.RESET_B(net405),
    .D(_0353_),
    .Q(\i_main_reg.data_d[320] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1464_ (.RESET_B(net405),
    .D(_0354_),
    .Q(\i_main_reg.data_d[321] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1465_ (.RESET_B(net405),
    .D(net513),
    .Q(\i_main_reg.data_d[322] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1466_ (.RESET_B(net408),
    .D(_0356_),
    .Q(\i_main_reg.data_d[323] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1467_ (.RESET_B(net408),
    .D(net220),
    .Q(\i_main_reg.data_d[324] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1468_ (.RESET_B(net408),
    .D(net620),
    .Q(\i_main_reg.data_d[325] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net408),
    .D(net53),
    .Q(\i_main_reg.data_d[326] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net408),
    .D(_0360_),
    .Q(\i_main_reg.data_d[327] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net408),
    .D(_0361_),
    .Q(\i_main_reg.data_d[328] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1472_ (.RESET_B(net408),
    .D(net95),
    .Q(\i_main_reg.data_d[329] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _1473_ (.RESET_B(net407),
    .D(net226),
    .Q(\i_main_reg.data_d[330] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1474_ (.RESET_B(net407),
    .D(net55),
    .Q(\i_main_reg.data_d[331] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1475_ (.RESET_B(net407),
    .D(_0365_),
    .Q(\i_main_reg.data_d[332] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1476_ (.RESET_B(net407),
    .D(_0366_),
    .Q(\i_main_reg.data_d[333] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1477_ (.RESET_B(net408),
    .D(_0367_),
    .Q(\i_main_reg.data_d[334] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _1478_ (.RESET_B(net409),
    .D(_0368_),
    .Q(\i_main_reg.data_d[335] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1479_ (.RESET_B(net415),
    .D(net217),
    .Q(\i_main_reg.data_d[336] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net415),
    .D(net65),
    .Q(\i_main_reg.data_d[337] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net415),
    .D(_0371_),
    .Q(\i_main_reg.data_d[338] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net415),
    .D(net148),
    .Q(\i_main_reg.data_d[339] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1483_ (.RESET_B(net415),
    .D(_0373_),
    .Q(\i_main_reg.data_d[340] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net416),
    .D(_0374_),
    .Q(\i_main_reg.data_d[341] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1485_ (.RESET_B(net416),
    .D(net511),
    .Q(\i_main_reg.data_d[342] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1486_ (.RESET_B(net415),
    .D(_0376_),
    .Q(\i_main_reg.data_d[343] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1487_ (.RESET_B(net415),
    .D(_0377_),
    .Q(\i_main_reg.data_d[344] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1488_ (.RESET_B(net415),
    .D(net229),
    .Q(\i_main_reg.data_d[345] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1489_ (.RESET_B(net416),
    .D(_0379_),
    .Q(\i_main_reg.data_d[346] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net416),
    .D(_0380_),
    .Q(\i_main_reg.data_d[347] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1491_ (.RESET_B(net416),
    .D(net109),
    .Q(\i_main_reg.data_d[348] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net416),
    .D(_0382_),
    .Q(\i_main_reg.data_d[349] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _1493_ (.RESET_B(net412),
    .D(net260),
    .Q(\i_main_reg.data_d[350] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net412),
    .D(net73),
    .Q(\i_main_reg.data_d[351] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1495_ (.RESET_B(net413),
    .D(_0385_),
    .Q(\i_main_reg.data_d[352] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1496_ (.RESET_B(net413),
    .D(net141),
    .Q(\i_main_reg.data_d[353] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _1497_ (.RESET_B(net413),
    .D(_0387_),
    .Q(\i_main_reg.data_d[354] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net417),
    .D(net297),
    .Q(\i_main_reg.data_d[355] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1499_ (.RESET_B(net417),
    .D(net286),
    .Q(\i_main_reg.data_d[356] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1500_ (.RESET_B(net417),
    .D(_0390_),
    .Q(\i_main_reg.data_d[357] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1501_ (.RESET_B(net417),
    .D(net79),
    .Q(\i_main_reg.data_d[358] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net417),
    .D(net624),
    .Q(\i_main_reg.data_d[359] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1503_ (.RESET_B(net417),
    .D(net712),
    .Q(\i_main_reg.data_d[360] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _1504_ (.RESET_B(net418),
    .D(net702),
    .Q(\i_main_reg.data_d[361] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _1505_ (.RESET_B(net417),
    .D(net622),
    .Q(\i_main_reg.data_d[362] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net441),
    .D(net164),
    .Q(\i_main_reg.data_d[363] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _1507_ (.RESET_B(net441),
    .D(_0397_),
    .Q(\i_main_reg.data_d[364] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net442),
    .D(_0398_),
    .Q(\i_main_reg.data_d[365] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1509_ (.RESET_B(net442),
    .D(_0399_),
    .Q(\i_main_reg.data_d[366] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1510_ (.RESET_B(net442),
    .D(net257),
    .Q(\i_main_reg.data_d[367] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1511_ (.RESET_B(net442),
    .D(_0401_),
    .Q(\i_main_reg.data_d[368] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net442),
    .D(_0402_),
    .Q(\i_main_reg.data_d[369] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1513_ (.RESET_B(net441),
    .D(net191),
    .Q(\i_main_reg.data_d[370] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1514_ (.RESET_B(net444),
    .D(_0404_),
    .Q(\i_main_reg.data_d[371] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _1515_ (.RESET_B(net444),
    .D(_0405_),
    .Q(\i_main_reg.data_d[372] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1516_ (.RESET_B(net444),
    .D(_0406_),
    .Q(\i_main_reg.data_d[373] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _1517_ (.RESET_B(net443),
    .D(net294),
    .Q(\i_main_reg.data_d[374] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1518_ (.RESET_B(net443),
    .D(net539),
    .Q(\i_main_reg.data_d[375] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1519_ (.RESET_B(net443),
    .D(net488),
    .Q(\i_main_reg.data_d[376] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1520_ (.RESET_B(net443),
    .D(_0410_),
    .Q(\i_main_reg.data_d[377] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _1521_ (.RESET_B(net450),
    .D(net81),
    .Q(\i_main_reg.data_d[378] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1522_ (.RESET_B(net450),
    .D(net63),
    .Q(\i_main_reg.data_d[379] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1523_ (.RESET_B(net450),
    .D(_0413_),
    .Q(\i_main_reg.data_d[380] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1524_ (.RESET_B(net450),
    .D(net93),
    .Q(\i_main_reg.data_d[381] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _1525_ (.RESET_B(net448),
    .D(_0415_),
    .Q(\i_main_reg.data_d[382] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _1526_ (.RESET_B(net449),
    .D(net32),
    .Q(\one_count_q[0] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _1527_ (.RESET_B(net449),
    .D(net754),
    .Q(\one_count_q[1] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_6 (.L_LO(net6));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_7 (.L_LO(net7));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_8 (.L_LO(net8));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_9 (.L_LO(net9));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_10 (.L_LO(net10));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_11 (.L_LO(net11));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_12 (.L_LO(net12));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_13 (.L_LO(net13));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_14 (.L_LO(net14));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_15 (.L_LO(net15));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_16 (.L_LO(net16));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_17 (.L_LO(net17));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_18 (.L_LO(net18));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_19 (.L_LO(net19));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_20 (.L_LO(net20));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_21 (.L_LO(net21));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_22 (.L_LO(net22));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_23 (.L_LO(net23));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_24 (.L_LO(net24));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _1548_ (.A(\i_main_reg.data_o ),
    .X(uo_out[0]));
 sg13g2_buf_1 _1549_ (.A(\i_step_counter.data_o ),
    .X(uo_out[1]));
 sg13g2_buf_1 _1550_ (.A(finished_q),
    .X(uo_out[2]));
 sg13g2_buf_1 _1551_ (.A(overflow_q),
    .X(uo_out[3]));
 sg13g2_buf_8 fanout303 (.A(net304),
    .X(net303));
 sg13g2_buf_8 fanout304 (.A(net311),
    .X(net304));
 sg13g2_buf_8 fanout305 (.A(net311),
    .X(net305));
 sg13g2_buf_1 fanout306 (.A(net311),
    .X(net306));
 sg13g2_buf_8 fanout307 (.A(net310),
    .X(net307));
 sg13g2_buf_8 fanout308 (.A(net310),
    .X(net308));
 sg13g2_buf_8 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_8 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_8 fanout311 (.A(net340),
    .X(net311));
 sg13g2_buf_8 fanout312 (.A(net316),
    .X(net312));
 sg13g2_buf_8 fanout313 (.A(net316),
    .X(net313));
 sg13g2_buf_8 fanout314 (.A(net316),
    .X(net314));
 sg13g2_buf_2 fanout315 (.A(net316),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(net340),
    .X(net316));
 sg13g2_buf_8 fanout317 (.A(net320),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(net320),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_8 fanout320 (.A(net340),
    .X(net320));
 sg13g2_buf_8 fanout321 (.A(net323),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(net323),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(net332),
    .X(net323));
 sg13g2_buf_8 fanout324 (.A(net332),
    .X(net324));
 sg13g2_buf_1 fanout325 (.A(net332),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(net327),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_8 fanout328 (.A(net331),
    .X(net328));
 sg13g2_buf_8 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_8 fanout330 (.A(net331),
    .X(net330));
 sg13g2_buf_8 fanout331 (.A(net332),
    .X(net331));
 sg13g2_buf_2 fanout332 (.A(net340),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(net335),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(net335),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(net340),
    .X(net335));
 sg13g2_buf_8 fanout336 (.A(net339),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(net339),
    .X(net337));
 sg13g2_buf_8 fanout338 (.A(net339),
    .X(net338));
 sg13g2_buf_8 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_8 fanout340 (.A(_0552_),
    .X(net340));
 sg13g2_buf_8 fanout341 (.A(net344),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(net344),
    .X(net342));
 sg13g2_buf_8 fanout343 (.A(net344),
    .X(net343));
 sg13g2_buf_8 fanout344 (.A(net358),
    .X(net344));
 sg13g2_buf_8 fanout345 (.A(net348),
    .X(net345));
 sg13g2_buf_1 fanout346 (.A(net348),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(net358),
    .X(net348));
 sg13g2_buf_8 fanout349 (.A(net350),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net358),
    .X(net350));
 sg13g2_buf_8 fanout351 (.A(net353),
    .X(net351));
 sg13g2_buf_8 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_8 fanout353 (.A(net358),
    .X(net353));
 sg13g2_buf_8 fanout354 (.A(net357),
    .X(net354));
 sg13g2_buf_8 fanout355 (.A(net356),
    .X(net355));
 sg13g2_buf_8 fanout356 (.A(net357),
    .X(net356));
 sg13g2_buf_8 fanout357 (.A(net358),
    .X(net357));
 sg13g2_buf_8 fanout358 (.A(net370),
    .X(net358));
 sg13g2_buf_8 fanout359 (.A(net363),
    .X(net359));
 sg13g2_buf_1 fanout360 (.A(net363),
    .X(net360));
 sg13g2_buf_8 fanout361 (.A(net363),
    .X(net361));
 sg13g2_buf_1 fanout362 (.A(net363),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(net370),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net367),
    .X(net364));
 sg13g2_buf_8 fanout365 (.A(net367),
    .X(net365));
 sg13g2_buf_8 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_8 fanout367 (.A(net370),
    .X(net367));
 sg13g2_buf_8 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_8 fanout369 (.A(net370),
    .X(net369));
 sg13g2_buf_8 fanout370 (.A(_0552_),
    .X(net370));
 sg13g2_buf_8 fanout371 (.A(_0452_),
    .X(net371));
 sg13g2_buf_8 fanout372 (.A(_0449_),
    .X(net372));
 sg13g2_buf_2 fanout373 (.A(_0449_),
    .X(net373));
 sg13g2_buf_8 fanout374 (.A(net375),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(_0447_),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(_0441_),
    .X(net376));
 sg13g2_buf_1 fanout377 (.A(_0441_),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(\i_main_reg.data_o ),
    .X(net378));
 sg13g2_buf_1 fanout379 (.A(\i_main_reg.data_o ),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(net381),
    .X(net380));
 sg13g2_buf_8 fanout381 (.A(net389),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(net383),
    .X(net382));
 sg13g2_buf_8 fanout383 (.A(net389),
    .X(net383));
 sg13g2_buf_8 fanout384 (.A(net386),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(net388),
    .X(net386));
 sg13g2_buf_8 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_8 fanout389 (.A(net419),
    .X(net389));
 sg13g2_buf_8 fanout390 (.A(net394),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(net394),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(net394),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(net394),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(net419),
    .X(net394));
 sg13g2_buf_8 fanout395 (.A(net398),
    .X(net395));
 sg13g2_buf_8 fanout396 (.A(net398),
    .X(net396));
 sg13g2_buf_8 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(net419),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(net401),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(net401),
    .X(net400));
 sg13g2_buf_8 fanout401 (.A(net410),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(net410),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(net410),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_8 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_8 fanout406 (.A(net410),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(net409),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(net409),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(net410),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net418),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(net412),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(net414),
    .X(net412));
 sg13g2_buf_8 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_8 fanout414 (.A(net418),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(net416),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(net418),
    .X(net417));
 sg13g2_buf_8 fanout418 (.A(net419),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(rst_n),
    .X(net419));
 sg13g2_buf_8 fanout420 (.A(net428),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net428),
    .X(net421));
 sg13g2_buf_8 fanout422 (.A(net423),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(net428),
    .X(net423));
 sg13g2_buf_8 fanout424 (.A(net427),
    .X(net424));
 sg13g2_buf_8 fanout425 (.A(net427),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(net427),
    .X(net426));
 sg13g2_buf_8 fanout427 (.A(net428),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(net452),
    .X(net428));
 sg13g2_buf_8 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_8 fanout430 (.A(net433),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net433),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(net433),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(net452),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(net437),
    .X(net434));
 sg13g2_buf_1 fanout435 (.A(net437),
    .X(net435));
 sg13g2_buf_8 fanout436 (.A(net437),
    .X(net436));
 sg13g2_buf_8 fanout437 (.A(net452),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(net440),
    .X(net438));
 sg13g2_buf_8 fanout439 (.A(net440),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(net452),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(net444),
    .X(net441));
 sg13g2_buf_8 fanout442 (.A(net444),
    .X(net442));
 sg13g2_buf_8 fanout443 (.A(net444),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net452),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(net447),
    .X(net445));
 sg13g2_buf_8 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_8 fanout447 (.A(net451),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(net451),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(net450),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(net451),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(net452),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(rst_n),
    .X(net452));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_themightyduckofdoom_bitserial_collatz_checker_5 (.L_LO(net5));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_8 clkload3 (.A(clknet_leaf_52_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(overflow_q),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0517_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0017_),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold4 (.A(\bit_counter_q[4] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0540_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0024_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold7 (.A(\one_count_q[0] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0416_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold9 (.A(\bit_counter_q[9] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_step_counter.data_d[3] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0004_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold12 (.A(finished_q),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0512_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0016_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_main_reg.data_d[0] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0554_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_step_counter.data_d[6] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0006_),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold19 (.A(\bit_counter_q[5] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0543_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_main_reg.data_d[193] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0225_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold23 (.A(\bit_counter_q[1] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0533_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0021_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_main_reg.data_d[21] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0053_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_main_reg.data_d[327] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0359_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_main_reg.data_d[332] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0364_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_main_reg.data_d[243] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0275_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_main_reg.data_d[188] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0220_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_main_reg.data_d[289] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0321_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_main_reg.data_d[380] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0412_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_main_reg.data_d[338] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0370_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_main_reg.data_d[67] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0100_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_main_reg.data_d[268] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0300_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_main_reg.data_d[164] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0196_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_main_reg.data_d[352] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0384_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_main_reg.data_d[136] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0169_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_main_reg.data_d[147] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0179_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_main_reg.data_d[358] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0391_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_main_reg.data_d[378] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0411_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_main_reg.data_d[273] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0306_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_main_reg.data_d[219] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0251_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_main_reg.data_d[213] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0245_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_main_reg.data_d[244] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold65 (.A(\bit_counter_q[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0538_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0023_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_main_reg.data_d[382] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0414_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_main_reg.data_d[329] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0362_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_main_reg.data_d[63] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold73 (.A(_0096_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_main_reg.data_d[271] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0304_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_main_reg.data_d[104] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0137_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_main_reg.data_d[47] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0080_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_main_reg.data_d[25] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0057_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_main_reg.data_d[262] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0295_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_main_reg.data_d[348] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0381_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_main_reg.data_d[70] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0103_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_main_reg.data_d[220] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_main_reg.data_d[27] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0060_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_main_reg.data_d[287] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0320_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_main_reg.data_d[106] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0138_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_main_reg.data_d[185] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0217_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_main_reg.data_d[190] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold98 (.A(_0223_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_main_reg.data_d[309] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0341_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_main_reg.data_d[304] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0336_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_main_reg.data_d[57] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0090_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_main_reg.data_d[111] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0143_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_main_reg.data_d[173] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold108 (.A(_0206_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_main_reg.data_d[146] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0178_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_main_reg.data_d[65] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0098_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_main_reg.data_d[381] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_main_reg.data_d[138] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0170_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_main_reg.data_d[354] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0386_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_main_reg.data_d[286] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_main_reg.data_d[245] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_main_reg.data_d[103] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_main_reg.data_d[231] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0264_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_main_reg.data_d[340] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0372_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_main_reg.data_d[109] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0142_),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_main_reg.data_d[30] ),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0062_),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold129 (.A(\i_main_reg.data_d[277] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold130 (.A(_0309_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_main_reg.data_d[61] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0094_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_main_reg.data_d[64] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_main_reg.data_d[88] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0121_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold136 (.A(\i_main_reg.data_d[189] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_main_reg.data_d[194] ),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_main_reg.data_d[186] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_main_reg.data_d[364] ),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold140 (.A(_0396_),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_main_reg.data_d[183] ),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0215_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_main_reg.data_d[341] ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_main_reg.data_d[121] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0154_),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_main_reg.data_d[290] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_main_reg.data_d[168] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0201_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_main_reg.data_d[59] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0091_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_main_reg.data_d[31] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_main_reg.data_d[217] ),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0250_),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_main_reg.data_d[264] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0296_),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_main_reg.data_d[339] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_main_reg.data_d[328] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_step_counter.data_d[14] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0509_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0015_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_main_reg.data_d[274] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0307_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_main_reg.data_d[333] ),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold164 (.A(\i_main_reg.data_d[191] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0224_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_main_reg.data_d[370] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0403_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_main_reg.data_d[120] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0152_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_main_reg.data_d[222] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0255_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_main_reg.data_d[161] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0193_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_main_reg.data_d[179] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0212_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_main_reg.data_d[206] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0238_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_main_reg.data_d[305] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_main_reg.data_d[238] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0270_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_main_reg.data_d[167] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_main_reg.data_d[255] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0287_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_main_reg.data_d[248] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0280_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_main_reg.data_d[108] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0140_),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_main_reg.data_d[199] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0232_),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_main_reg.data_d[75] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0108_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_main_reg.data_d[336] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0369_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_main_reg.data_d[60] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_main_reg.data_d[324] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold196 (.A(_0357_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_main_reg.data_d[283] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0316_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_main_reg.data_d[81] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0113_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_main_reg.data_d[330] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0363_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_main_reg.data_d[62] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_main_reg.data_d[345] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0378_),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_main_reg.data_d[26] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_main_reg.data_d[211] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0243_),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_main_reg.data_d[85] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0118_),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_main_reg.data_d[113] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0146_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_main_reg.data_d[22] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold214 (.A(_0055_),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_main_reg.data_d[261] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_main_reg.data_d[272] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_main_reg.data_d[1] ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0034_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_main_reg.data_d[107] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_main_reg.data_d[224] ),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0256_),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_main_reg.data_d[285] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_main_reg.data_d[158] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0191_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_main_reg.data_d[156] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0189_),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_main_reg.data_d[214] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_main_reg.data_d[181] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0213_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_main_reg.data_d[41] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0074_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_main_reg.data_d[367] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0400_),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_main_reg.data_d[207] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_main_reg.data_d[350] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0383_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_main_reg.data_d[249] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_main_reg.data_d[366] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_main_reg.data_d[221] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold240 (.A(carry_q),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0525_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold242 (.A(_0018_),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_main_reg.data_d[117] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0150_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_main_reg.data_d[172] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0204_),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_main_reg.data_d[195] ),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_main_reg.data_d[29] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0061_),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_main_reg.data_d[182] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_main_reg.data_d[365] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_main_reg.data_d[129] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0161_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_main_reg.data_d[198] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_main_reg.data_d[148] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold256 (.A(_0181_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_main_reg.data_d[270] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0302_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_main_reg.data_d[18] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold260 (.A(_0051_),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_main_reg.data_d[357] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold262 (.A(_0389_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_main_reg.data_d[349] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_main_reg.data_d[178] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_main_reg.data_d[134] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0166_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_main_reg.data_d[131] ),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0164_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_main_reg.data_d[374] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0407_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_main_reg.data_d[306] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_main_reg.data_d[355] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0388_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_main_reg.data_d[256] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_main_reg.data_d[284] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_main_reg.data_d[2] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0035_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_main_reg.data_d[44] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold279 (.A(_0077_),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_main_reg.data_d[34] ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0067_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_main_reg.data_d[369] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold283 (.A(\i_main_reg.data_d[116] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_main_reg.data_d[139] ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0172_),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_main_reg.data_d[225] ),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0258_),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_main_reg.data_d[282] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0314_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_main_reg.data_d[171] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0203_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_main_reg.data_d[203] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold293 (.A(_0236_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_main_reg.data_d[162] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold295 (.A(\i_main_reg.data_d[204] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0237_),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_main_reg.data_d[82] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0115_),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_main_reg.data_d[269] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_main_reg.data_d[299] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold301 (.A(_0332_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold302 (.A(\i_main_reg.data_d[10] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0042_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_main_reg.data_d[216] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0248_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold306 (.A(\i_main_reg.data_d[368] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_main_reg.data_d[66] ),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold308 (.A(\i_main_reg.data_d[279] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0311_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold310 (.A(\i_main_reg.data_d[166] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_main_reg.data_d[54] ),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0087_),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_main_reg.data_d[377] ),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0409_),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_main_reg.data_d[46] ),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_main_reg.data_d[42] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold317 (.A(_0075_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold318 (.A(\i_main_reg.data_d[320] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold319 (.A(_0352_),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold320 (.A(\i_main_reg.data_d[14] ),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0047_),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold322 (.A(\i_main_reg.data_d[150] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0183_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold324 (.A(\i_main_reg.data_d[177] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold325 (.A(\i_main_reg.data_d[53] ),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold326 (.A(\i_main_reg.data_d[87] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold327 (.A(\i_main_reg.data_d[101] ),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold328 (.A(_0133_),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold329 (.A(\i_main_reg.data_d[196] ),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold330 (.A(\i_main_reg.data_d[23] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold331 (.A(_0056_),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold332 (.A(\i_main_reg.data_d[130] ),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold333 (.A(\i_main_reg.data_d[74] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold334 (.A(\i_main_reg.data_d[135] ),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold335 (.A(\i_main_reg.data_d[11] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold336 (.A(\i_main_reg.data_d[342] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0375_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold338 (.A(\i_main_reg.data_d[322] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0355_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold340 (.A(\i_main_reg.data_d[200] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0233_),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold342 (.A(\i_main_reg.data_d[313] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold343 (.A(_0345_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold344 (.A(\i_main_reg.data_d[55] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold345 (.A(_0088_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold346 (.A(\i_main_reg.data_d[373] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold347 (.A(\i_main_reg.data_d[157] ),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold348 (.A(\i_main_reg.data_d[73] ),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0105_),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold350 (.A(\i_main_reg.data_d[275] ),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0308_),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold352 (.A(\i_main_reg.data_d[187] ),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold353 (.A(\i_main_reg.data_d[49] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold354 (.A(_0082_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold355 (.A(\i_main_reg.data_d[202] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold356 (.A(\i_main_reg.data_d[122] ),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0155_),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold358 (.A(\i_main_reg.data_d[165] ),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold359 (.A(\i_main_reg.data_d[310] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold360 (.A(\i_main_reg.data_d[12] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold361 (.A(\i_main_reg.data_d[112] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold362 (.A(\i_main_reg.data_d[252] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold363 (.A(_0285_),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold364 (.A(\i_main_reg.data_d[375] ),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0408_),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold366 (.A(\i_main_reg.data_d[56] ),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold367 (.A(\i_main_reg.data_d[169] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold368 (.A(_0202_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold369 (.A(\i_main_reg.data_d[77] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0110_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold371 (.A(\i_main_reg.data_d[100] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0132_),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold373 (.A(\i_main_reg.data_d[149] ),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold374 (.A(\i_main_reg.data_d[215] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold375 (.A(\i_main_reg.data_d[278] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold376 (.A(\i_main_reg.data_d[334] ),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold377 (.A(\i_main_reg.data_d[230] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold378 (.A(\i_main_reg.data_d[208] ),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold379 (.A(\i_main_reg.data_d[233] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0265_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold381 (.A(\i_main_reg.data_d[43] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold382 (.A(\i_main_reg.data_d[314] ),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold383 (.A(\i_main_reg.data_d[69] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold384 (.A(\i_main_reg.data_d[246] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0279_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold386 (.A(\i_main_reg.data_d[176] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold387 (.A(\i_main_reg.data_d[76] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold388 (.A(\i_main_reg.data_d[50] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0083_),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold390 (.A(\i_main_reg.data_d[259] ),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0292_),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold392 (.A(\i_main_reg.data_d[68] ),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold393 (.A(\i_main_reg.data_d[312] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0344_),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold395 (.A(\i_main_reg.data_d[115] ),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold396 (.A(\i_main_reg.data_d[197] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold397 (.A(\i_main_reg.data_d[353] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold398 (.A(\i_main_reg.data_d[241] ),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0274_),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold400 (.A(\i_main_reg.data_d[311] ),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold401 (.A(\i_main_reg.data_d[335] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold402 (.A(\i_main_reg.data_d[184] ),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold403 (.A(\i_main_reg.data_d[37] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0070_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold405 (.A(\i_main_reg.data_d[291] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold406 (.A(\i_main_reg.data_d[323] ),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold407 (.A(\i_main_reg.data_d[265] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold408 (.A(\i_main_reg.data_d[16] ),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0048_),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold410 (.A(\i_main_reg.data_d[45] ),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold411 (.A(\i_main_reg.data_d[295] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0327_),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_main_reg.data_d[19] ),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0052_),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold415 (.A(\i_main_reg.data_d[280] ),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold416 (.A(\i_main_reg.data_d[102] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold417 (.A(\i_main_reg.data_d[239] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0272_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold419 (.A(\i_main_reg.data_d[114] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold420 (.A(\i_main_reg.data_d[163] ),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold421 (.A(\i_main_reg.data_d[344] ),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_main_reg.data_d[13] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold423 (.A(\i_main_reg.data_d[347] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold424 (.A(\i_main_reg.data_d[95] ),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0128_),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold426 (.A(\i_main_reg.data_d[99] ),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0131_),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold428 (.A(\i_main_reg.data_d[316] ),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold429 (.A(_0348_),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold430 (.A(\i_main_reg.data_d[317] ),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold431 (.A(_0350_),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold432 (.A(\i_main_reg.data_d[36] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold433 (.A(\i_main_reg.data_d[123] ),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold434 (.A(_0156_),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold435 (.A(\i_main_reg.data_d[40] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold436 (.A(\i_main_reg.data_d[258] ),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold437 (.A(\i_main_reg.data_d[133] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0165_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_main_reg.data_d[17] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold440 (.A(\i_main_reg.data_d[94] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold441 (.A(\i_main_reg.data_d[267] ),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0299_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold443 (.A(\i_main_reg.data_d[84] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0116_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold445 (.A(\i_main_reg.data_d[325] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0358_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_main_reg.data_d[363] ),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0395_),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold449 (.A(\i_main_reg.data_d[359] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0392_),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold451 (.A(\i_main_reg.data_d[307] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold452 (.A(\i_main_reg.data_d[209] ),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold453 (.A(_0242_),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold454 (.A(\i_main_reg.data_d[372] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold455 (.A(\i_main_reg.data_d[89] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0122_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold457 (.A(\i_main_reg.data_d[32] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0065_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold459 (.A(\i_main_reg.data_d[302] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0334_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold461 (.A(\i_main_reg.data_d[212] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold462 (.A(\i_main_reg.data_d[229] ),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold463 (.A(\i_main_reg.data_d[174] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0207_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold465 (.A(\i_main_reg.data_d[292] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold466 (.A(\i_main_reg.data_d[143] ),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold467 (.A(_0175_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold468 (.A(\i_main_reg.data_d[260] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold469 (.A(\i_main_reg.data_d[52] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold470 (.A(\i_main_reg.data_d[293] ),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold471 (.A(\i_main_reg.data_d[93] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold472 (.A(\i_main_reg.data_d[153] ),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold473 (.A(_0185_),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold474 (.A(\i_main_reg.data_d[240] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold475 (.A(\i_main_reg.data_d[254] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0286_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold477 (.A(\i_main_reg.data_d[321] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold478 (.A(\i_main_reg.data_d[251] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold479 (.A(\i_main_reg.data_d[201] ),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold480 (.A(\i_main_reg.data_d[126] ),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold481 (.A(_0159_),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold482 (.A(\i_main_reg.data_d[308] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold483 (.A(\i_main_reg.data_d[128] ),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0160_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold485 (.A(\i_main_reg.data_d[155] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold486 (.A(\i_main_reg.data_d[343] ),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold487 (.A(\i_main_reg.data_d[315] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold488 (.A(\i_main_reg.data_d[281] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold489 (.A(\i_main_reg.data_d[125] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0157_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold491 (.A(\i_main_reg.data_d[72] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold492 (.A(_0104_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold493 (.A(\i_main_reg.data_d[80] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0112_),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold495 (.A(\i_main_reg.data_d[235] ),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0268_),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold497 (.A(\i_main_reg.data_d[266] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold498 (.A(\i_main_reg.data_d[159] ),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0192_),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold500 (.A(\i_main_reg.data_d[48] ),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold501 (.A(\i_main_reg.data_d[4] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0037_),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold503 (.A(\i_main_reg.data_d[234] ),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold504 (.A(\i_main_reg.data_d[175] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold505 (.A(\i_main_reg.data_d[151] ),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0184_),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold507 (.A(\i_main_reg.data_d[237] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0269_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold509 (.A(\i_main_reg.data_d[3] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold510 (.A(\i_main_reg.data_d[119] ),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0151_),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold512 (.A(\i_main_reg.data_d[154] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold513 (.A(\i_main_reg.data_d[303] ),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold514 (.A(\i_main_reg.data_d[250] ),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold515 (.A(\i_main_reg.data_d[298] ),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold516 (.A(\i_main_reg.data_d[79] ),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold517 (.A(_0111_),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold518 (.A(\i_main_reg.data_d[33] ),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold519 (.A(\i_main_reg.data_d[35] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold520 (.A(\i_main_reg.data_d[38] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold521 (.A(_0071_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold522 (.A(\i_main_reg.data_d[228] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold523 (.A(\i_main_reg.data_d[6] ),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold524 (.A(_0039_),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold525 (.A(\i_main_reg.data_d[8] ),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold526 (.A(_0040_),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold527 (.A(\i_main_reg.data_d[362] ),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold528 (.A(_0394_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold529 (.A(\i_main_reg.data_d[346] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold530 (.A(\i_main_reg.data_d[92] ),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0124_),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold532 (.A(\i_main_reg.data_d[51] ),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold533 (.A(\i_main_reg.data_d[96] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold534 (.A(_0129_),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold535 (.A(\i_step_counter.data_o ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold536 (.A(_0000_),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold537 (.A(\i_main_reg.data_d[360] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold538 (.A(_0393_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold539 (.A(\i_main_reg.data_d[318] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0351_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold541 (.A(\bit_counter_q[8] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0028_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold543 (.A(\i_main_reg.data_d[227] ),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0259_),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold545 (.A(\i_step_counter.data_d[11] ),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0501_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0013_),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold548 (.A(\i_main_reg.data_d[296] ),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold549 (.A(_0329_),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold550 (.A(\i_main_reg.data_d[86] ),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold551 (.A(\i_step_counter.data_d[2] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold552 (.A(_0002_),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold553 (.A(\i_main_reg.data_d[140] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold554 (.A(_0173_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold555 (.A(\i_main_reg.data_d[5] ),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold556 (.A(\i_main_reg.data_d[98] ),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold557 (.A(_0130_),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold558 (.A(\i_main_reg.data_d[141] ),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0174_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold560 (.A(\i_main_reg.data_d[9] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold561 (.A(\i_main_reg.data_d[300] ),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold562 (.A(_0333_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold563 (.A(\i_main_reg.data_d[257] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold564 (.A(\i_main_reg.data_d[297] ),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold565 (.A(\i_main_reg.data_d[39] ),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_step_counter.data_d[9] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold567 (.A(_0492_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold568 (.A(_0011_),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold569 (.A(\i_main_reg.data_d[91] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold570 (.A(_0123_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold571 (.A(\bit_counter_q[7] ),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold572 (.A(_0547_),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold573 (.A(_0027_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold574 (.A(\i_main_reg.data_d[144] ),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold575 (.A(\bit_counter_q[6] ),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold576 (.A(_0545_),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold577 (.A(\i_main_reg.data_d[371] ),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold578 (.A(\i_main_reg.data_d[145] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold579 (.A(\one_count_q[1] ),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold580 (.A(_0417_),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold581 (.A(\i_step_counter.data_d[13] ),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold582 (.A(_0014_),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold583 (.A(\i_main_reg.data_d[294] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold584 (.A(previous_bit_q),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold585 (.A(_0526_),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold586 (.A(\bit_counter_q[0] ),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold587 (.A(\state_q[0] ),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold588 (.A(_0421_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold589 (.A(\bit_counter_q[2] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold590 (.A(\i_step_counter.data_d[1] ),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold591 (.A(_0001_),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold592 (.A(\i_step_counter.data_d[8] ),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold593 (.A(_0491_),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold594 (.A(_0010_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_step_counter.data_d[0] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold596 (.A(\i_step_counter.data_d[7] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_step_counter.data_d[4] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold598 (.A(_0472_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold599 (.A(\i_step_counter.data_d[5] ),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold600 (.A(\state_q[1] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold601 (.A(\i_step_counter.data_d[12] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold602 (.A(_0012_),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold603 (.A(\state_q[0] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold604 (.A(\state_q[1] ),
    .X(net778));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_126 ();
 sg13g2_decap_4 FILLER_0_209 ();
 sg13g2_fill_2 FILLER_0_250 ();
 sg13g2_fill_1 FILLER_0_252 ();
 sg13g2_fill_1 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_fill_1 FILLER_1_119 ();
 sg13g2_decap_4 FILLER_1_192 ();
 sg13g2_decap_4 FILLER_1_214 ();
 sg13g2_fill_2 FILLER_1_218 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_fill_2 FILLER_2_112 ();
 sg13g2_fill_1 FILLER_2_114 ();
 sg13g2_decap_8 FILLER_2_143 ();
 sg13g2_fill_2 FILLER_2_159 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_fill_2 FILLER_2_189 ();
 sg13g2_fill_1 FILLER_2_191 ();
 sg13g2_fill_2 FILLER_2_201 ();
 sg13g2_fill_1 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_222 ();
 sg13g2_decap_4 FILLER_2_250 ();
 sg13g2_fill_2 FILLER_2_254 ();
 sg13g2_decap_4 FILLER_2_346 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_4 FILLER_3_98 ();
 sg13g2_fill_2 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_3_176 ();
 sg13g2_decap_4 FILLER_3_193 ();
 sg13g2_decap_4 FILLER_3_206 ();
 sg13g2_decap_4 FILLER_3_247 ();
 sg13g2_fill_1 FILLER_3_261 ();
 sg13g2_fill_1 FILLER_3_272 ();
 sg13g2_fill_2 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_fill_1 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_fill_2 FILLER_4_207 ();
 sg13g2_decap_4 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_242 ();
 sg13g2_decap_4 FILLER_4_317 ();
 sg13g2_fill_2 FILLER_4_321 ();
 sg13g2_fill_2 FILLER_4_360 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_fill_1 FILLER_5_145 ();
 sg13g2_decap_4 FILLER_5_237 ();
 sg13g2_fill_2 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_253 ();
 sg13g2_decap_4 FILLER_5_277 ();
 sg13g2_fill_1 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_fill_1 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_96 ();
 sg13g2_decap_4 FILLER_6_171 ();
 sg13g2_fill_2 FILLER_6_212 ();
 sg13g2_decap_4 FILLER_6_321 ();
 sg13g2_fill_2 FILLER_6_362 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_fill_2 FILLER_7_96 ();
 sg13g2_fill_1 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_109 ();
 sg13g2_decap_4 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_164 ();
 sg13g2_fill_1 FILLER_7_166 ();
 sg13g2_fill_1 FILLER_7_200 ();
 sg13g2_fill_1 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_fill_1 FILLER_7_362 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_4 FILLER_8_63 ();
 sg13g2_fill_1 FILLER_8_95 ();
 sg13g2_fill_2 FILLER_8_159 ();
 sg13g2_fill_1 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_236 ();
 sg13g2_fill_2 FILLER_8_240 ();
 sg13g2_decap_4 FILLER_8_282 ();
 sg13g2_fill_2 FILLER_8_326 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_4 FILLER_9_56 ();
 sg13g2_fill_2 FILLER_9_60 ();
 sg13g2_decap_4 FILLER_9_125 ();
 sg13g2_fill_2 FILLER_9_129 ();
 sg13g2_decap_8 FILLER_9_184 ();
 sg13g2_decap_4 FILLER_9_218 ();
 sg13g2_fill_2 FILLER_9_222 ();
 sg13g2_fill_1 FILLER_9_251 ();
 sg13g2_fill_1 FILLER_9_279 ();
 sg13g2_fill_1 FILLER_9_290 ();
 sg13g2_fill_1 FILLER_9_340 ();
 sg13g2_fill_1 FILLER_9_368 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_fill_2 FILLER_10_49 ();
 sg13g2_fill_1 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_140 ();
 sg13g2_decap_4 FILLER_10_205 ();
 sg13g2_fill_1 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_decap_4 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_4 FILLER_10_365 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_4 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_60 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_fill_1 FILLER_11_133 ();
 sg13g2_decap_4 FILLER_11_160 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_decap_4 FILLER_11_205 ();
 sg13g2_fill_1 FILLER_11_209 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_decap_4 FILLER_11_270 ();
 sg13g2_fill_2 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_303 ();
 sg13g2_fill_1 FILLER_11_305 ();
 sg13g2_decap_4 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_96 ();
 sg13g2_decap_4 FILLER_12_144 ();
 sg13g2_fill_1 FILLER_12_148 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_213 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_decap_8 FILLER_12_271 ();
 sg13g2_decap_4 FILLER_12_305 ();
 sg13g2_fill_1 FILLER_12_309 ();
 sg13g2_decap_8 FILLER_12_401 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_4 FILLER_13_49 ();
 sg13g2_fill_2 FILLER_13_127 ();
 sg13g2_fill_1 FILLER_13_156 ();
 sg13g2_decap_4 FILLER_13_170 ();
 sg13g2_decap_8 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_decap_4 FILLER_13_229 ();
 sg13g2_fill_1 FILLER_13_243 ();
 sg13g2_decap_8 FILLER_13_290 ();
 sg13g2_decap_4 FILLER_13_310 ();
 sg13g2_fill_2 FILLER_13_314 ();
 sg13g2_decap_4 FILLER_13_356 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_4 FILLER_14_49 ();
 sg13g2_fill_2 FILLER_14_98 ();
 sg13g2_fill_1 FILLER_14_100 ();
 sg13g2_fill_1 FILLER_14_141 ();
 sg13g2_fill_2 FILLER_14_329 ();
 sg13g2_fill_1 FILLER_14_331 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_121 ();
 sg13g2_fill_1 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_205 ();
 sg13g2_decap_4 FILLER_15_216 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_decap_4 FILLER_15_248 ();
 sg13g2_fill_1 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_4 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_60 ();
 sg13g2_decap_4 FILLER_16_269 ();
 sg13g2_fill_1 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_4 FILLER_17_56 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_fill_2 FILLER_17_102 ();
 sg13g2_decap_4 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_234 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_fill_1 FILLER_17_304 ();
 sg13g2_decap_4 FILLER_17_342 ();
 sg13g2_fill_2 FILLER_17_346 ();
 sg13g2_decap_8 FILLER_17_402 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_fill_2 FILLER_18_42 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_159 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_185 ();
 sg13g2_fill_1 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_fill_1 FILLER_18_224 ();
 sg13g2_fill_1 FILLER_18_235 ();
 sg13g2_fill_1 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_316 ();
 sg13g2_fill_1 FILLER_18_318 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_decap_4 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_239 ();
 sg13g2_fill_1 FILLER_19_241 ();
 sg13g2_decap_4 FILLER_19_283 ();
 sg13g2_fill_2 FILLER_19_314 ();
 sg13g2_fill_1 FILLER_19_316 ();
 sg13g2_fill_2 FILLER_19_344 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_4 FILLER_20_35 ();
 sg13g2_decap_4 FILLER_20_95 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_2 FILLER_20_196 ();
 sg13g2_fill_2 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_fill_1 FILLER_20_299 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_1 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_99 ();
 sg13g2_decap_4 FILLER_21_127 ();
 sg13g2_fill_2 FILLER_21_131 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_fill_1 FILLER_21_207 ();
 sg13g2_fill_2 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_4 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_decap_4 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_228 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_fill_2 FILLER_23_42 ();
 sg13g2_fill_1 FILLER_23_44 ();
 sg13g2_fill_2 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_101 ();
 sg13g2_fill_2 FILLER_23_195 ();
 sg13g2_fill_1 FILLER_23_197 ();
 sg13g2_fill_1 FILLER_23_266 ();
 sg13g2_fill_2 FILLER_23_307 ();
 sg13g2_fill_1 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_4 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_fill_2 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_44 ();
 sg13g2_decap_4 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_2 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_303 ();
 sg13g2_fill_1 FILLER_25_310 ();
 sg13g2_decap_8 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_372 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_39 ();
 sg13g2_decap_8 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_148 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_200 ();
 sg13g2_fill_2 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_4 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_fill_1 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_227 ();
 sg13g2_fill_1 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_fill_1 FILLER_27_252 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_fill_2 FILLER_27_406 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_fill_1 FILLER_28_49 ();
 sg13g2_fill_2 FILLER_28_104 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_fill_1 FILLER_28_182 ();
 sg13g2_decap_4 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_267 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_decap_4 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_104 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_260 ();
 sg13g2_decap_8 FILLER_29_350 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_4 FILLER_30_35 ();
 sg13g2_fill_1 FILLER_30_39 ();
 sg13g2_fill_2 FILLER_30_177 ();
 sg13g2_decap_4 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_decap_8 FILLER_31_101 ();
 sg13g2_fill_1 FILLER_31_108 ();
 sg13g2_fill_1 FILLER_31_149 ();
 sg13g2_decap_4 FILLER_31_214 ();
 sg13g2_fill_1 FILLER_31_218 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_fill_2 FILLER_32_49 ();
 sg13g2_fill_2 FILLER_32_141 ();
 sg13g2_decap_8 FILLER_32_216 ();
 sg13g2_decap_8 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_297 ();
 sg13g2_decap_8 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_371 ();
 sg13g2_decap_8 FILLER_32_378 ();
 sg13g2_decap_8 FILLER_32_385 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_399 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_fill_2 FILLER_33_104 ();
 sg13g2_fill_1 FILLER_33_106 ();
 sg13g2_fill_2 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_217 ();
 sg13g2_decap_4 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_245 ();
 sg13g2_fill_2 FILLER_33_300 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_344 ();
 sg13g2_decap_8 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_33_358 ();
 sg13g2_decap_8 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_33_372 ();
 sg13g2_decap_8 FILLER_33_379 ();
 sg13g2_decap_8 FILLER_33_386 ();
 sg13g2_decap_8 FILLER_33_393 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_63 ();
 sg13g2_decap_4 FILLER_34_103 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_fill_1 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_decap_4 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_358 ();
 sg13g2_decap_8 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_fill_2 FILLER_35_56 ();
 sg13g2_fill_1 FILLER_35_58 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_208 ();
 sg13g2_decap_4 FILLER_35_276 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_361 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_fill_2 FILLER_36_153 ();
 sg13g2_decap_4 FILLER_36_232 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_decap_8 FILLER_37_138 ();
 sg13g2_fill_2 FILLER_37_172 ();
 sg13g2_decap_4 FILLER_37_211 ();
 sg13g2_fill_2 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_227 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_fill_2 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_decap_8 FILLER_37_351 ();
 sg13g2_decap_8 FILLER_37_358 ();
 sg13g2_decap_8 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_372 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_77 ();
 sg13g2_decap_4 FILLER_38_120 ();
 sg13g2_decap_8 FILLER_38_178 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_fill_1 FILLER_38_236 ();
 sg13g2_decap_4 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_351 ();
 sg13g2_decap_8 FILLER_38_358 ();
 sg13g2_decap_8 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_372 ();
 sg13g2_decap_8 FILLER_38_379 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_fill_1 FILLER_39_63 ();
 sg13g2_fill_1 FILLER_39_119 ();
 sg13g2_decap_4 FILLER_39_152 ();
 sg13g2_fill_1 FILLER_39_166 ();
 sg13g2_fill_2 FILLER_39_204 ();
 sg13g2_fill_1 FILLER_39_206 ();
 sg13g2_decap_8 FILLER_39_234 ();
 sg13g2_fill_1 FILLER_39_241 ();
 sg13g2_decap_8 FILLER_39_360 ();
 sg13g2_decap_8 FILLER_39_367 ();
 sg13g2_decap_8 FILLER_39_374 ();
 sg13g2_decap_8 FILLER_39_381 ();
 sg13g2_decap_8 FILLER_39_388 ();
 sg13g2_decap_8 FILLER_39_395 ();
 sg13g2_decap_8 FILLER_39_402 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_4 FILLER_40_56 ();
 sg13g2_fill_2 FILLER_40_60 ();
 sg13g2_decap_4 FILLER_40_117 ();
 sg13g2_fill_2 FILLER_40_121 ();
 sg13g2_fill_2 FILLER_40_143 ();
 sg13g2_decap_8 FILLER_40_165 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_decap_8 FILLER_40_351 ();
 sg13g2_decap_8 FILLER_40_358 ();
 sg13g2_decap_8 FILLER_40_365 ();
 sg13g2_decap_8 FILLER_40_372 ();
 sg13g2_decap_8 FILLER_40_379 ();
 sg13g2_decap_8 FILLER_40_386 ();
 sg13g2_decap_8 FILLER_40_393 ();
 sg13g2_decap_8 FILLER_40_400 ();
 sg13g2_fill_2 FILLER_40_407 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_4 FILLER_41_70 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_decap_8 FILLER_41_103 ();
 sg13g2_fill_2 FILLER_41_146 ();
 sg13g2_decap_4 FILLER_41_175 ();
 sg13g2_fill_2 FILLER_41_266 ();
 sg13g2_decap_4 FILLER_41_278 ();
 sg13g2_fill_1 FILLER_41_282 ();
 sg13g2_decap_8 FILLER_41_355 ();
 sg13g2_decap_8 FILLER_41_362 ();
 sg13g2_decap_8 FILLER_41_369 ();
 sg13g2_decap_8 FILLER_41_376 ();
 sg13g2_decap_8 FILLER_41_383 ();
 sg13g2_decap_8 FILLER_41_390 ();
 sg13g2_decap_8 FILLER_41_397 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_decap_8 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_70 ();
 sg13g2_decap_4 FILLER_42_116 ();
 sg13g2_fill_2 FILLER_42_120 ();
 sg13g2_decap_4 FILLER_42_251 ();
 sg13g2_fill_2 FILLER_42_255 ();
 sg13g2_decap_8 FILLER_42_294 ();
 sg13g2_fill_1 FILLER_42_301 ();
 sg13g2_decap_8 FILLER_42_342 ();
 sg13g2_decap_8 FILLER_42_349 ();
 sg13g2_decap_8 FILLER_42_356 ();
 sg13g2_decap_8 FILLER_42_363 ();
 sg13g2_decap_8 FILLER_42_370 ();
 sg13g2_decap_8 FILLER_42_377 ();
 sg13g2_decap_8 FILLER_42_384 ();
 sg13g2_decap_8 FILLER_42_391 ();
 sg13g2_decap_8 FILLER_42_398 ();
 sg13g2_decap_4 FILLER_42_405 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_244 ();
 sg13g2_fill_1 FILLER_43_251 ();
 sg13g2_fill_1 FILLER_43_265 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_fill_2 FILLER_43_406 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_decap_8 FILLER_44_49 ();
 sg13g2_decap_4 FILLER_44_56 ();
 sg13g2_fill_1 FILLER_44_60 ();
 sg13g2_decap_8 FILLER_44_116 ();
 sg13g2_fill_1 FILLER_44_123 ();
 sg13g2_fill_2 FILLER_44_179 ();
 sg13g2_decap_8 FILLER_44_258 ();
 sg13g2_fill_1 FILLER_44_265 ();
 sg13g2_fill_2 FILLER_44_293 ();
 sg13g2_decap_8 FILLER_44_350 ();
 sg13g2_decap_8 FILLER_44_357 ();
 sg13g2_decap_8 FILLER_44_364 ();
 sg13g2_decap_8 FILLER_44_371 ();
 sg13g2_decap_8 FILLER_44_378 ();
 sg13g2_decap_8 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_392 ();
 sg13g2_decap_8 FILLER_44_399 ();
 sg13g2_fill_2 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_408 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_4 FILLER_45_63 ();
 sg13g2_fill_2 FILLER_45_67 ();
 sg13g2_decap_4 FILLER_45_123 ();
 sg13g2_fill_1 FILLER_45_149 ();
 sg13g2_fill_1 FILLER_45_183 ();
 sg13g2_fill_2 FILLER_45_221 ();
 sg13g2_fill_2 FILLER_45_264 ();
 sg13g2_fill_1 FILLER_45_266 ();
 sg13g2_decap_4 FILLER_45_277 ();
 sg13g2_fill_2 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_396 ();
 sg13g2_decap_4 FILLER_45_403 ();
 sg13g2_fill_2 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_4 FILLER_46_70 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_fill_2 FILLER_46_157 ();
 sg13g2_fill_1 FILLER_46_159 ();
 sg13g2_decap_4 FILLER_46_187 ();
 sg13g2_decap_8 FILLER_46_272 ();
 sg13g2_fill_1 FILLER_46_279 ();
 sg13g2_fill_2 FILLER_46_320 ();
 sg13g2_decap_8 FILLER_46_367 ();
 sg13g2_decap_8 FILLER_46_374 ();
 sg13g2_decap_8 FILLER_46_381 ();
 sg13g2_decap_8 FILLER_46_388 ();
 sg13g2_decap_8 FILLER_46_395 ();
 sg13g2_decap_8 FILLER_46_402 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_4 FILLER_47_63 ();
 sg13g2_fill_2 FILLER_47_118 ();
 sg13g2_fill_1 FILLER_47_120 ();
 sg13g2_decap_8 FILLER_47_185 ();
 sg13g2_fill_1 FILLER_47_192 ();
 sg13g2_fill_2 FILLER_47_222 ();
 sg13g2_fill_1 FILLER_47_224 ();
 sg13g2_fill_2 FILLER_47_235 ();
 sg13g2_fill_2 FILLER_47_284 ();
 sg13g2_fill_1 FILLER_47_286 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_decap_8 FILLER_47_397 ();
 sg13g2_decap_4 FILLER_47_404 ();
 sg13g2_fill_1 FILLER_47_408 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_117 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_160 ();
 sg13g2_decap_4 FILLER_48_190 ();
 sg13g2_fill_1 FILLER_48_194 ();
 sg13g2_decap_4 FILLER_48_283 ();
 sg13g2_fill_1 FILLER_48_287 ();
 sg13g2_fill_1 FILLER_48_321 ();
 sg13g2_decap_8 FILLER_48_367 ();
 sg13g2_decap_8 FILLER_48_374 ();
 sg13g2_decap_8 FILLER_48_381 ();
 sg13g2_decap_8 FILLER_48_388 ();
 sg13g2_decap_8 FILLER_48_395 ();
 sg13g2_decap_8 FILLER_48_402 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_4 FILLER_49_56 ();
 sg13g2_fill_2 FILLER_49_60 ();
 sg13g2_fill_2 FILLER_49_116 ();
 sg13g2_fill_1 FILLER_49_118 ();
 sg13g2_fill_2 FILLER_49_156 ();
 sg13g2_decap_4 FILLER_49_185 ();
 sg13g2_fill_1 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_257 ();
 sg13g2_fill_2 FILLER_49_296 ();
 sg13g2_fill_1 FILLER_49_298 ();
 sg13g2_fill_2 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_fill_1 FILLER_50_56 ();
 sg13g2_decap_4 FILLER_50_140 ();
 sg13g2_fill_2 FILLER_50_167 ();
 sg13g2_fill_1 FILLER_50_216 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_fill_2 FILLER_50_258 ();
 sg13g2_decap_8 FILLER_50_377 ();
 sg13g2_decap_8 FILLER_50_384 ();
 sg13g2_decap_8 FILLER_50_391 ();
 sg13g2_decap_8 FILLER_50_398 ();
 sg13g2_decap_4 FILLER_50_405 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_8 FILLER_51_49 ();
 sg13g2_fill_2 FILLER_51_56 ();
 sg13g2_fill_1 FILLER_51_58 ();
 sg13g2_fill_1 FILLER_51_115 ();
 sg13g2_decap_8 FILLER_51_183 ();
 sg13g2_fill_2 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_219 ();
 sg13g2_decap_4 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_309 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_4 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_56 ();
 sg13g2_fill_2 FILLER_52_156 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_2 FILLER_52_219 ();
 sg13g2_fill_1 FILLER_52_221 ();
 sg13g2_decap_8 FILLER_52_235 ();
 sg13g2_fill_1 FILLER_52_242 ();
 sg13g2_decap_8 FILLER_52_395 ();
 sg13g2_decap_8 FILLER_52_402 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_4 FILLER_53_56 ();
 sg13g2_fill_1 FILLER_53_115 ();
 sg13g2_decap_4 FILLER_53_169 ();
 sg13g2_fill_1 FILLER_53_173 ();
 sg13g2_fill_2 FILLER_53_228 ();
 sg13g2_decap_8 FILLER_53_381 ();
 sg13g2_decap_8 FILLER_53_388 ();
 sg13g2_decap_8 FILLER_53_395 ();
 sg13g2_decap_8 FILLER_53_402 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_decap_4 FILLER_54_56 ();
 sg13g2_decap_8 FILLER_54_154 ();
 sg13g2_fill_1 FILLER_54_161 ();
 sg13g2_fill_1 FILLER_54_189 ();
 sg13g2_decap_4 FILLER_54_250 ();
 sg13g2_fill_1 FILLER_54_331 ();
 sg13g2_decap_8 FILLER_54_379 ();
 sg13g2_decap_8 FILLER_54_386 ();
 sg13g2_decap_8 FILLER_54_393 ();
 sg13g2_decap_8 FILLER_54_400 ();
 sg13g2_fill_2 FILLER_54_407 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_63 ();
 sg13g2_fill_1 FILLER_55_65 ();
 sg13g2_decap_4 FILLER_55_139 ();
 sg13g2_fill_1 FILLER_55_143 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_fill_1 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_373 ();
 sg13g2_decap_8 FILLER_55_380 ();
 sg13g2_decap_8 FILLER_55_387 ();
 sg13g2_decap_8 FILLER_55_394 ();
 sg13g2_decap_8 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_decap_8 FILLER_56_56 ();
 sg13g2_decap_4 FILLER_56_63 ();
 sg13g2_fill_2 FILLER_56_67 ();
 sg13g2_fill_1 FILLER_56_207 ();
 sg13g2_fill_1 FILLER_56_221 ();
 sg13g2_decap_4 FILLER_56_252 ();
 sg13g2_fill_1 FILLER_56_256 ();
 sg13g2_fill_1 FILLER_56_327 ();
 sg13g2_decap_8 FILLER_56_373 ();
 sg13g2_decap_8 FILLER_56_380 ();
 sg13g2_decap_8 FILLER_56_387 ();
 sg13g2_decap_8 FILLER_56_394 ();
 sg13g2_decap_8 FILLER_56_401 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_4 FILLER_57_70 ();
 sg13g2_decap_4 FILLER_57_110 ();
 sg13g2_fill_2 FILLER_57_114 ();
 sg13g2_fill_2 FILLER_57_129 ();
 sg13g2_fill_1 FILLER_57_131 ();
 sg13g2_decap_8 FILLER_57_205 ();
 sg13g2_fill_1 FILLER_57_239 ();
 sg13g2_fill_1 FILLER_57_256 ();
 sg13g2_fill_1 FILLER_57_297 ();
 sg13g2_fill_2 FILLER_57_317 ();
 sg13g2_decap_8 FILLER_57_373 ();
 sg13g2_decap_8 FILLER_57_380 ();
 sg13g2_decap_8 FILLER_57_387 ();
 sg13g2_decap_8 FILLER_57_394 ();
 sg13g2_decap_8 FILLER_57_401 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_fill_1 FILLER_58_63 ();
 sg13g2_decap_4 FILLER_58_128 ();
 sg13g2_fill_2 FILLER_58_145 ();
 sg13g2_fill_1 FILLER_58_147 ();
 sg13g2_fill_2 FILLER_58_175 ();
 sg13g2_fill_1 FILLER_58_177 ();
 sg13g2_decap_4 FILLER_58_205 ();
 sg13g2_fill_2 FILLER_58_209 ();
 sg13g2_fill_2 FILLER_58_238 ();
 sg13g2_fill_1 FILLER_58_240 ();
 sg13g2_decap_8 FILLER_58_379 ();
 sg13g2_decap_8 FILLER_58_386 ();
 sg13g2_decap_8 FILLER_58_393 ();
 sg13g2_decap_8 FILLER_58_400 ();
 sg13g2_fill_2 FILLER_58_407 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_fill_2 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_110 ();
 sg13g2_fill_1 FILLER_59_117 ();
 sg13g2_fill_2 FILLER_59_145 ();
 sg13g2_fill_1 FILLER_59_147 ();
 sg13g2_decap_4 FILLER_59_175 ();
 sg13g2_fill_1 FILLER_59_236 ();
 sg13g2_fill_1 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_346 ();
 sg13g2_decap_8 FILLER_59_384 ();
 sg13g2_decap_8 FILLER_59_391 ();
 sg13g2_decap_8 FILLER_59_398 ();
 sg13g2_decap_4 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_fill_2 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_110 ();
 sg13g2_decap_8 FILLER_60_389 ();
 sg13g2_decap_8 FILLER_60_396 ();
 sg13g2_decap_4 FILLER_60_403 ();
 sg13g2_fill_2 FILLER_60_407 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_fill_2 FILLER_61_49 ();
 sg13g2_decap_4 FILLER_61_106 ();
 sg13g2_fill_1 FILLER_61_110 ();
 sg13g2_fill_2 FILLER_61_121 ();
 sg13g2_fill_1 FILLER_61_123 ();
 sg13g2_fill_1 FILLER_61_137 ();
 sg13g2_decap_4 FILLER_61_158 ();
 sg13g2_decap_8 FILLER_61_204 ();
 sg13g2_fill_1 FILLER_61_211 ();
 sg13g2_decap_8 FILLER_61_399 ();
 sg13g2_fill_2 FILLER_61_406 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_fill_2 FILLER_62_159 ();
 sg13g2_decap_4 FILLER_62_207 ();
 sg13g2_fill_2 FILLER_62_211 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_56 ();
 sg13g2_fill_1 FILLER_63_111 ();
 sg13g2_fill_2 FILLER_63_139 ();
 sg13g2_fill_1 FILLER_63_141 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_fill_2 FILLER_64_70 ();
 sg13g2_decap_4 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_177 ();
 sg13g2_fill_1 FILLER_64_179 ();
 sg13g2_fill_2 FILLER_64_289 ();
 sg13g2_fill_2 FILLER_64_331 ();
 sg13g2_decap_4 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_4 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_125 ();
 sg13g2_fill_1 FILLER_65_132 ();
 sg13g2_fill_2 FILLER_65_293 ();
 sg13g2_fill_1 FILLER_65_317 ();
 sg13g2_fill_1 FILLER_65_360 ();
 sg13g2_decap_8 FILLER_65_394 ();
 sg13g2_decap_8 FILLER_65_401 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_4 FILLER_66_49 ();
 sg13g2_fill_1 FILLER_66_53 ();
 sg13g2_fill_2 FILLER_66_147 ();
 sg13g2_fill_1 FILLER_66_149 ();
 sg13g2_fill_1 FILLER_66_257 ();
 sg13g2_decap_8 FILLER_66_390 ();
 sg13g2_decap_8 FILLER_66_397 ();
 sg13g2_decap_4 FILLER_66_404 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_4 FILLER_67_63 ();
 sg13g2_fill_2 FILLER_67_67 ();
 sg13g2_fill_2 FILLER_67_173 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_393 ();
 sg13g2_decap_8 FILLER_67_400 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_4 FILLER_68_63 ();
 sg13g2_fill_1 FILLER_68_67 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_fill_1 FILLER_68_174 ();
 sg13g2_fill_2 FILLER_68_336 ();
 sg13g2_decap_8 FILLER_68_392 ();
 sg13g2_decap_8 FILLER_68_399 ();
 sg13g2_fill_2 FILLER_68_406 ();
 sg13g2_fill_1 FILLER_68_408 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_4 FILLER_69_70 ();
 sg13g2_fill_2 FILLER_69_74 ();
 sg13g2_decap_4 FILLER_69_139 ();
 sg13g2_fill_1 FILLER_69_143 ();
 sg13g2_fill_1 FILLER_69_157 ();
 sg13g2_fill_2 FILLER_69_198 ();
 sg13g2_fill_1 FILLER_69_200 ();
 sg13g2_decap_8 FILLER_69_384 ();
 sg13g2_decap_8 FILLER_69_391 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_decap_4 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_4 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_fill_1 FILLER_70_176 ();
 sg13g2_fill_2 FILLER_70_202 ();
 sg13g2_fill_1 FILLER_70_237 ();
 sg13g2_fill_2 FILLER_70_269 ();
 sg13g2_decap_8 FILLER_70_382 ();
 sg13g2_decap_8 FILLER_70_389 ();
 sg13g2_decap_8 FILLER_70_396 ();
 sg13g2_decap_4 FILLER_70_403 ();
 sg13g2_fill_2 FILLER_70_407 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_fill_2 FILLER_71_70 ();
 sg13g2_fill_2 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_173 ();
 sg13g2_fill_1 FILLER_71_264 ();
 sg13g2_decap_8 FILLER_71_389 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_decap_4 FILLER_71_403 ();
 sg13g2_fill_2 FILLER_71_407 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_77 ();
 sg13g2_fill_1 FILLER_72_79 ();
 sg13g2_decap_4 FILLER_72_116 ();
 sg13g2_fill_2 FILLER_72_151 ();
 sg13g2_fill_2 FILLER_72_207 ();
 sg13g2_decap_8 FILLER_72_380 ();
 sg13g2_decap_8 FILLER_72_387 ();
 sg13g2_decap_8 FILLER_72_394 ();
 sg13g2_decap_8 FILLER_72_401 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_fill_2 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_144 ();
 sg13g2_fill_1 FILLER_73_182 ();
 sg13g2_decap_8 FILLER_73_375 ();
 sg13g2_decap_8 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_decap_4 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_fill_1 FILLER_74_70 ();
 sg13g2_fill_1 FILLER_74_153 ();
 sg13g2_fill_1 FILLER_74_230 ();
 sg13g2_decap_8 FILLER_74_377 ();
 sg13g2_decap_8 FILLER_74_384 ();
 sg13g2_decap_8 FILLER_74_391 ();
 sg13g2_decap_8 FILLER_74_398 ();
 sg13g2_decap_4 FILLER_74_405 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_63 ();
 sg13g2_fill_2 FILLER_75_167 ();
 sg13g2_fill_1 FILLER_75_169 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_213 ();
 sg13g2_fill_2 FILLER_75_347 ();
 sg13g2_fill_1 FILLER_75_349 ();
 sg13g2_decap_8 FILLER_75_368 ();
 sg13g2_decap_8 FILLER_75_375 ();
 sg13g2_decap_8 FILLER_75_382 ();
 sg13g2_decap_8 FILLER_75_389 ();
 sg13g2_decap_8 FILLER_75_396 ();
 sg13g2_decap_4 FILLER_75_403 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_4 FILLER_76_63 ();
 sg13g2_fill_2 FILLER_76_67 ();
 sg13g2_fill_2 FILLER_76_129 ();
 sg13g2_fill_1 FILLER_76_293 ();
 sg13g2_decap_8 FILLER_76_362 ();
 sg13g2_decap_8 FILLER_76_369 ();
 sg13g2_decap_8 FILLER_76_376 ();
 sg13g2_decap_8 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_390 ();
 sg13g2_decap_8 FILLER_76_397 ();
 sg13g2_decap_4 FILLER_76_404 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_fill_1 FILLER_77_160 ();
 sg13g2_fill_1 FILLER_77_234 ();
 sg13g2_decap_8 FILLER_77_358 ();
 sg13g2_decap_8 FILLER_77_365 ();
 sg13g2_decap_8 FILLER_77_372 ();
 sg13g2_decap_8 FILLER_77_379 ();
 sg13g2_decap_8 FILLER_77_386 ();
 sg13g2_decap_8 FILLER_77_393 ();
 sg13g2_decap_8 FILLER_77_400 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_fill_2 FILLER_78_63 ();
 sg13g2_fill_1 FILLER_78_65 ();
 sg13g2_fill_2 FILLER_78_143 ();
 sg13g2_fill_1 FILLER_78_269 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_decap_8 FILLER_78_355 ();
 sg13g2_decap_8 FILLER_78_362 ();
 sg13g2_decap_8 FILLER_78_369 ();
 sg13g2_decap_8 FILLER_78_376 ();
 sg13g2_decap_8 FILLER_78_383 ();
 sg13g2_decap_8 FILLER_78_390 ();
 sg13g2_decap_8 FILLER_78_397 ();
 sg13g2_decap_4 FILLER_78_404 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_4 FILLER_79_49 ();
 sg13g2_fill_2 FILLER_79_53 ();
 sg13g2_fill_2 FILLER_79_198 ();
 sg13g2_fill_1 FILLER_79_286 ();
 sg13g2_decap_8 FILLER_79_349 ();
 sg13g2_decap_8 FILLER_79_356 ();
 sg13g2_decap_8 FILLER_79_363 ();
 sg13g2_decap_8 FILLER_79_370 ();
 sg13g2_decap_8 FILLER_79_377 ();
 sg13g2_decap_8 FILLER_79_384 ();
 sg13g2_decap_8 FILLER_79_391 ();
 sg13g2_decap_8 FILLER_79_398 ();
 sg13g2_decap_4 FILLER_79_405 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_4 FILLER_80_42 ();
 sg13g2_fill_1 FILLER_80_46 ();
 sg13g2_decap_4 FILLER_80_356 ();
 sg13g2_decap_4 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_372 ();
 sg13g2_decap_8 FILLER_80_379 ();
 sg13g2_decap_8 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_393 ();
 sg13g2_decap_8 FILLER_80_400 ();
 sg13g2_fill_2 FILLER_80_407 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net13;
 assign uio_out[1] = net14;
 assign uio_out[2] = net15;
 assign uio_out[3] = net16;
 assign uio_out[4] = net17;
 assign uio_out[5] = net18;
 assign uio_out[6] = net19;
 assign uio_out[7] = net20;
 assign uo_out[4] = net21;
 assign uo_out[5] = net22;
 assign uo_out[6] = net23;
 assign uo_out[7] = net24;
endmodule
