module tt_um_dranoel06_SAP1 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire clknet_0_clk;
 wire \cpu0.a_reg[0] ;
 wire \cpu0.a_reg[1] ;
 wire \cpu0.a_reg[2] ;
 wire \cpu0.a_reg[3] ;
 wire \cpu0.a_reg[4] ;
 wire \cpu0.a_reg[5] ;
 wire \cpu0.a_reg[6] ;
 wire \cpu0.a_reg[7] ;
 wire \cpu0.b_reg[0] ;
 wire \cpu0.b_reg[1] ;
 wire \cpu0.b_reg[2] ;
 wire \cpu0.b_reg[3] ;
 wire \cpu0.b_reg[4] ;
 wire \cpu0.b_reg[5] ;
 wire \cpu0.b_reg[6] ;
 wire \cpu0.b_reg[7] ;
 wire \cpu0.ir[0] ;
 wire \cpu0.ir[1] ;
 wire \cpu0.ir[2] ;
 wire \cpu0.ir[3] ;
 wire \cpu0.ir[4] ;
 wire \cpu0.ir[5] ;
 wire \cpu0.ir[6] ;
 wire \cpu0.ir[7] ;
 wire \cpu0.mar[0] ;
 wire \cpu0.mar[1] ;
 wire \cpu0.mar[2] ;
 wire \cpu0.mar[3] ;
 wire \cpu0.pc[0] ;
 wire \cpu0.pc[1] ;
 wire \cpu0.pc[2] ;
 wire \cpu0.pc[3] ;
 wire \cpu0.ram[0][0] ;
 wire \cpu0.ram[0][1] ;
 wire \cpu0.ram[0][2] ;
 wire \cpu0.ram[0][3] ;
 wire \cpu0.ram[0][4] ;
 wire \cpu0.ram[0][5] ;
 wire \cpu0.ram[0][6] ;
 wire \cpu0.ram[0][7] ;
 wire \cpu0.ram[10][0] ;
 wire \cpu0.ram[10][1] ;
 wire \cpu0.ram[10][2] ;
 wire \cpu0.ram[10][3] ;
 wire \cpu0.ram[10][4] ;
 wire \cpu0.ram[10][5] ;
 wire \cpu0.ram[10][6] ;
 wire \cpu0.ram[10][7] ;
 wire \cpu0.ram[11][0] ;
 wire \cpu0.ram[11][1] ;
 wire \cpu0.ram[11][2] ;
 wire \cpu0.ram[11][3] ;
 wire \cpu0.ram[11][4] ;
 wire \cpu0.ram[11][5] ;
 wire \cpu0.ram[11][6] ;
 wire \cpu0.ram[11][7] ;
 wire \cpu0.ram[12][0] ;
 wire \cpu0.ram[12][1] ;
 wire \cpu0.ram[12][2] ;
 wire \cpu0.ram[12][3] ;
 wire \cpu0.ram[12][4] ;
 wire \cpu0.ram[12][5] ;
 wire \cpu0.ram[12][6] ;
 wire \cpu0.ram[12][7] ;
 wire \cpu0.ram[13][0] ;
 wire \cpu0.ram[13][1] ;
 wire \cpu0.ram[13][2] ;
 wire \cpu0.ram[13][3] ;
 wire \cpu0.ram[13][4] ;
 wire \cpu0.ram[13][5] ;
 wire \cpu0.ram[13][6] ;
 wire \cpu0.ram[13][7] ;
 wire \cpu0.ram[14][0] ;
 wire \cpu0.ram[14][1] ;
 wire \cpu0.ram[14][2] ;
 wire \cpu0.ram[14][3] ;
 wire \cpu0.ram[14][4] ;
 wire \cpu0.ram[14][5] ;
 wire \cpu0.ram[14][6] ;
 wire \cpu0.ram[14][7] ;
 wire \cpu0.ram[15][0] ;
 wire \cpu0.ram[15][1] ;
 wire \cpu0.ram[15][2] ;
 wire \cpu0.ram[15][3] ;
 wire \cpu0.ram[15][4] ;
 wire \cpu0.ram[15][5] ;
 wire \cpu0.ram[15][6] ;
 wire \cpu0.ram[15][7] ;
 wire \cpu0.ram[1][0] ;
 wire \cpu0.ram[1][1] ;
 wire \cpu0.ram[1][2] ;
 wire \cpu0.ram[1][3] ;
 wire \cpu0.ram[1][4] ;
 wire \cpu0.ram[1][5] ;
 wire \cpu0.ram[1][6] ;
 wire \cpu0.ram[1][7] ;
 wire \cpu0.ram[2][0] ;
 wire \cpu0.ram[2][1] ;
 wire \cpu0.ram[2][2] ;
 wire \cpu0.ram[2][3] ;
 wire \cpu0.ram[2][4] ;
 wire \cpu0.ram[2][5] ;
 wire \cpu0.ram[2][6] ;
 wire \cpu0.ram[2][7] ;
 wire \cpu0.ram[3][0] ;
 wire \cpu0.ram[3][1] ;
 wire \cpu0.ram[3][2] ;
 wire \cpu0.ram[3][3] ;
 wire \cpu0.ram[3][4] ;
 wire \cpu0.ram[3][5] ;
 wire \cpu0.ram[3][6] ;
 wire \cpu0.ram[3][7] ;
 wire \cpu0.ram[4][0] ;
 wire \cpu0.ram[4][1] ;
 wire \cpu0.ram[4][2] ;
 wire \cpu0.ram[4][3] ;
 wire \cpu0.ram[4][4] ;
 wire \cpu0.ram[4][5] ;
 wire \cpu0.ram[4][6] ;
 wire \cpu0.ram[4][7] ;
 wire \cpu0.ram[5][0] ;
 wire \cpu0.ram[5][1] ;
 wire \cpu0.ram[5][2] ;
 wire \cpu0.ram[5][3] ;
 wire \cpu0.ram[5][4] ;
 wire \cpu0.ram[5][5] ;
 wire \cpu0.ram[5][6] ;
 wire \cpu0.ram[5][7] ;
 wire \cpu0.ram[6][0] ;
 wire \cpu0.ram[6][1] ;
 wire \cpu0.ram[6][2] ;
 wire \cpu0.ram[6][3] ;
 wire \cpu0.ram[6][4] ;
 wire \cpu0.ram[6][5] ;
 wire \cpu0.ram[6][6] ;
 wire \cpu0.ram[6][7] ;
 wire \cpu0.ram[7][0] ;
 wire \cpu0.ram[7][1] ;
 wire \cpu0.ram[7][2] ;
 wire \cpu0.ram[7][3] ;
 wire \cpu0.ram[7][4] ;
 wire \cpu0.ram[7][5] ;
 wire \cpu0.ram[7][6] ;
 wire \cpu0.ram[7][7] ;
 wire \cpu0.ram[8][0] ;
 wire \cpu0.ram[8][1] ;
 wire \cpu0.ram[8][2] ;
 wire \cpu0.ram[8][3] ;
 wire \cpu0.ram[8][4] ;
 wire \cpu0.ram[8][5] ;
 wire \cpu0.ram[8][6] ;
 wire \cpu0.ram[8][7] ;
 wire \cpu0.ram[9][0] ;
 wire \cpu0.ram[9][1] ;
 wire \cpu0.ram[9][2] ;
 wire \cpu0.ram[9][3] ;
 wire \cpu0.ram[9][4] ;
 wire \cpu0.ram[9][5] ;
 wire \cpu0.ram[9][6] ;
 wire \cpu0.ram[9][7] ;
 wire \cpu0.step[0] ;
 wire \cpu0.step[1] ;
 wire \cpu0.step[2] ;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;

 sg13g2_inv_1 _0778_ (.Y(_0179_),
    .A(\cpu0.a_reg[1] ));
 sg13g2_inv_1 _0779_ (.Y(_0180_),
    .A(\cpu0.ir[7] ));
 sg13g2_inv_1 _0780_ (.Y(_0181_),
    .A(net468));
 sg13g2_inv_1 _0781_ (.Y(_0182_),
    .A(net207));
 sg13g2_inv_1 _0782_ (.Y(_0183_),
    .A(net188));
 sg13g2_inv_1 _0783_ (.Y(_0184_),
    .A(net180));
 sg13g2_inv_1 _0784_ (.Y(_0185_),
    .A(\cpu0.ram[9][1] ));
 sg13g2_inv_1 _0785_ (.Y(_0186_),
    .A(net283));
 sg13g2_inv_1 _0786_ (.Y(_0187_),
    .A(net288));
 sg13g2_inv_1 _0787_ (.Y(_0188_),
    .A(\cpu0.ram[1][2] ));
 sg13g2_inv_1 _0788_ (.Y(_0189_),
    .A(net286));
 sg13g2_inv_1 _0789_ (.Y(_0190_),
    .A(net285));
 sg13g2_inv_1 _0790_ (.Y(_0191_),
    .A(\cpu0.ram[13][2] ));
 sg13g2_inv_1 _0791_ (.Y(_0192_),
    .A(\cpu0.ram[5][3] ));
 sg13g2_inv_1 _0792_ (.Y(_0193_),
    .A(\cpu0.ram[7][3] ));
 sg13g2_inv_1 _0793_ (.Y(_0194_),
    .A(net281));
 sg13g2_inv_1 _0794_ (.Y(_0195_),
    .A(net280));
 sg13g2_inv_1 _0795_ (.Y(_0196_),
    .A(net284));
 sg13g2_inv_1 _0796_ (.Y(_0197_),
    .A(\cpu0.ram[13][4] ));
 sg13g2_inv_1 _0797_ (.Y(_0198_),
    .A(\cpu0.ram[15][5] ));
 sg13g2_inv_1 _0798_ (.Y(_0199_),
    .A(\cpu0.ram[13][6] ));
 sg13g2_inv_1 _0799_ (.Y(_0200_),
    .A(\cpu0.ram[13][7] ));
 sg13g2_nand2b_1 _0800_ (.Y(_0201_),
    .B(\cpu0.ir[6] ),
    .A_N(\cpu0.ir[7] ));
 sg13g2_nand2b_1 _0801_ (.Y(_0202_),
    .B(\cpu0.ir[4] ),
    .A_N(\cpu0.ir[5] ));
 sg13g2_nor4_1 _0802_ (.A(\cpu0.step[0] ),
    .B(\cpu0.step[1] ),
    .C(_0181_),
    .D(_0202_),
    .Y(_0203_));
 sg13g2_nand4_1 _0803_ (.B(\cpu0.ir[6] ),
    .C(net207),
    .A(_0180_),
    .Y(_0204_),
    .D(_0203_));
 sg13g2_nor2b_2 _0804_ (.A(net13),
    .B_N(_0204_),
    .Y(_0205_));
 sg13g2_nor2_1 _0805_ (.A(net13),
    .B(_0204_),
    .Y(_0206_));
 sg13g2_mux2_1 _0806_ (.A0(net9),
    .A1(\cpu0.mar[0] ),
    .S(net168),
    .X(_0207_));
 sg13g2_nor2b_2 _0807_ (.A(_0205_),
    .B_N(_0207_),
    .Y(_0208_));
 sg13g2_nor2b_1 _0808_ (.A(net168),
    .B_N(net10),
    .Y(_0209_));
 sg13g2_a21oi_2 _0809_ (.B1(_0209_),
    .Y(_0210_),
    .A2(net168),
    .A1(\cpu0.mar[1] ));
 sg13g2_a21o_2 _0810_ (.A2(net168),
    .A1(\cpu0.mar[1] ),
    .B1(_0209_),
    .X(_0211_));
 sg13g2_nand2_1 _0811_ (.Y(_0212_),
    .A(_0208_),
    .B(_0210_));
 sg13g2_mux2_1 _0812_ (.A0(net11),
    .A1(\cpu0.mar[2] ),
    .S(net168),
    .X(_0213_));
 sg13g2_mux2_1 _0813_ (.A0(net12),
    .A1(\cpu0.mar[3] ),
    .S(net168),
    .X(_0214_));
 sg13g2_nand2b_1 _0814_ (.Y(_0215_),
    .B(_0213_),
    .A_N(_0214_));
 sg13g2_or2_1 _0815_ (.X(_0216_),
    .B(_0215_),
    .A(_0212_));
 sg13g2_nand2_1 _0816_ (.Y(_0217_),
    .A(net450),
    .B(_0181_));
 sg13g2_nand2b_2 _0817_ (.Y(_0218_),
    .B(net450),
    .A_N(\cpu0.step[1] ));
 sg13g2_nor3_2 _0818_ (.A(\cpu0.step[2] ),
    .B(net202),
    .C(_0218_),
    .Y(_0219_));
 sg13g2_nand2_1 _0819_ (.Y(_0220_),
    .A(net450),
    .B(net472));
 sg13g2_nor2_1 _0820_ (.A(\cpu0.step[2] ),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_nor3_1 _0821_ (.A(net468),
    .B(net203),
    .C(_0220_),
    .Y(_0222_));
 sg13g2_nand2_1 _0822_ (.Y(_0223_),
    .A(net207),
    .B(_0221_));
 sg13g2_nor3_1 _0823_ (.A(\cpu0.a_reg[1] ),
    .B(\cpu0.a_reg[0] ),
    .C(\cpu0.ir[6] ),
    .Y(_0224_));
 sg13g2_nor2_1 _0824_ (.A(\cpu0.a_reg[7] ),
    .B(\cpu0.a_reg[6] ),
    .Y(_0225_));
 sg13g2_nor4_1 _0825_ (.A(\cpu0.a_reg[5] ),
    .B(\cpu0.a_reg[4] ),
    .C(\cpu0.a_reg[3] ),
    .D(\cpu0.a_reg[2] ),
    .Y(_0226_));
 sg13g2_nand3_1 _0826_ (.B(_0225_),
    .C(_0226_),
    .A(_0224_),
    .Y(_0227_));
 sg13g2_nor2_1 _0827_ (.A(\cpu0.ir[7] ),
    .B(\cpu0.ir[6] ),
    .Y(_0228_));
 sg13g2_nor2_1 _0828_ (.A(\cpu0.ir[5] ),
    .B(\cpu0.ir[4] ),
    .Y(_0229_));
 sg13g2_nand3b_1 _0829_ (.B(_0229_),
    .C(_0221_),
    .Y(_0230_),
    .A_N(_0228_));
 sg13g2_a21oi_1 _0830_ (.A1(\cpu0.ir[7] ),
    .A2(_0227_),
    .Y(_0231_),
    .B1(_0230_));
 sg13g2_nand2_2 _0831_ (.Y(_0232_),
    .A(\cpu0.ir[5] ),
    .B(\cpu0.ir[4] ));
 sg13g2_nor2_1 _0832_ (.A(\cpu0.ir[6] ),
    .B(_0232_),
    .Y(_0233_));
 sg13g2_nor3_1 _0833_ (.A(\cpu0.ir[7] ),
    .B(_0229_),
    .C(_0233_),
    .Y(_0234_));
 sg13g2_nor2_1 _0834_ (.A(_0231_),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_nor2_2 _0835_ (.A(_0223_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_nand2_1 _0836_ (.Y(_0237_),
    .A(\cpu0.ir[0] ),
    .B(_0236_));
 sg13g2_nor4_2 _0837_ (.A(\cpu0.ir[7] ),
    .B(\cpu0.ir[6] ),
    .C(_0223_),
    .Y(_0238_),
    .D(_0232_));
 sg13g2_nand4_1 _0838_ (.B(\cpu0.ir[4] ),
    .C(_0222_),
    .A(\cpu0.ir[5] ),
    .Y(_0239_),
    .D(_0228_));
 sg13g2_nand2_2 _0839_ (.Y(_0240_),
    .A(_0204_),
    .B(_0239_));
 sg13g2_nor2b_1 _0840_ (.A(\cpu0.ir[4] ),
    .B_N(\cpu0.ir[5] ),
    .Y(_0241_));
 sg13g2_nor2_1 _0841_ (.A(_0201_),
    .B(_0232_),
    .Y(_0242_));
 sg13g2_a21oi_1 _0842_ (.A1(_0228_),
    .A2(_0241_),
    .Y(_0243_),
    .B1(_0242_));
 sg13g2_nand2b_2 _0843_ (.Y(_0244_),
    .B(\cpu0.step[1] ),
    .A_N(net450));
 sg13g2_nand2_1 _0844_ (.Y(_0245_),
    .A(net468),
    .B(net207));
 sg13g2_nor3_2 _0845_ (.A(_0243_),
    .B(_0244_),
    .C(_0245_),
    .Y(_0246_));
 sg13g2_nor4_1 _0846_ (.A(net450),
    .B(\cpu0.step[1] ),
    .C(_0181_),
    .D(_0243_),
    .Y(_0247_));
 sg13g2_nand2_1 _0847_ (.Y(_0248_),
    .A(net204),
    .B(_0247_));
 sg13g2_nor2_2 _0848_ (.A(net473),
    .B(_0244_),
    .Y(_0249_));
 sg13g2_nor3_2 _0849_ (.A(net473),
    .B(net202),
    .C(_0244_),
    .Y(_0250_));
 sg13g2_nand2_2 _0850_ (.Y(_0251_),
    .A(net207),
    .B(_0249_));
 sg13g2_nand3_1 _0851_ (.B(_0203_),
    .C(_0228_),
    .A(net207),
    .Y(_0252_));
 sg13g2_and3_2 _0852_ (.X(_0253_),
    .A(net166),
    .B(net171),
    .C(_0252_));
 sg13g2_nand3_1 _0853_ (.B(net171),
    .C(_0252_),
    .A(net166),
    .Y(_0254_));
 sg13g2_nand2b_1 _0854_ (.Y(_0255_),
    .B(\cpu0.b_reg[0] ),
    .A_N(\cpu0.a_reg[0] ));
 sg13g2_xor2_1 _0855_ (.B(\cpu0.a_reg[0] ),
    .A(\cpu0.b_reg[0] ),
    .X(_0256_));
 sg13g2_a221oi_1 _0856_ (.B2(_0256_),
    .C1(_0254_),
    .B1(net167),
    .A1(\cpu0.a_reg[0] ),
    .Y(_0257_),
    .A2(_0240_));
 sg13g2_mux2_1 _0857_ (.A0(\cpu0.ram[12][0] ),
    .A1(\cpu0.ram[13][0] ),
    .S(net198),
    .X(_0258_));
 sg13g2_nand2_1 _0858_ (.Y(_0259_),
    .A(net174),
    .B(_0258_));
 sg13g2_mux2_1 _0859_ (.A0(\cpu0.ram[14][0] ),
    .A1(\cpu0.ram[15][0] ),
    .S(net200),
    .X(_0260_));
 sg13g2_a21oi_1 _0860_ (.A1(net187),
    .A2(_0260_),
    .Y(_0261_),
    .B1(_0184_));
 sg13g2_mux4_1 _0861_ (.S0(net191),
    .A0(\cpu0.ram[8][0] ),
    .A1(\cpu0.ram[9][0] ),
    .A2(\cpu0.ram[10][0] ),
    .A3(\cpu0.ram[11][0] ),
    .S1(net183),
    .X(_0262_));
 sg13g2_o21ai_1 _0862_ (.B1(net175),
    .Y(_0263_),
    .A1(net177),
    .A2(_0262_));
 sg13g2_a21oi_1 _0863_ (.A1(_0259_),
    .A2(_0261_),
    .Y(_0264_),
    .B1(_0263_));
 sg13g2_mux4_1 _0864_ (.S0(net192),
    .A0(\cpu0.ram[0][0] ),
    .A1(\cpu0.ram[1][0] ),
    .A2(\cpu0.ram[2][0] ),
    .A3(\cpu0.ram[3][0] ),
    .S1(net185),
    .X(_0265_));
 sg13g2_nor2_1 _0865_ (.A(net179),
    .B(_0265_),
    .Y(_0266_));
 sg13g2_mux2_1 _0866_ (.A0(\cpu0.ram[4][0] ),
    .A1(\cpu0.ram[5][0] ),
    .S(net198),
    .X(_0267_));
 sg13g2_nor2b_1 _0867_ (.A(\cpu0.ram[7][0] ),
    .B_N(net194),
    .Y(_0268_));
 sg13g2_o21ai_1 _0868_ (.B1(net187),
    .Y(_0269_),
    .A1(net194),
    .A2(\cpu0.ram[6][0] ));
 sg13g2_o21ai_1 _0869_ (.B1(net177),
    .Y(_0270_),
    .A1(_0268_),
    .A2(_0269_));
 sg13g2_a21oi_1 _0870_ (.A1(net173),
    .A2(_0267_),
    .Y(_0271_),
    .B1(_0270_));
 sg13g2_nor3_1 _0871_ (.A(net175),
    .B(_0266_),
    .C(_0271_),
    .Y(_0272_));
 sg13g2_nor2_1 _0872_ (.A(_0264_),
    .B(_0272_),
    .Y(_0273_));
 sg13g2_a221oi_1 _0873_ (.B2(net161),
    .C1(net172),
    .B1(_0273_),
    .A1(_0237_),
    .Y(_0274_),
    .A2(_0257_));
 sg13g2_a21o_2 _0874_ (.A2(net172),
    .A1(net442),
    .B1(_0274_),
    .X(_0275_));
 sg13g2_inv_4 _0875_ (.A(_0275_),
    .Y(_0276_));
 sg13g2_nor2_1 _0876_ (.A(net1),
    .B(net169),
    .Y(_0277_));
 sg13g2_a21oi_2 _0877_ (.B1(_0277_),
    .Y(_0278_),
    .A2(_0276_),
    .A1(net169));
 sg13g2_mux2_1 _0878_ (.A0(net150),
    .A1(net377),
    .S(net159),
    .X(_0004_));
 sg13g2_or4_1 _0879_ (.A(_0201_),
    .B(_0232_),
    .C(_0244_),
    .D(_0245_),
    .X(_0279_));
 sg13g2_nand3_1 _0880_ (.B(\cpu0.b_reg[0] ),
    .C(_0279_),
    .A(\cpu0.b_reg[1] ),
    .Y(_0280_));
 sg13g2_a21o_1 _0881_ (.A2(_0279_),
    .A1(\cpu0.b_reg[0] ),
    .B1(\cpu0.b_reg[1] ),
    .X(_0281_));
 sg13g2_a21oi_1 _0882_ (.A1(_0280_),
    .A2(_0281_),
    .Y(_0282_),
    .B1(_0179_));
 sg13g2_nand3_1 _0883_ (.B(_0280_),
    .C(_0281_),
    .A(_0179_),
    .Y(_0283_));
 sg13g2_nand2b_1 _0884_ (.Y(_0284_),
    .B(_0283_),
    .A_N(_0282_));
 sg13g2_xnor2_1 _0885_ (.Y(_0285_),
    .A(_0255_),
    .B(_0284_));
 sg13g2_a21oi_1 _0886_ (.A1(\cpu0.ir[1] ),
    .A2(_0236_),
    .Y(_0286_),
    .B1(net161));
 sg13g2_a22oi_1 _0887_ (.Y(_0287_),
    .B1(net167),
    .B2(_0285_),
    .A2(_0240_),
    .A1(\cpu0.a_reg[1] ));
 sg13g2_nand2b_1 _0888_ (.Y(_0288_),
    .B(net197),
    .A_N(\cpu0.ram[13][1] ));
 sg13g2_o21ai_1 _0889_ (.B1(_0288_),
    .Y(_0289_),
    .A1(net197),
    .A2(\cpu0.ram[12][1] ));
 sg13g2_o21ai_1 _0890_ (.B1(net188),
    .Y(_0290_),
    .A1(net200),
    .A2(\cpu0.ram[14][1] ));
 sg13g2_a21oi_1 _0891_ (.A1(net200),
    .A2(_0187_),
    .Y(_0291_),
    .B1(_0290_));
 sg13g2_o21ai_1 _0892_ (.B1(net182),
    .Y(_0292_),
    .A1(net187),
    .A2(_0289_));
 sg13g2_o21ai_1 _0893_ (.B1(net173),
    .Y(_0293_),
    .A1(net189),
    .A2(\cpu0.ram[8][1] ));
 sg13g2_a21oi_1 _0894_ (.A1(net190),
    .A2(_0185_),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_o21ai_1 _0895_ (.B1(net184),
    .Y(_0295_),
    .A1(net190),
    .A2(\cpu0.ram[10][1] ));
 sg13g2_a21oi_1 _0896_ (.A1(net190),
    .A2(_0186_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_nor3_1 _0897_ (.A(net177),
    .B(_0294_),
    .C(_0296_),
    .Y(_0297_));
 sg13g2_o21ai_1 _0898_ (.B1(net176),
    .Y(_0298_),
    .A1(_0291_),
    .A2(_0292_));
 sg13g2_nor2_1 _0899_ (.A(_0297_),
    .B(_0298_),
    .Y(_0299_));
 sg13g2_mux4_1 _0900_ (.S0(net192),
    .A0(\cpu0.ram[0][1] ),
    .A1(\cpu0.ram[1][1] ),
    .A2(\cpu0.ram[2][1] ),
    .A3(\cpu0.ram[3][1] ),
    .S1(net185),
    .X(_0300_));
 sg13g2_nor2_1 _0901_ (.A(net179),
    .B(_0300_),
    .Y(_0301_));
 sg13g2_mux2_1 _0902_ (.A0(\cpu0.ram[4][1] ),
    .A1(\cpu0.ram[5][1] ),
    .S(net198),
    .X(_0302_));
 sg13g2_nor2b_1 _0903_ (.A(\cpu0.ram[7][1] ),
    .B_N(net194),
    .Y(_0303_));
 sg13g2_o21ai_1 _0904_ (.B1(net187),
    .Y(_0304_),
    .A1(net194),
    .A2(\cpu0.ram[6][1] ));
 sg13g2_o21ai_1 _0905_ (.B1(net177),
    .Y(_0305_),
    .A1(_0303_),
    .A2(_0304_));
 sg13g2_a21oi_1 _0906_ (.A1(net173),
    .A2(_0302_),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_nor3_1 _0907_ (.A(net175),
    .B(_0301_),
    .C(_0306_),
    .Y(_0307_));
 sg13g2_nor2_1 _0908_ (.A(_0299_),
    .B(_0307_),
    .Y(_0308_));
 sg13g2_a221oi_1 _0909_ (.B2(net161),
    .C1(net172),
    .B1(_0308_),
    .A1(_0286_),
    .Y(_0309_),
    .A2(_0287_));
 sg13g2_a21oi_2 _0910_ (.B1(_0309_),
    .Y(_0310_),
    .A2(net172),
    .A1(net457));
 sg13g2_nor2_1 _0911_ (.A(net2),
    .B(net169),
    .Y(_0311_));
 sg13g2_a21oi_1 _0912_ (.A1(net169),
    .A2(_0310_),
    .Y(_0312_),
    .B1(_0311_));
 sg13g2_mux2_1 _0913_ (.A0(net154),
    .A1(net416),
    .S(net159),
    .X(_0005_));
 sg13g2_a21o_1 _0914_ (.A2(_0283_),
    .A1(_0255_),
    .B1(_0282_),
    .X(_0313_));
 sg13g2_or2_1 _0915_ (.X(_0314_),
    .B(\cpu0.b_reg[0] ),
    .A(\cpu0.b_reg[1] ));
 sg13g2_nand2_1 _0916_ (.Y(_0315_),
    .A(_0279_),
    .B(_0314_));
 sg13g2_xnor2_1 _0917_ (.Y(_0316_),
    .A(\cpu0.b_reg[2] ),
    .B(_0315_));
 sg13g2_nand2b_1 _0918_ (.Y(_0317_),
    .B(\cpu0.a_reg[2] ),
    .A_N(_0316_));
 sg13g2_xnor2_1 _0919_ (.Y(_0318_),
    .A(\cpu0.a_reg[2] ),
    .B(_0316_));
 sg13g2_nand2_1 _0920_ (.Y(_0319_),
    .A(_0313_),
    .B(_0318_));
 sg13g2_o21ai_1 _0921_ (.B1(net167),
    .Y(_0320_),
    .A1(_0313_),
    .A2(_0318_));
 sg13g2_nand2b_1 _0922_ (.Y(_0321_),
    .B(_0319_),
    .A_N(_0320_));
 sg13g2_a221oi_1 _0923_ (.B2(\cpu0.a_reg[2] ),
    .C1(net161),
    .B1(_0240_),
    .A1(\cpu0.ir[2] ),
    .Y(_0322_),
    .A2(_0236_));
 sg13g2_a21oi_1 _0924_ (.A1(net192),
    .A2(_0188_),
    .Y(_0323_),
    .B1(net185));
 sg13g2_o21ai_1 _0925_ (.B1(_0323_),
    .Y(_0324_),
    .A1(net193),
    .A2(\cpu0.ram[0][2] ));
 sg13g2_o21ai_1 _0926_ (.B1(net186),
    .Y(_0325_),
    .A1(net193),
    .A2(\cpu0.ram[2][2] ));
 sg13g2_a21oi_1 _0927_ (.A1(net193),
    .A2(_0189_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_nor2_1 _0928_ (.A(net179),
    .B(_0326_),
    .Y(_0327_));
 sg13g2_o21ai_1 _0929_ (.B1(net174),
    .Y(_0328_),
    .A1(net198),
    .A2(\cpu0.ram[4][2] ));
 sg13g2_a21oi_1 _0930_ (.A1(net198),
    .A2(_0190_),
    .Y(_0329_),
    .B1(_0328_));
 sg13g2_nor2b_1 _0931_ (.A(\cpu0.ram[7][2] ),
    .B_N(net194),
    .Y(_0330_));
 sg13g2_o21ai_1 _0932_ (.B1(net187),
    .Y(_0331_),
    .A1(net194),
    .A2(\cpu0.ram[6][2] ));
 sg13g2_o21ai_1 _0933_ (.B1(net178),
    .Y(_0332_),
    .A1(_0330_),
    .A2(_0331_));
 sg13g2_or2_1 _0934_ (.X(_0333_),
    .B(_0332_),
    .A(_0329_));
 sg13g2_a21oi_1 _0935_ (.A1(_0324_),
    .A2(_0327_),
    .Y(_0334_),
    .B1(net176));
 sg13g2_mux4_1 _0936_ (.S0(net189),
    .A0(\cpu0.ram[8][2] ),
    .A1(\cpu0.ram[9][2] ),
    .A2(\cpu0.ram[10][2] ),
    .A3(\cpu0.ram[11][2] ),
    .S1(net184),
    .X(_0335_));
 sg13g2_nor2_1 _0937_ (.A(net177),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_o21ai_1 _0938_ (.B1(net174),
    .Y(_0337_),
    .A1(net198),
    .A2(\cpu0.ram[12][2] ));
 sg13g2_a21oi_1 _0939_ (.A1(net198),
    .A2(_0191_),
    .Y(_0338_),
    .B1(_0337_));
 sg13g2_nor2b_1 _0940_ (.A(\cpu0.ram[15][2] ),
    .B_N(net199),
    .Y(_0339_));
 sg13g2_o21ai_1 _0941_ (.B1(net187),
    .Y(_0340_),
    .A1(net197),
    .A2(\cpu0.ram[14][2] ));
 sg13g2_o21ai_1 _0942_ (.B1(net182),
    .Y(_0341_),
    .A1(_0339_),
    .A2(_0340_));
 sg13g2_o21ai_1 _0943_ (.B1(net176),
    .Y(_0342_),
    .A1(_0338_),
    .A2(_0341_));
 sg13g2_nor2_1 _0944_ (.A(_0336_),
    .B(_0342_),
    .Y(_0343_));
 sg13g2_a21oi_1 _0945_ (.A1(_0333_),
    .A2(_0334_),
    .Y(_0344_),
    .B1(_0343_));
 sg13g2_a221oi_1 _0946_ (.B2(net161),
    .C1(net172),
    .B1(_0344_),
    .A1(_0321_),
    .Y(_0345_),
    .A2(_0322_));
 sg13g2_a21oi_2 _0947_ (.B1(_0345_),
    .Y(_0346_),
    .A2(net172),
    .A1(net459));
 sg13g2_nor2_1 _0948_ (.A(net3),
    .B(net169),
    .Y(_0347_));
 sg13g2_a21oi_1 _0949_ (.A1(net169),
    .A2(_0346_),
    .Y(_0348_),
    .B1(_0347_));
 sg13g2_nor2_1 _0950_ (.A(net159),
    .B(net152),
    .Y(_0349_));
 sg13g2_a21oi_1 _0951_ (.A1(_0190_),
    .A2(net159),
    .Y(_0006_),
    .B1(_0349_));
 sg13g2_a221oi_1 _0952_ (.B2(\cpu0.a_reg[3] ),
    .C1(net161),
    .B1(_0240_),
    .A1(\cpu0.ir[3] ),
    .Y(_0350_),
    .A2(_0236_));
 sg13g2_o21ai_1 _0953_ (.B1(_0279_),
    .Y(_0351_),
    .A1(\cpu0.b_reg[2] ),
    .A2(_0314_));
 sg13g2_nand2_1 _0954_ (.Y(_0352_),
    .A(\cpu0.b_reg[3] ),
    .B(_0279_));
 sg13g2_xor2_1 _0955_ (.B(_0351_),
    .A(\cpu0.b_reg[3] ),
    .X(_0353_));
 sg13g2_nand2_1 _0956_ (.Y(_0354_),
    .A(\cpu0.a_reg[3] ),
    .B(_0353_));
 sg13g2_xnor2_1 _0957_ (.Y(_0355_),
    .A(\cpu0.a_reg[3] ),
    .B(_0353_));
 sg13g2_nand3_1 _0958_ (.B(_0319_),
    .C(_0355_),
    .A(_0317_),
    .Y(_0356_));
 sg13g2_a21o_2 _0959_ (.A2(_0319_),
    .A1(_0317_),
    .B1(_0355_),
    .X(_0357_));
 sg13g2_nand3_1 _0960_ (.B(_0356_),
    .C(_0357_),
    .A(net167),
    .Y(_0358_));
 sg13g2_mux4_1 _0961_ (.S0(net192),
    .A0(\cpu0.ram[0][3] ),
    .A1(\cpu0.ram[1][3] ),
    .A2(\cpu0.ram[2][3] ),
    .A3(\cpu0.ram[3][3] ),
    .S1(net185),
    .X(_0359_));
 sg13g2_nand2b_1 _0962_ (.Y(_0360_),
    .B(_0184_),
    .A_N(_0359_));
 sg13g2_a21oi_1 _0963_ (.A1(net197),
    .A2(_0192_),
    .Y(_0361_),
    .B1(net188));
 sg13g2_o21ai_1 _0964_ (.B1(_0361_),
    .Y(_0362_),
    .A1(net195),
    .A2(\cpu0.ram[4][3] ));
 sg13g2_o21ai_1 _0965_ (.B1(net184),
    .Y(_0363_),
    .A1(net190),
    .A2(\cpu0.ram[6][3] ));
 sg13g2_a21oi_1 _0966_ (.A1(net195),
    .A2(_0193_),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_nor2_1 _0967_ (.A(_0184_),
    .B(_0364_),
    .Y(_0365_));
 sg13g2_a21oi_1 _0968_ (.A1(_0362_),
    .A2(_0365_),
    .Y(_0366_),
    .B1(net175));
 sg13g2_a21oi_1 _0969_ (.A1(net190),
    .A2(_0194_),
    .Y(_0367_),
    .B1(net184));
 sg13g2_o21ai_1 _0970_ (.B1(_0367_),
    .Y(_0368_),
    .A1(net190),
    .A2(\cpu0.ram[8][3] ));
 sg13g2_o21ai_1 _0971_ (.B1(net183),
    .Y(_0369_),
    .A1(net191),
    .A2(\cpu0.ram[10][3] ));
 sg13g2_a21oi_1 _0972_ (.A1(net190),
    .A2(_0195_),
    .Y(_0370_),
    .B1(_0369_));
 sg13g2_nor2_1 _0973_ (.A(net179),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_o21ai_1 _0974_ (.B1(net174),
    .Y(_0372_),
    .A1(net199),
    .A2(\cpu0.ram[12][3] ));
 sg13g2_a21oi_1 _0975_ (.A1(net199),
    .A2(_0196_),
    .Y(_0373_),
    .B1(_0372_));
 sg13g2_nor2b_1 _0976_ (.A(\cpu0.ram[15][3] ),
    .B_N(net197),
    .Y(_0374_));
 sg13g2_o21ai_1 _0977_ (.B1(net188),
    .Y(_0375_),
    .A1(net197),
    .A2(\cpu0.ram[14][3] ));
 sg13g2_o21ai_1 _0978_ (.B1(net182),
    .Y(_0376_),
    .A1(_0374_),
    .A2(_0375_));
 sg13g2_o21ai_1 _0979_ (.B1(net176),
    .Y(_0377_),
    .A1(_0373_),
    .A2(_0376_));
 sg13g2_a21oi_1 _0980_ (.A1(_0368_),
    .A2(_0371_),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_a21oi_1 _0981_ (.A1(_0360_),
    .A2(_0366_),
    .Y(_0379_),
    .B1(_0378_));
 sg13g2_a221oi_1 _0982_ (.B2(net161),
    .C1(net172),
    .B1(_0379_),
    .A1(_0350_),
    .Y(_0380_),
    .A2(_0358_));
 sg13g2_a21oi_2 _0983_ (.B1(_0380_),
    .Y(_0381_),
    .A2(net172),
    .A1(net461));
 sg13g2_nor2_1 _0984_ (.A(net4),
    .B(net169),
    .Y(_0382_));
 sg13g2_a21oi_2 _0985_ (.B1(_0382_),
    .Y(_0383_),
    .A2(_0381_),
    .A1(net170));
 sg13g2_mux2_1 _0986_ (.A0(net148),
    .A1(net333),
    .S(_0216_),
    .X(_0007_));
 sg13g2_nor2_1 _0987_ (.A(net5),
    .B(net169),
    .Y(_0384_));
 sg13g2_nand2_1 _0988_ (.Y(_0385_),
    .A(_0351_),
    .B(_0352_));
 sg13g2_xor2_1 _0989_ (.B(_0385_),
    .A(\cpu0.b_reg[4] ),
    .X(_0386_));
 sg13g2_nand2b_1 _0990_ (.Y(_0387_),
    .B(\cpu0.a_reg[4] ),
    .A_N(_0386_));
 sg13g2_xor2_1 _0991_ (.B(_0386_),
    .A(\cpu0.a_reg[4] ),
    .X(_0388_));
 sg13g2_a21o_1 _0992_ (.A2(_0357_),
    .A1(_0354_),
    .B1(_0388_),
    .X(_0389_));
 sg13g2_nand3_1 _0993_ (.B(_0357_),
    .C(_0388_),
    .A(_0354_),
    .Y(_0390_));
 sg13g2_and2_1 _0994_ (.A(net167),
    .B(_0390_),
    .X(_0391_));
 sg13g2_a22oi_1 _0995_ (.Y(_0392_),
    .B1(_0389_),
    .B2(_0391_),
    .A2(_0240_),
    .A1(\cpu0.a_reg[4] ));
 sg13g2_o21ai_1 _0996_ (.B1(net174),
    .Y(_0393_),
    .A1(net197),
    .A2(\cpu0.ram[12][4] ));
 sg13g2_a21oi_1 _0997_ (.A1(net197),
    .A2(_0197_),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_nor2b_1 _0998_ (.A(\cpu0.ram[15][4] ),
    .B_N(net200),
    .Y(_0395_));
 sg13g2_o21ai_1 _0999_ (.B1(net188),
    .Y(_0396_),
    .A1(net201),
    .A2(\cpu0.ram[14][4] ));
 sg13g2_o21ai_1 _1000_ (.B1(net182),
    .Y(_0397_),
    .A1(_0395_),
    .A2(_0396_));
 sg13g2_mux4_1 _1001_ (.S0(net191),
    .A0(\cpu0.ram[8][4] ),
    .A1(\cpu0.ram[9][4] ),
    .A2(\cpu0.ram[10][4] ),
    .A3(\cpu0.ram[11][4] ),
    .S1(net183),
    .X(_0398_));
 sg13g2_nor2_1 _1002_ (.A(net180),
    .B(_0398_),
    .Y(_0399_));
 sg13g2_o21ai_1 _1003_ (.B1(_0003_),
    .Y(_0400_),
    .A1(_0394_),
    .A2(_0397_));
 sg13g2_nor2_1 _1004_ (.A(_0399_),
    .B(_0400_),
    .Y(_0401_));
 sg13g2_mux4_1 _1005_ (.S0(net192),
    .A0(\cpu0.ram[0][4] ),
    .A1(\cpu0.ram[1][4] ),
    .A2(\cpu0.ram[2][4] ),
    .A3(\cpu0.ram[3][4] ),
    .S1(net185),
    .X(_0402_));
 sg13g2_nor2_1 _1006_ (.A(net179),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_mux2_1 _1007_ (.A0(\cpu0.ram[4][4] ),
    .A1(\cpu0.ram[5][4] ),
    .S(net196),
    .X(_0404_));
 sg13g2_nor2b_1 _1008_ (.A(\cpu0.ram[7][4] ),
    .B_N(net195),
    .Y(_0405_));
 sg13g2_o21ai_1 _1009_ (.B1(net187),
    .Y(_0406_),
    .A1(net195),
    .A2(\cpu0.ram[6][4] ));
 sg13g2_o21ai_1 _1010_ (.B1(net178),
    .Y(_0407_),
    .A1(_0405_),
    .A2(_0406_));
 sg13g2_a21oi_1 _1011_ (.A1(net173),
    .A2(_0404_),
    .Y(_0408_),
    .B1(_0407_));
 sg13g2_nor3_1 _1012_ (.A(net176),
    .B(_0403_),
    .C(_0408_),
    .Y(_0409_));
 sg13g2_nor3_1 _1013_ (.A(_0253_),
    .B(_0401_),
    .C(_0409_),
    .Y(_0410_));
 sg13g2_a21o_2 _1014_ (.A2(_0392_),
    .A1(_0253_),
    .B1(_0410_),
    .X(_0411_));
 sg13g2_inv_1 _1015_ (.Y(_0412_),
    .A(_0411_));
 sg13g2_a21oi_2 _1016_ (.B1(_0384_),
    .Y(_0413_),
    .A2(_0411_),
    .A1(net170));
 sg13g2_mux2_1 _1017_ (.A0(net146),
    .A1(net311),
    .S(net159),
    .X(_0008_));
 sg13g2_nand2_1 _1018_ (.Y(_0414_),
    .A(\cpu0.b_reg[4] ),
    .B(_0279_));
 sg13g2_nand3_1 _1019_ (.B(_0352_),
    .C(_0414_),
    .A(_0351_),
    .Y(_0415_));
 sg13g2_xnor2_1 _1020_ (.Y(_0416_),
    .A(\cpu0.b_reg[5] ),
    .B(_0415_));
 sg13g2_or2_1 _1021_ (.X(_0417_),
    .B(_0416_),
    .A(\cpu0.a_reg[5] ));
 sg13g2_nand2_1 _1022_ (.Y(_0418_),
    .A(\cpu0.a_reg[5] ),
    .B(_0416_));
 sg13g2_nand2_1 _1023_ (.Y(_0419_),
    .A(_0417_),
    .B(_0418_));
 sg13g2_nand2_1 _1024_ (.Y(_0420_),
    .A(_0387_),
    .B(_0389_));
 sg13g2_xnor2_1 _1025_ (.Y(_0421_),
    .A(_0419_),
    .B(_0420_));
 sg13g2_a221oi_1 _1026_ (.B2(_0421_),
    .C1(_0254_),
    .B1(net167),
    .A1(\cpu0.a_reg[5] ),
    .Y(_0422_),
    .A2(_0240_));
 sg13g2_mux4_1 _1027_ (.S0(net191),
    .A0(\cpu0.ram[8][5] ),
    .A1(\cpu0.ram[9][5] ),
    .A2(\cpu0.ram[10][5] ),
    .A3(\cpu0.ram[11][5] ),
    .S1(net183),
    .X(_0423_));
 sg13g2_nor2_1 _1028_ (.A(net179),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_nor2b_1 _1029_ (.A(\cpu0.ram[13][5] ),
    .B_N(net195),
    .Y(_0425_));
 sg13g2_o21ai_1 _1030_ (.B1(net174),
    .Y(_0426_),
    .A1(net195),
    .A2(\cpu0.ram[12][5] ));
 sg13g2_o21ai_1 _1031_ (.B1(net188),
    .Y(_0427_),
    .A1(net201),
    .A2(\cpu0.ram[14][5] ));
 sg13g2_a21oi_1 _1032_ (.A1(net201),
    .A2(_0198_),
    .Y(_0428_),
    .B1(_0427_));
 sg13g2_o21ai_1 _1033_ (.B1(net182),
    .Y(_0429_),
    .A1(_0425_),
    .A2(_0426_));
 sg13g2_o21ai_1 _1034_ (.B1(net176),
    .Y(_0430_),
    .A1(_0428_),
    .A2(_0429_));
 sg13g2_mux4_1 _1035_ (.S0(net192),
    .A0(\cpu0.ram[0][5] ),
    .A1(\cpu0.ram[1][5] ),
    .A2(\cpu0.ram[2][5] ),
    .A3(\cpu0.ram[3][5] ),
    .S1(net185),
    .X(_0431_));
 sg13g2_mux2_1 _1036_ (.A0(\cpu0.ram[4][5] ),
    .A1(\cpu0.ram[5][5] ),
    .S(net194),
    .X(_0432_));
 sg13g2_nor2b_1 _1037_ (.A(\cpu0.ram[7][5] ),
    .B_N(net189),
    .Y(_0433_));
 sg13g2_o21ai_1 _1038_ (.B1(net187),
    .Y(_0434_),
    .A1(net189),
    .A2(\cpu0.ram[6][5] ));
 sg13g2_o21ai_1 _1039_ (.B1(net178),
    .Y(_0435_),
    .A1(_0433_),
    .A2(_0434_));
 sg13g2_a21oi_1 _1040_ (.A1(net173),
    .A2(_0432_),
    .Y(_0436_),
    .B1(_0435_));
 sg13g2_nor2_1 _1041_ (.A(net175),
    .B(_0436_),
    .Y(_0437_));
 sg13g2_o21ai_1 _1042_ (.B1(_0437_),
    .Y(_0438_),
    .A1(net180),
    .A2(_0431_));
 sg13g2_o21ai_1 _1043_ (.B1(_0438_),
    .Y(_0439_),
    .A1(_0424_),
    .A2(_0430_));
 sg13g2_nor2_1 _1044_ (.A(_0253_),
    .B(_0439_),
    .Y(_0440_));
 sg13g2_nor2_2 _1045_ (.A(_0422_),
    .B(_0440_),
    .Y(_0441_));
 sg13g2_mux2_1 _1046_ (.A0(net6),
    .A1(_0441_),
    .S(net170),
    .X(_0442_));
 sg13g2_mux2_1 _1047_ (.A0(net144),
    .A1(net366),
    .S(net159),
    .X(_0009_));
 sg13g2_a21o_1 _1048_ (.A2(_0279_),
    .A1(\cpu0.b_reg[5] ),
    .B1(_0415_),
    .X(_0443_));
 sg13g2_xnor2_1 _1049_ (.Y(_0444_),
    .A(\cpu0.b_reg[6] ),
    .B(_0443_));
 sg13g2_and2_1 _1050_ (.A(\cpu0.a_reg[6] ),
    .B(_0444_),
    .X(_0445_));
 sg13g2_xnor2_1 _1051_ (.Y(_0446_),
    .A(\cpu0.a_reg[6] ),
    .B(_0444_));
 sg13g2_nand2b_1 _1052_ (.Y(_0447_),
    .B(_0417_),
    .A_N(_0387_));
 sg13g2_and2_1 _1053_ (.A(_0418_),
    .B(_0447_),
    .X(_0448_));
 sg13g2_nand3b_1 _1054_ (.B(_0417_),
    .C(_0418_),
    .Y(_0449_),
    .A_N(_0388_));
 sg13g2_a21o_1 _1055_ (.A2(_0357_),
    .A1(_0354_),
    .B1(_0449_),
    .X(_0450_));
 sg13g2_and2_1 _1056_ (.A(_0448_),
    .B(_0450_),
    .X(_0451_));
 sg13g2_a21oi_1 _1057_ (.A1(_0448_),
    .A2(_0450_),
    .Y(_0452_),
    .B1(_0446_));
 sg13g2_xor2_1 _1058_ (.B(_0451_),
    .A(_0446_),
    .X(_0453_));
 sg13g2_a22oi_1 _1059_ (.Y(_0454_),
    .B1(_0246_),
    .B2(_0453_),
    .A2(_0240_),
    .A1(\cpu0.a_reg[6] ));
 sg13g2_mux4_1 _1060_ (.S0(net191),
    .A0(\cpu0.ram[8][6] ),
    .A1(\cpu0.ram[9][6] ),
    .A2(\cpu0.ram[10][6] ),
    .A3(\cpu0.ram[11][6] ),
    .S1(net183),
    .X(_0455_));
 sg13g2_nor2_1 _1061_ (.A(net177),
    .B(_0455_),
    .Y(_0456_));
 sg13g2_o21ai_1 _1062_ (.B1(net173),
    .Y(_0457_),
    .A1(net195),
    .A2(\cpu0.ram[12][6] ));
 sg13g2_a21oi_1 _1063_ (.A1(net195),
    .A2(_0199_),
    .Y(_0458_),
    .B1(_0457_));
 sg13g2_nor2b_1 _1064_ (.A(\cpu0.ram[15][6] ),
    .B_N(net200),
    .Y(_0459_));
 sg13g2_o21ai_1 _1065_ (.B1(_0001_),
    .Y(_0460_),
    .A1(net200),
    .A2(\cpu0.ram[14][6] ));
 sg13g2_o21ai_1 _1066_ (.B1(net180),
    .Y(_0461_),
    .A1(_0459_),
    .A2(_0460_));
 sg13g2_o21ai_1 _1067_ (.B1(net176),
    .Y(_0462_),
    .A1(_0458_),
    .A2(_0461_));
 sg13g2_mux4_1 _1068_ (.S0(net192),
    .A0(\cpu0.ram[0][6] ),
    .A1(\cpu0.ram[1][6] ),
    .A2(\cpu0.ram[2][6] ),
    .A3(\cpu0.ram[3][6] ),
    .S1(net185),
    .X(_0463_));
 sg13g2_mux2_1 _1069_ (.A0(\cpu0.ram[4][6] ),
    .A1(\cpu0.ram[5][6] ),
    .S(net196),
    .X(_0464_));
 sg13g2_nor2b_1 _1070_ (.A(\cpu0.ram[7][6] ),
    .B_N(net189),
    .Y(_0465_));
 sg13g2_o21ai_1 _1071_ (.B1(net183),
    .Y(_0466_),
    .A1(net189),
    .A2(\cpu0.ram[6][6] ));
 sg13g2_o21ai_1 _1072_ (.B1(net177),
    .Y(_0467_),
    .A1(_0465_),
    .A2(_0466_));
 sg13g2_a21oi_1 _1073_ (.A1(net173),
    .A2(_0464_),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_nor2_1 _1074_ (.A(net175),
    .B(_0468_),
    .Y(_0469_));
 sg13g2_o21ai_1 _1075_ (.B1(_0469_),
    .Y(_0470_),
    .A1(net179),
    .A2(_0463_));
 sg13g2_o21ai_1 _1076_ (.B1(_0470_),
    .Y(_0471_),
    .A1(_0456_),
    .A2(_0462_));
 sg13g2_nor2_1 _1077_ (.A(_0253_),
    .B(_0471_),
    .Y(_0472_));
 sg13g2_a21o_2 _1078_ (.A2(_0454_),
    .A1(_0253_),
    .B1(_0472_),
    .X(_0473_));
 sg13g2_nor2_1 _1079_ (.A(net7),
    .B(net170),
    .Y(_0474_));
 sg13g2_a21oi_2 _1080_ (.B1(_0474_),
    .Y(_0475_),
    .A2(_0473_),
    .A1(net168));
 sg13g2_mux2_1 _1081_ (.A0(net142),
    .A1(net317),
    .S(net159),
    .X(_0010_));
 sg13g2_a21oi_1 _1082_ (.A1(\cpu0.a_reg[7] ),
    .A2(_0240_),
    .Y(_0476_),
    .B1(_0254_));
 sg13g2_o21ai_1 _1083_ (.B1(_0279_),
    .Y(_0477_),
    .A1(\cpu0.b_reg[6] ),
    .A2(_0443_));
 sg13g2_xnor2_1 _1084_ (.Y(_0478_),
    .A(\cpu0.b_reg[7] ),
    .B(\cpu0.a_reg[7] ));
 sg13g2_xnor2_1 _1085_ (.Y(_0479_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_o21ai_1 _1086_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0445_),
    .A2(_0452_));
 sg13g2_or3_1 _1087_ (.A(_0445_),
    .B(_0452_),
    .C(_0479_),
    .X(_0481_));
 sg13g2_nand3_1 _1088_ (.B(_0480_),
    .C(_0481_),
    .A(net167),
    .Y(_0482_));
 sg13g2_mux4_1 _1089_ (.S0(net191),
    .A0(\cpu0.ram[8][7] ),
    .A1(\cpu0.ram[9][7] ),
    .A2(\cpu0.ram[10][7] ),
    .A3(\cpu0.ram[11][7] ),
    .S1(net183),
    .X(_0483_));
 sg13g2_nor2_1 _1090_ (.A(net177),
    .B(_0483_),
    .Y(_0484_));
 sg13g2_o21ai_1 _1091_ (.B1(net173),
    .Y(_0485_),
    .A1(net196),
    .A2(\cpu0.ram[12][7] ));
 sg13g2_a21oi_1 _1092_ (.A1(net196),
    .A2(_0200_),
    .Y(_0486_),
    .B1(_0485_));
 sg13g2_nor2b_1 _1093_ (.A(\cpu0.ram[15][7] ),
    .B_N(net200),
    .Y(_0487_));
 sg13g2_o21ai_1 _1094_ (.B1(net188),
    .Y(_0488_),
    .A1(net200),
    .A2(\cpu0.ram[14][7] ));
 sg13g2_o21ai_1 _1095_ (.B1(net182),
    .Y(_0489_),
    .A1(_0487_),
    .A2(_0488_));
 sg13g2_o21ai_1 _1096_ (.B1(net175),
    .Y(_0490_),
    .A1(_0486_),
    .A2(_0489_));
 sg13g2_nor2_1 _1097_ (.A(_0484_),
    .B(_0490_),
    .Y(_0491_));
 sg13g2_mux4_1 _1098_ (.S0(net192),
    .A0(\cpu0.ram[0][7] ),
    .A1(\cpu0.ram[1][7] ),
    .A2(\cpu0.ram[2][7] ),
    .A3(\cpu0.ram[3][7] ),
    .S1(net185),
    .X(_0492_));
 sg13g2_nor2_1 _1099_ (.A(net179),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_mux2_1 _1100_ (.A0(\cpu0.ram[4][7] ),
    .A1(\cpu0.ram[5][7] ),
    .S(net194),
    .X(_0494_));
 sg13g2_nor2b_1 _1101_ (.A(\cpu0.ram[7][7] ),
    .B_N(net189),
    .Y(_0495_));
 sg13g2_o21ai_1 _1102_ (.B1(net183),
    .Y(_0496_),
    .A1(net189),
    .A2(\cpu0.ram[6][7] ));
 sg13g2_o21ai_1 _1103_ (.B1(net178),
    .Y(_0497_),
    .A1(_0495_),
    .A2(_0496_));
 sg13g2_a21oi_1 _1104_ (.A1(net174),
    .A2(_0494_),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_nor3_1 _1105_ (.A(net175),
    .B(_0493_),
    .C(_0498_),
    .Y(_0499_));
 sg13g2_nor2_1 _1106_ (.A(_0491_),
    .B(_0499_),
    .Y(_0500_));
 sg13g2_a21o_1 _1107_ (.A2(_0500_),
    .A1(net161),
    .B1(_0219_),
    .X(_0501_));
 sg13g2_a21o_2 _1108_ (.A2(_0482_),
    .A1(_0476_),
    .B1(_0501_),
    .X(_0502_));
 sg13g2_nor2_1 _1109_ (.A(net8),
    .B(net170),
    .Y(_0503_));
 sg13g2_a21oi_2 _1110_ (.B1(_0503_),
    .Y(_0504_),
    .A2(_0502_),
    .A1(net168));
 sg13g2_mux2_1 _1111_ (.A0(net140),
    .A1(net353),
    .S(net159),
    .X(_0011_));
 sg13g2_o21ai_1 _1112_ (.B1(_0243_),
    .Y(_0505_),
    .A1(\cpu0.ir[7] ),
    .A2(_0202_));
 sg13g2_a21o_2 _1113_ (.A2(_0505_),
    .A1(_0222_),
    .B1(_0219_),
    .X(_0506_));
 sg13g2_o21ai_1 _1114_ (.B1(net205),
    .Y(_0507_),
    .A1(net467),
    .A2(net162));
 sg13g2_a21oi_1 _1115_ (.A1(_0276_),
    .A2(net162),
    .Y(_0012_),
    .B1(_0507_));
 sg13g2_o21ai_1 _1116_ (.B1(net204),
    .Y(_0508_),
    .A1(net469),
    .A2(net162));
 sg13g2_a21oi_1 _1117_ (.A1(_0310_),
    .A2(net162),
    .Y(_0013_),
    .B1(_0508_));
 sg13g2_o21ai_1 _1118_ (.B1(net205),
    .Y(_0509_),
    .A1(net464),
    .A2(net163));
 sg13g2_a21oi_1 _1119_ (.A1(_0346_),
    .A2(net163),
    .Y(_0014_),
    .B1(_0509_));
 sg13g2_o21ai_1 _1120_ (.B1(net204),
    .Y(_0510_),
    .A1(net463),
    .A2(net162));
 sg13g2_a21oi_1 _1121_ (.A1(_0381_),
    .A2(net162),
    .Y(_0015_),
    .B1(_0510_));
 sg13g2_nand2_1 _1122_ (.Y(_0511_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_nor2_2 _1123_ (.A(_0205_),
    .B(_0207_),
    .Y(_0512_));
 sg13g2_nand2_1 _1124_ (.Y(_0513_),
    .A(_0210_),
    .B(_0512_));
 sg13g2_or2_1 _1125_ (.X(_0514_),
    .B(_0513_),
    .A(_0511_));
 sg13g2_mux2_1 _1126_ (.A0(net150),
    .A1(net360),
    .S(_0514_),
    .X(_0016_));
 sg13g2_mux2_1 _1127_ (.A0(net154),
    .A1(net328),
    .S(_0514_),
    .X(_0017_));
 sg13g2_mux2_1 _1128_ (.A0(net152),
    .A1(net362),
    .S(_0514_),
    .X(_0018_));
 sg13g2_mux2_1 _1129_ (.A0(net148),
    .A1(net352),
    .S(_0514_),
    .X(_0019_));
 sg13g2_mux2_1 _1130_ (.A0(net146),
    .A1(net405),
    .S(_0514_),
    .X(_0020_));
 sg13g2_mux2_1 _1131_ (.A0(net144),
    .A1(net349),
    .S(_0514_),
    .X(_0021_));
 sg13g2_mux2_1 _1132_ (.A0(net142),
    .A1(net326),
    .S(_0514_),
    .X(_0022_));
 sg13g2_mux2_1 _1133_ (.A0(net140),
    .A1(net387),
    .S(_0514_),
    .X(_0023_));
 sg13g2_a21oi_1 _1134_ (.A1(net451),
    .A2(_0244_),
    .Y(_0024_),
    .B1(net203));
 sg13g2_nor2b_1 _1135_ (.A(_0245_),
    .B_N(_0220_),
    .Y(_0515_));
 sg13g2_or2_1 _1136_ (.X(_0025_),
    .B(_0515_),
    .A(_0222_));
 sg13g2_and3_1 _1137_ (.X(_0026_),
    .A(net207),
    .B(_0217_),
    .C(net451));
 sg13g2_or2_1 _1138_ (.X(_0516_),
    .B(_0513_),
    .A(_0215_));
 sg13g2_mux2_1 _1139_ (.A0(net150),
    .A1(net308),
    .S(_0516_),
    .X(_0027_));
 sg13g2_mux2_1 _1140_ (.A0(net154),
    .A1(net391),
    .S(_0516_),
    .X(_0028_));
 sg13g2_mux2_1 _1141_ (.A0(net152),
    .A1(net332),
    .S(_0516_),
    .X(_0029_));
 sg13g2_mux2_1 _1142_ (.A0(net148),
    .A1(net361),
    .S(_0516_),
    .X(_0030_));
 sg13g2_mux2_1 _1143_ (.A0(net146),
    .A1(net431),
    .S(_0516_),
    .X(_0031_));
 sg13g2_mux2_1 _1144_ (.A0(net144),
    .A1(net430),
    .S(_0516_),
    .X(_0032_));
 sg13g2_mux2_1 _1145_ (.A0(net142),
    .A1(net374),
    .S(_0516_),
    .X(_0033_));
 sg13g2_mux2_1 _1146_ (.A0(net140),
    .A1(net303),
    .S(_0516_),
    .X(_0034_));
 sg13g2_nand2_1 _1147_ (.Y(_0517_),
    .A(_0211_),
    .B(_0512_));
 sg13g2_or2_1 _1148_ (.X(_0518_),
    .B(_0517_),
    .A(_0511_));
 sg13g2_mux2_1 _1149_ (.A0(net150),
    .A1(net334),
    .S(_0518_),
    .X(_0035_));
 sg13g2_mux2_1 _1150_ (.A0(net154),
    .A1(net385),
    .S(_0518_),
    .X(_0036_));
 sg13g2_mux2_1 _1151_ (.A0(net152),
    .A1(net410),
    .S(_0518_),
    .X(_0037_));
 sg13g2_mux2_1 _1152_ (.A0(net148),
    .A1(net331),
    .S(_0518_),
    .X(_0038_));
 sg13g2_mux2_1 _1153_ (.A0(net146),
    .A1(net392),
    .S(_0518_),
    .X(_0039_));
 sg13g2_mux2_1 _1154_ (.A0(net144),
    .A1(net382),
    .S(_0518_),
    .X(_0040_));
 sg13g2_mux2_1 _1155_ (.A0(net142),
    .A1(net330),
    .S(_0518_),
    .X(_0041_));
 sg13g2_mux2_1 _1156_ (.A0(net140),
    .A1(net376),
    .S(_0518_),
    .X(_0042_));
 sg13g2_or2_1 _1157_ (.X(_0519_),
    .B(_0511_),
    .A(_0212_));
 sg13g2_mux2_1 _1158_ (.A0(net150),
    .A1(net316),
    .S(net158),
    .X(_0043_));
 sg13g2_mux2_1 _1159_ (.A0(net154),
    .A1(net304),
    .S(net158),
    .X(_0044_));
 sg13g2_mux2_1 _1160_ (.A0(net152),
    .A1(net324),
    .S(net158),
    .X(_0045_));
 sg13g2_nor2_1 _1161_ (.A(net148),
    .B(net158),
    .Y(_0520_));
 sg13g2_a21oi_1 _1162_ (.A1(_0196_),
    .A2(net158),
    .Y(_0046_),
    .B1(_0520_));
 sg13g2_mux2_1 _1163_ (.A0(net146),
    .A1(net307),
    .S(_0519_),
    .X(_0047_));
 sg13g2_mux2_1 _1164_ (.A0(net144),
    .A1(net344),
    .S(net158),
    .X(_0048_));
 sg13g2_mux2_1 _1165_ (.A0(net142),
    .A1(net367),
    .S(net158),
    .X(_0049_));
 sg13g2_mux2_1 _1166_ (.A0(net140),
    .A1(net389),
    .S(net158),
    .X(_0050_));
 sg13g2_nor2_2 _1167_ (.A(_0213_),
    .B(_0214_),
    .Y(_0521_));
 sg13g2_nand2_1 _1168_ (.Y(_0522_),
    .A(_0208_),
    .B(_0211_));
 sg13g2_inv_2 _1169_ (.Y(_0523_),
    .A(_0522_));
 sg13g2_nand2_2 _1170_ (.Y(_0524_),
    .A(_0521_),
    .B(_0523_));
 sg13g2_mux2_1 _1171_ (.A0(net149),
    .A1(net336),
    .S(net156),
    .X(_0051_));
 sg13g2_mux2_1 _1172_ (.A0(net153),
    .A1(net348),
    .S(net156),
    .X(_0052_));
 sg13g2_nor2_1 _1173_ (.A(net151),
    .B(net156),
    .Y(_0525_));
 sg13g2_a21oi_1 _1174_ (.A1(_0189_),
    .A2(_0524_),
    .Y(_0053_),
    .B1(_0525_));
 sg13g2_mux2_1 _1175_ (.A0(net147),
    .A1(net365),
    .S(net156),
    .X(_0054_));
 sg13g2_mux2_1 _1176_ (.A0(net145),
    .A1(net414),
    .S(net156),
    .X(_0055_));
 sg13g2_mux2_1 _1177_ (.A0(net143),
    .A1(net399),
    .S(net156),
    .X(_0056_));
 sg13g2_mux2_1 _1178_ (.A0(net141),
    .A1(net363),
    .S(net156),
    .X(_0057_));
 sg13g2_mux2_1 _1179_ (.A0(net139),
    .A1(net335),
    .S(net156),
    .X(_0058_));
 sg13g2_nand3_1 _1180_ (.B(_0512_),
    .C(_0521_),
    .A(_0211_),
    .Y(_0526_));
 sg13g2_mux2_1 _1181_ (.A0(net149),
    .A1(net386),
    .S(_0526_),
    .X(_0059_));
 sg13g2_mux2_1 _1182_ (.A0(net153),
    .A1(net397),
    .S(_0526_),
    .X(_0060_));
 sg13g2_mux2_1 _1183_ (.A0(net151),
    .A1(net394),
    .S(_0526_),
    .X(_0061_));
 sg13g2_mux2_1 _1184_ (.A0(net147),
    .A1(net370),
    .S(_0526_),
    .X(_0062_));
 sg13g2_mux2_1 _1185_ (.A0(net145),
    .A1(net347),
    .S(_0526_),
    .X(_0063_));
 sg13g2_mux2_1 _1186_ (.A0(net143),
    .A1(net395),
    .S(_0526_),
    .X(_0064_));
 sg13g2_mux2_1 _1187_ (.A0(net141),
    .A1(net408),
    .S(_0526_),
    .X(_0065_));
 sg13g2_mux2_1 _1188_ (.A0(net139),
    .A1(net419),
    .S(_0526_),
    .X(_0066_));
 sg13g2_nand3_1 _1189_ (.B(_0210_),
    .C(_0521_),
    .A(_0208_),
    .Y(_0527_));
 sg13g2_mux2_1 _1190_ (.A0(net149),
    .A1(net413),
    .S(_0527_),
    .X(_0067_));
 sg13g2_mux2_1 _1191_ (.A0(net154),
    .A1(net320),
    .S(_0527_),
    .X(_0068_));
 sg13g2_mux2_1 _1192_ (.A0(net152),
    .A1(net319),
    .S(_0527_),
    .X(_0069_));
 sg13g2_mux2_1 _1193_ (.A0(net147),
    .A1(net424),
    .S(_0527_),
    .X(_0070_));
 sg13g2_mux2_1 _1194_ (.A0(net145),
    .A1(net329),
    .S(_0527_),
    .X(_0071_));
 sg13g2_mux2_1 _1195_ (.A0(net143),
    .A1(net318),
    .S(_0527_),
    .X(_0072_));
 sg13g2_mux2_1 _1196_ (.A0(net141),
    .A1(net425),
    .S(_0527_),
    .X(_0073_));
 sg13g2_mux2_1 _1197_ (.A0(net139),
    .A1(net388),
    .S(_0527_),
    .X(_0074_));
 sg13g2_or2_1 _1198_ (.X(_0528_),
    .B(_0522_),
    .A(_0511_));
 sg13g2_mux2_1 _1199_ (.A0(net150),
    .A1(net402),
    .S(net157),
    .X(_0075_));
 sg13g2_nor2_1 _1200_ (.A(_0312_),
    .B(net157),
    .Y(_0529_));
 sg13g2_a21oi_1 _1201_ (.A1(_0187_),
    .A2(net157),
    .Y(_0076_),
    .B1(_0529_));
 sg13g2_mux2_1 _1202_ (.A0(_0348_),
    .A1(net436),
    .S(net157),
    .X(_0077_));
 sg13g2_mux2_1 _1203_ (.A0(_0383_),
    .A1(net381),
    .S(net157),
    .X(_0078_));
 sg13g2_mux2_1 _1204_ (.A0(net146),
    .A1(net339),
    .S(_0528_),
    .X(_0079_));
 sg13g2_mux2_1 _1205_ (.A0(net144),
    .A1(net369),
    .S(net157),
    .X(_0080_));
 sg13g2_mux2_1 _1206_ (.A0(net142),
    .A1(net393),
    .S(net157),
    .X(_0081_));
 sg13g2_mux2_1 _1207_ (.A0(net140),
    .A1(net314),
    .S(net157),
    .X(_0082_));
 sg13g2_nor2_2 _1208_ (.A(net202),
    .B(_0249_),
    .Y(_0530_));
 sg13g2_a22oi_1 _1209_ (.Y(_0531_),
    .B1(_0530_),
    .B2(net297),
    .A2(_0275_),
    .A1(_0250_));
 sg13g2_inv_1 _1210_ (.Y(_0083_),
    .A(net298));
 sg13g2_nand2_1 _1211_ (.Y(_0532_),
    .A(net276),
    .B(_0530_));
 sg13g2_o21ai_1 _1212_ (.B1(_0532_),
    .Y(_0084_),
    .A1(net171),
    .A2(_0310_));
 sg13g2_nand2_1 _1213_ (.Y(_0533_),
    .A(net274),
    .B(_0530_));
 sg13g2_o21ai_1 _1214_ (.B1(_0533_),
    .Y(_0085_),
    .A1(_0251_),
    .A2(_0346_));
 sg13g2_nand2_1 _1215_ (.Y(_0534_),
    .A(net278),
    .B(_0530_));
 sg13g2_o21ai_1 _1216_ (.B1(_0534_),
    .Y(_0086_),
    .A1(_0251_),
    .A2(_0381_));
 sg13g2_nand2_1 _1217_ (.Y(_0535_),
    .A(net440),
    .B(_0530_));
 sg13g2_o21ai_1 _1218_ (.B1(_0535_),
    .Y(_0087_),
    .A1(net171),
    .A2(_0411_));
 sg13g2_a22oi_1 _1219_ (.Y(_0536_),
    .B1(_0530_),
    .B2(net444),
    .A2(_0441_),
    .A1(_0250_));
 sg13g2_inv_1 _1220_ (.Y(_0088_),
    .A(net445));
 sg13g2_nand2_1 _1221_ (.Y(_0537_),
    .A(net446),
    .B(_0530_));
 sg13g2_o21ai_1 _1222_ (.B1(_0537_),
    .Y(_0089_),
    .A1(net171),
    .A2(_0473_));
 sg13g2_nand2_1 _1223_ (.Y(_0538_),
    .A(net448),
    .B(_0530_));
 sg13g2_o21ai_1 _1224_ (.B1(_0538_),
    .Y(_0090_),
    .A1(net171),
    .A2(_0502_));
 sg13g2_nor2_2 _1225_ (.A(net202),
    .B(_0238_),
    .Y(_0539_));
 sg13g2_a22oi_1 _1226_ (.Y(_0540_),
    .B1(_0539_),
    .B2(net434),
    .A2(_0275_),
    .A1(_0238_));
 sg13g2_inv_1 _1227_ (.Y(_0091_),
    .A(net435));
 sg13g2_nand2_1 _1228_ (.Y(_0541_),
    .A(net322),
    .B(_0539_));
 sg13g2_o21ai_1 _1229_ (.B1(_0541_),
    .Y(_0092_),
    .A1(_0239_),
    .A2(_0310_));
 sg13g2_nand2_1 _1230_ (.Y(_0542_),
    .A(net301),
    .B(_0539_));
 sg13g2_o21ai_1 _1231_ (.B1(_0542_),
    .Y(_0093_),
    .A1(_0239_),
    .A2(_0346_));
 sg13g2_nand2_1 _1232_ (.Y(_0543_),
    .A(net289),
    .B(_0539_));
 sg13g2_o21ai_1 _1233_ (.B1(_0543_),
    .Y(_0094_),
    .A1(_0239_),
    .A2(_0381_));
 sg13g2_nand2_1 _1234_ (.Y(_0544_),
    .A(net305),
    .B(_0539_));
 sg13g2_o21ai_1 _1235_ (.B1(_0544_),
    .Y(_0095_),
    .A1(_0239_),
    .A2(_0411_));
 sg13g2_a22oi_1 _1236_ (.Y(_0545_),
    .B1(_0539_),
    .B2(net420),
    .A2(_0441_),
    .A1(_0238_));
 sg13g2_inv_1 _1237_ (.Y(_0096_),
    .A(net421));
 sg13g2_nand2_1 _1238_ (.Y(_0546_),
    .A(net291),
    .B(_0539_));
 sg13g2_o21ai_1 _1239_ (.B1(_0546_),
    .Y(_0097_),
    .A1(_0239_),
    .A2(_0473_));
 sg13g2_nand2_1 _1240_ (.Y(_0547_),
    .A(net293),
    .B(_0539_));
 sg13g2_o21ai_1 _1241_ (.B1(_0547_),
    .Y(_0098_),
    .A1(_0239_),
    .A2(_0502_));
 sg13g2_nand2b_2 _1242_ (.Y(_0548_),
    .B(_0252_),
    .A_N(net167));
 sg13g2_inv_1 _1243_ (.Y(_0549_),
    .A(_0548_));
 sg13g2_and4_1 _1244_ (.A(_0180_),
    .B(\cpu0.ir[6] ),
    .C(_0222_),
    .D(_0241_),
    .X(_0550_));
 sg13g2_nor2_1 _1245_ (.A(_0548_),
    .B(_0550_),
    .Y(_0551_));
 sg13g2_or2_1 _1246_ (.X(_0552_),
    .B(_0550_),
    .A(_0548_));
 sg13g2_o21ai_1 _1247_ (.B1(net205),
    .Y(_0553_),
    .A1(net465),
    .A2(_0552_));
 sg13g2_a21oi_1 _1248_ (.A1(_0276_),
    .A2(_0552_),
    .Y(_0099_),
    .B1(_0553_));
 sg13g2_o21ai_1 _1249_ (.B1(net205),
    .Y(_0554_),
    .A1(net453),
    .A2(_0552_));
 sg13g2_a21oi_1 _1250_ (.A1(_0310_),
    .A2(_0552_),
    .Y(_0100_),
    .B1(_0554_));
 sg13g2_o21ai_1 _1251_ (.B1(net204),
    .Y(_0555_),
    .A1(net466),
    .A2(_0552_));
 sg13g2_a21oi_1 _1252_ (.A1(_0346_),
    .A2(_0552_),
    .Y(_0101_),
    .B1(_0555_));
 sg13g2_o21ai_1 _1253_ (.B1(net204),
    .Y(_0556_),
    .A1(net462),
    .A2(_0552_));
 sg13g2_a21oi_1 _1254_ (.A1(_0381_),
    .A2(_0552_),
    .Y(_0102_),
    .B1(_0556_));
 sg13g2_a22oi_1 _1255_ (.Y(_0557_),
    .B1(_0551_),
    .B2(net447),
    .A2(_0548_),
    .A1(_0412_));
 sg13g2_nor2_1 _1256_ (.A(net203),
    .B(_0557_),
    .Y(_0103_));
 sg13g2_a22oi_1 _1257_ (.Y(_0558_),
    .B1(_0551_),
    .B2(net441),
    .A2(_0548_),
    .A1(_0441_));
 sg13g2_nor2_1 _1258_ (.A(net203),
    .B(_0558_),
    .Y(_0104_));
 sg13g2_nand2_1 _1259_ (.Y(_0559_),
    .A(net471),
    .B(_0551_));
 sg13g2_o21ai_1 _1260_ (.B1(_0559_),
    .Y(_0560_),
    .A1(_0473_),
    .A2(_0549_));
 sg13g2_and2_1 _1261_ (.A(net204),
    .B(_0560_),
    .X(_0105_));
 sg13g2_nand2_1 _1262_ (.Y(_0561_),
    .A(net470),
    .B(_0551_));
 sg13g2_o21ai_1 _1263_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0502_),
    .A2(_0549_));
 sg13g2_and2_1 _1264_ (.A(net206),
    .B(_0562_),
    .X(_0106_));
 sg13g2_nand3_1 _1265_ (.B(net205),
    .C(net164),
    .A(net437),
    .Y(_0563_));
 sg13g2_o21ai_1 _1266_ (.B1(_0563_),
    .Y(_0107_),
    .A1(net164),
    .A2(_0276_));
 sg13g2_nand3_1 _1267_ (.B(net205),
    .C(net164),
    .A(net371),
    .Y(_0564_));
 sg13g2_o21ai_1 _1268_ (.B1(_0564_),
    .Y(_0108_),
    .A1(net164),
    .A2(_0310_));
 sg13g2_nand3_1 _1269_ (.B(net205),
    .C(net164),
    .A(net299),
    .Y(_0565_));
 sg13g2_o21ai_1 _1270_ (.B1(_0565_),
    .Y(_0109_),
    .A1(net164),
    .A2(_0346_));
 sg13g2_nand3_1 _1271_ (.B(net205),
    .C(net165),
    .A(net357),
    .Y(_0566_));
 sg13g2_o21ai_1 _1272_ (.B1(_0566_),
    .Y(_0110_),
    .A1(net164),
    .A2(_0381_));
 sg13g2_nand3_1 _1273_ (.B(net206),
    .C(net165),
    .A(net400),
    .Y(_0567_));
 sg13g2_o21ai_1 _1274_ (.B1(_0567_),
    .Y(_0111_),
    .A1(net164),
    .A2(_0411_));
 sg13g2_nor2_1 _1275_ (.A(net166),
    .B(_0441_),
    .Y(_0568_));
 sg13g2_o21ai_1 _1276_ (.B1(net204),
    .Y(_0569_),
    .A1(net455),
    .A2(_0247_));
 sg13g2_nor2_1 _1277_ (.A(_0568_),
    .B(net456),
    .Y(_0112_));
 sg13g2_nand3_1 _1278_ (.B(net206),
    .C(net165),
    .A(net309),
    .Y(_0570_));
 sg13g2_o21ai_1 _1279_ (.B1(_0570_),
    .Y(_0113_),
    .A1(net165),
    .A2(_0473_));
 sg13g2_nand2_1 _1280_ (.Y(_0571_),
    .A(net295),
    .B(net204));
 sg13g2_a22oi_1 _1281_ (.Y(_0114_),
    .B1(_0571_),
    .B2(net166),
    .A2(_0502_),
    .A1(_0247_));
 sg13g2_or2_1 _1282_ (.X(_0572_),
    .B(_0517_),
    .A(_0215_));
 sg13g2_mux2_1 _1283_ (.A0(_0278_),
    .A1(net364),
    .S(_0572_),
    .X(_0115_));
 sg13g2_mux2_1 _1284_ (.A0(net153),
    .A1(net383),
    .S(_0572_),
    .X(_0116_));
 sg13g2_mux2_1 _1285_ (.A0(net151),
    .A1(net337),
    .S(_0572_),
    .X(_0117_));
 sg13g2_mux2_1 _1286_ (.A0(net148),
    .A1(net368),
    .S(_0572_),
    .X(_0118_));
 sg13g2_mux2_1 _1287_ (.A0(net146),
    .A1(net345),
    .S(_0572_),
    .X(_0119_));
 sg13g2_mux2_1 _1288_ (.A0(net144),
    .A1(net384),
    .S(_0572_),
    .X(_0120_));
 sg13g2_mux2_1 _1289_ (.A0(net142),
    .A1(net417),
    .S(_0572_),
    .X(_0121_));
 sg13g2_mux2_1 _1290_ (.A0(net140),
    .A1(net380),
    .S(_0572_),
    .X(_0122_));
 sg13g2_nor2b_2 _1291_ (.A(_0213_),
    .B_N(_0214_),
    .Y(_0573_));
 sg13g2_nand3_1 _1292_ (.B(_0512_),
    .C(_0573_),
    .A(_0211_),
    .Y(_0574_));
 sg13g2_mux2_1 _1293_ (.A0(net149),
    .A1(net356),
    .S(_0574_),
    .X(_0123_));
 sg13g2_mux2_1 _1294_ (.A0(net153),
    .A1(net378),
    .S(_0574_),
    .X(_0124_));
 sg13g2_mux2_1 _1295_ (.A0(net151),
    .A1(net398),
    .S(_0574_),
    .X(_0125_));
 sg13g2_mux2_1 _1296_ (.A0(net147),
    .A1(net355),
    .S(_0574_),
    .X(_0126_));
 sg13g2_mux2_1 _1297_ (.A0(net145),
    .A1(net429),
    .S(_0574_),
    .X(_0127_));
 sg13g2_mux2_1 _1298_ (.A0(net143),
    .A1(net354),
    .S(_0574_),
    .X(_0128_));
 sg13g2_mux2_1 _1299_ (.A0(net141),
    .A1(net407),
    .S(_0574_),
    .X(_0129_));
 sg13g2_mux2_1 _1300_ (.A0(net139),
    .A1(net422),
    .S(_0574_),
    .X(_0130_));
 sg13g2_nand3_1 _1301_ (.B(_0512_),
    .C(_0573_),
    .A(_0210_),
    .Y(_0575_));
 sg13g2_mux2_1 _1302_ (.A0(net149),
    .A1(net406),
    .S(_0575_),
    .X(_0131_));
 sg13g2_mux2_1 _1303_ (.A0(net153),
    .A1(net340),
    .S(_0575_),
    .X(_0132_));
 sg13g2_mux2_1 _1304_ (.A0(net151),
    .A1(net338),
    .S(_0575_),
    .X(_0133_));
 sg13g2_mux2_1 _1305_ (.A0(net147),
    .A1(net415),
    .S(_0575_),
    .X(_0134_));
 sg13g2_mux2_1 _1306_ (.A0(net145),
    .A1(net404),
    .S(_0575_),
    .X(_0135_));
 sg13g2_mux2_1 _1307_ (.A0(net143),
    .A1(net411),
    .S(_0575_),
    .X(_0136_));
 sg13g2_mux2_1 _1308_ (.A0(net141),
    .A1(net390),
    .S(_0575_),
    .X(_0137_));
 sg13g2_mux2_1 _1309_ (.A0(net139),
    .A1(net310),
    .S(_0575_),
    .X(_0138_));
 sg13g2_nand3_1 _1310_ (.B(_0512_),
    .C(_0521_),
    .A(_0210_),
    .Y(_0576_));
 sg13g2_mux2_1 _1311_ (.A0(net150),
    .A1(net327),
    .S(_0576_),
    .X(_0139_));
 sg13g2_mux2_1 _1312_ (.A0(net154),
    .A1(net427),
    .S(_0576_),
    .X(_0140_));
 sg13g2_mux2_1 _1313_ (.A0(net152),
    .A1(net428),
    .S(_0576_),
    .X(_0141_));
 sg13g2_mux2_1 _1314_ (.A0(net147),
    .A1(net432),
    .S(_0576_),
    .X(_0142_));
 sg13g2_mux2_1 _1315_ (.A0(net145),
    .A1(net312),
    .S(_0576_),
    .X(_0143_));
 sg13g2_mux2_1 _1316_ (.A0(net143),
    .A1(net350),
    .S(_0576_),
    .X(_0144_));
 sg13g2_mux2_1 _1317_ (.A0(net141),
    .A1(net412),
    .S(_0576_),
    .X(_0145_));
 sg13g2_mux2_1 _1318_ (.A0(net139),
    .A1(net423),
    .S(_0576_),
    .X(_0146_));
 sg13g2_or2_1 _1319_ (.X(_0577_),
    .B(_0522_),
    .A(_0215_));
 sg13g2_mux2_1 _1320_ (.A0(net149),
    .A1(net433),
    .S(_0577_),
    .X(_0147_));
 sg13g2_mux2_1 _1321_ (.A0(net153),
    .A1(net426),
    .S(_0577_),
    .X(_0148_));
 sg13g2_mux2_1 _1322_ (.A0(net151),
    .A1(net439),
    .S(_0577_),
    .X(_0149_));
 sg13g2_mux2_1 _1323_ (.A0(net148),
    .A1(net342),
    .S(_0577_),
    .X(_0150_));
 sg13g2_mux2_1 _1324_ (.A0(net146),
    .A1(net375),
    .S(_0577_),
    .X(_0151_));
 sg13g2_mux2_1 _1325_ (.A0(net144),
    .A1(net325),
    .S(_0577_),
    .X(_0152_));
 sg13g2_mux2_1 _1326_ (.A0(net142),
    .A1(net351),
    .S(_0577_),
    .X(_0153_));
 sg13g2_mux2_1 _1327_ (.A0(net140),
    .A1(net373),
    .S(_0577_),
    .X(_0154_));
 sg13g2_nand2_2 _1328_ (.Y(_0578_),
    .A(_0523_),
    .B(_0573_));
 sg13g2_mux2_1 _1329_ (.A0(net149),
    .A1(net359),
    .S(net155),
    .X(_0155_));
 sg13g2_nor2_1 _1330_ (.A(net153),
    .B(net155),
    .Y(_0579_));
 sg13g2_a21oi_1 _1331_ (.A1(_0186_),
    .A2(net155),
    .Y(_0156_),
    .B1(_0579_));
 sg13g2_mux2_1 _1332_ (.A0(net151),
    .A1(net315),
    .S(net155),
    .X(_0157_));
 sg13g2_nor2_1 _1333_ (.A(net147),
    .B(_0578_),
    .Y(_0580_));
 sg13g2_a21oi_1 _1334_ (.A1(_0195_),
    .A2(_0578_),
    .Y(_0158_),
    .B1(_0580_));
 sg13g2_mux2_1 _1335_ (.A0(net145),
    .A1(net341),
    .S(net155),
    .X(_0159_));
 sg13g2_mux2_1 _1336_ (.A0(net143),
    .A1(net346),
    .S(net155),
    .X(_0160_));
 sg13g2_mux2_1 _1337_ (.A0(net141),
    .A1(net321),
    .S(net155),
    .X(_0161_));
 sg13g2_mux2_1 _1338_ (.A0(net139),
    .A1(net403),
    .S(net155),
    .X(_0162_));
 sg13g2_or2_1 _1339_ (.X(_0581_),
    .B(_0249_),
    .A(_0231_));
 sg13g2_inv_1 _1340_ (.Y(_0582_),
    .A(_0581_));
 sg13g2_nand2_1 _1341_ (.Y(_0583_),
    .A(net207),
    .B(_0581_));
 sg13g2_a21oi_1 _1342_ (.A1(net442),
    .A2(_0249_),
    .Y(_0584_),
    .B1(_0583_));
 sg13g2_o21ai_1 _1343_ (.B1(_0584_),
    .Y(_0585_),
    .A1(_0249_),
    .A2(_0275_));
 sg13g2_nand2_1 _1344_ (.Y(_0586_),
    .A(net442),
    .B(_0582_));
 sg13g2_a21oi_1 _1345_ (.A1(_0585_),
    .A2(_0586_),
    .Y(_0163_),
    .B1(net202));
 sg13g2_xnor2_1 _1346_ (.Y(_0587_),
    .A(net457),
    .B(net442));
 sg13g2_nand2_1 _1347_ (.Y(_0588_),
    .A(_0250_),
    .B(_0587_));
 sg13g2_a21oi_1 _1348_ (.A1(net171),
    .A2(_0310_),
    .Y(_0589_),
    .B1(_0583_));
 sg13g2_a22oi_1 _1349_ (.Y(_0590_),
    .B1(_0588_),
    .B2(_0589_),
    .A2(_0582_),
    .A1(net457));
 sg13g2_nor2_1 _1350_ (.A(net202),
    .B(net458),
    .Y(_0164_));
 sg13g2_a21oi_1 _1351_ (.A1(\cpu0.pc[1] ),
    .A2(\cpu0.pc[0] ),
    .Y(_0591_),
    .B1(net459));
 sg13g2_nand3_1 _1352_ (.B(\cpu0.pc[1] ),
    .C(\cpu0.pc[0] ),
    .A(net459),
    .Y(_0592_));
 sg13g2_nor2_1 _1353_ (.A(net171),
    .B(_0591_),
    .Y(_0593_));
 sg13g2_a21oi_1 _1354_ (.A1(_0592_),
    .A2(_0593_),
    .Y(_0594_),
    .B1(_0583_));
 sg13g2_o21ai_1 _1355_ (.B1(_0594_),
    .Y(_0595_),
    .A1(_0250_),
    .A2(_0346_));
 sg13g2_o21ai_1 _1356_ (.B1(_0595_),
    .Y(_0596_),
    .A1(net459),
    .A2(_0581_));
 sg13g2_nor2_1 _1357_ (.A(net202),
    .B(net460),
    .Y(_0165_));
 sg13g2_xnor2_1 _1358_ (.Y(_0597_),
    .A(net461),
    .B(_0592_));
 sg13g2_a21oi_1 _1359_ (.A1(_0250_),
    .A2(_0597_),
    .Y(_0598_),
    .B1(_0583_));
 sg13g2_o21ai_1 _1360_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0250_),
    .A2(_0381_));
 sg13g2_o21ai_1 _1361_ (.B1(_0599_),
    .Y(_0600_),
    .A1(net461),
    .A2(_0581_));
 sg13g2_nor2_1 _1362_ (.A(net202),
    .B(_0600_),
    .Y(_0166_));
 sg13g2_nand3_1 _1363_ (.B(_0210_),
    .C(_0573_),
    .A(_0208_),
    .Y(_0601_));
 sg13g2_mux2_1 _1364_ (.A0(net149),
    .A1(net396),
    .S(net160),
    .X(_0167_));
 sg13g2_mux2_1 _1365_ (.A0(net153),
    .A1(net313),
    .S(net160),
    .X(_0168_));
 sg13g2_mux2_1 _1366_ (.A0(net151),
    .A1(net343),
    .S(net160),
    .X(_0169_));
 sg13g2_nor2_1 _1367_ (.A(net147),
    .B(net160),
    .Y(_0602_));
 sg13g2_a21oi_1 _1368_ (.A1(_0194_),
    .A2(_0601_),
    .Y(_0170_),
    .B1(_0602_));
 sg13g2_mux2_1 _1369_ (.A0(net145),
    .A1(net418),
    .S(net160),
    .X(_0171_));
 sg13g2_mux2_1 _1370_ (.A0(net143),
    .A1(net379),
    .S(net160),
    .X(_0172_));
 sg13g2_mux2_1 _1371_ (.A0(net141),
    .A1(net401),
    .S(net160),
    .X(_0173_));
 sg13g2_mux2_1 _1372_ (.A0(net139),
    .A1(net409),
    .S(net160),
    .X(_0174_));
 sg13g2_a21oi_1 _1373_ (.A1(_0276_),
    .A2(net163),
    .Y(_0175_),
    .B1(_0507_));
 sg13g2_a21oi_1 _1374_ (.A1(_0310_),
    .A2(net162),
    .Y(_0176_),
    .B1(_0508_));
 sg13g2_a21oi_1 _1375_ (.A1(_0346_),
    .A2(net163),
    .Y(_0177_),
    .B1(_0509_));
 sg13g2_a21oi_1 _1376_ (.A1(_0381_),
    .A2(net162),
    .Y(_0178_),
    .B1(_0510_));
 sg13g2_dfrbpq_1 _1377_ (.RESET_B(net116),
    .D(_0004_),
    .Q(\cpu0.ram[5][0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net52),
    .D(_0005_),
    .Q(\cpu0.ram[5][1] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1379_ (.RESET_B(net51),
    .D(_0006_),
    .Q(\cpu0.ram[5][2] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net50),
    .D(_0007_),
    .Q(\cpu0.ram[5][3] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1381_ (.RESET_B(net49),
    .D(_0008_),
    .Q(\cpu0.ram[5][4] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1382_ (.RESET_B(net48),
    .D(_0009_),
    .Q(\cpu0.ram[5][5] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1383_ (.RESET_B(net47),
    .D(_0010_),
    .Q(\cpu0.ram[5][6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1384_ (.RESET_B(net46),
    .D(_0011_),
    .Q(\cpu0.ram[5][7] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1385_ (.RESET_B(net45),
    .D(_0012_),
    .Q(_0000_),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1386_ (.RESET_B(net44),
    .D(_0013_),
    .Q(_0001_),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net43),
    .D(_0014_),
    .Q(_0002_),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1388_ (.RESET_B(net42),
    .D(_0015_),
    .Q(_0003_),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1389_ (.RESET_B(net41),
    .D(_0016_),
    .Q(\cpu0.ram[12][0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1390_ (.RESET_B(net40),
    .D(_0017_),
    .Q(\cpu0.ram[12][1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net39),
    .D(_0018_),
    .Q(\cpu0.ram[12][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1392_ (.RESET_B(net38),
    .D(_0019_),
    .Q(\cpu0.ram[12][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1393_ (.RESET_B(net37),
    .D(_0020_),
    .Q(\cpu0.ram[12][4] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1394_ (.RESET_B(net36),
    .D(_0021_),
    .Q(\cpu0.ram[12][5] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net35),
    .D(_0022_),
    .Q(\cpu0.ram[12][6] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net34),
    .D(_0023_),
    .Q(\cpu0.ram[12][7] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1397_ (.RESET_B(net33),
    .D(net452),
    .Q(\cpu0.step[1] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1398_ (.RESET_B(net32),
    .D(_0025_),
    .Q(\cpu0.step[2] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1399_ (.RESET_B(net31),
    .D(_0026_),
    .Q(\cpu0.step[0] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1400_ (.RESET_B(net30),
    .D(_0027_),
    .Q(\cpu0.ram[4][0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1401_ (.RESET_B(net273),
    .D(_0028_),
    .Q(\cpu0.ram[4][1] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1402_ (.RESET_B(net272),
    .D(_0029_),
    .Q(\cpu0.ram[4][2] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1403_ (.RESET_B(net271),
    .D(_0030_),
    .Q(\cpu0.ram[4][3] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1404_ (.RESET_B(net270),
    .D(_0031_),
    .Q(\cpu0.ram[4][4] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1405_ (.RESET_B(net269),
    .D(_0032_),
    .Q(\cpu0.ram[4][5] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1406_ (.RESET_B(net268),
    .D(_0033_),
    .Q(\cpu0.ram[4][6] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1407_ (.RESET_B(net267),
    .D(_0034_),
    .Q(\cpu0.ram[4][7] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1408_ (.RESET_B(net266),
    .D(_0035_),
    .Q(\cpu0.ram[14][0] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1409_ (.RESET_B(net265),
    .D(_0036_),
    .Q(\cpu0.ram[14][1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1410_ (.RESET_B(net264),
    .D(_0037_),
    .Q(\cpu0.ram[14][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1411_ (.RESET_B(net263),
    .D(_0038_),
    .Q(\cpu0.ram[14][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1412_ (.RESET_B(net262),
    .D(_0039_),
    .Q(\cpu0.ram[14][4] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net261),
    .D(_0040_),
    .Q(\cpu0.ram[14][5] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net260),
    .D(_0041_),
    .Q(\cpu0.ram[14][6] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1415_ (.RESET_B(net259),
    .D(_0042_),
    .Q(\cpu0.ram[14][7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1416_ (.RESET_B(net258),
    .D(_0043_),
    .Q(\cpu0.ram[13][0] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1417_ (.RESET_B(net257),
    .D(_0044_),
    .Q(\cpu0.ram[13][1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1418_ (.RESET_B(net256),
    .D(_0045_),
    .Q(\cpu0.ram[13][2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1419_ (.RESET_B(net255),
    .D(_0046_),
    .Q(\cpu0.ram[13][3] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net254),
    .D(_0047_),
    .Q(\cpu0.ram[13][4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1421_ (.RESET_B(net253),
    .D(_0048_),
    .Q(\cpu0.ram[13][5] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net252),
    .D(_0049_),
    .Q(\cpu0.ram[13][6] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1423_ (.RESET_B(net251),
    .D(_0050_),
    .Q(\cpu0.ram[13][7] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net250),
    .D(_0051_),
    .Q(\cpu0.ram[3][0] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1425_ (.RESET_B(net249),
    .D(_0052_),
    .Q(\cpu0.ram[3][1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1426_ (.RESET_B(net248),
    .D(net287),
    .Q(\cpu0.ram[3][2] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1427_ (.RESET_B(net247),
    .D(_0054_),
    .Q(\cpu0.ram[3][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net246),
    .D(_0055_),
    .Q(\cpu0.ram[3][4] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net245),
    .D(_0056_),
    .Q(\cpu0.ram[3][5] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net244),
    .D(_0057_),
    .Q(\cpu0.ram[3][6] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1431_ (.RESET_B(net243),
    .D(_0058_),
    .Q(\cpu0.ram[3][7] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1432_ (.RESET_B(net242),
    .D(_0059_),
    .Q(\cpu0.ram[2][0] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1433_ (.RESET_B(net241),
    .D(_0060_),
    .Q(\cpu0.ram[2][1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1434_ (.RESET_B(net240),
    .D(_0061_),
    .Q(\cpu0.ram[2][2] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1435_ (.RESET_B(net239),
    .D(_0062_),
    .Q(\cpu0.ram[2][3] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1436_ (.RESET_B(net238),
    .D(_0063_),
    .Q(\cpu0.ram[2][4] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1437_ (.RESET_B(net237),
    .D(_0064_),
    .Q(\cpu0.ram[2][5] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1438_ (.RESET_B(net236),
    .D(_0065_),
    .Q(\cpu0.ram[2][6] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1439_ (.RESET_B(net235),
    .D(_0066_),
    .Q(\cpu0.ram[2][7] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1440_ (.RESET_B(net234),
    .D(_0067_),
    .Q(\cpu0.ram[1][0] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1441_ (.RESET_B(net233),
    .D(_0068_),
    .Q(\cpu0.ram[1][1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1442_ (.RESET_B(net232),
    .D(_0069_),
    .Q(\cpu0.ram[1][2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1443_ (.RESET_B(net231),
    .D(_0070_),
    .Q(\cpu0.ram[1][3] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net230),
    .D(_0071_),
    .Q(\cpu0.ram[1][4] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net229),
    .D(_0072_),
    .Q(\cpu0.ram[1][5] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net228),
    .D(_0073_),
    .Q(\cpu0.ram[1][6] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net227),
    .D(_0074_),
    .Q(\cpu0.ram[1][7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1448_ (.RESET_B(net226),
    .D(_0075_),
    .Q(\cpu0.ram[15][0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net225),
    .D(_0076_),
    .Q(\cpu0.ram[15][1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net224),
    .D(_0077_),
    .Q(\cpu0.ram[15][2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net223),
    .D(_0078_),
    .Q(\cpu0.ram[15][3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1452_ (.RESET_B(net222),
    .D(_0079_),
    .Q(\cpu0.ram[15][4] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net221),
    .D(_0080_),
    .Q(\cpu0.ram[15][5] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net220),
    .D(_0081_),
    .Q(\cpu0.ram[15][6] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net219),
    .D(_0082_),
    .Q(\cpu0.ram[15][7] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1456_ (.RESET_B(net218),
    .D(_0083_),
    .Q(\cpu0.ir[0] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net216),
    .D(net277),
    .Q(\cpu0.ir[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net214),
    .D(net275),
    .Q(\cpu0.ir[2] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net212),
    .D(net279),
    .Q(\cpu0.ir[3] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1460_ (.RESET_B(net210),
    .D(_0087_),
    .Q(\cpu0.ir[4] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1461_ (.RESET_B(net208),
    .D(_0088_),
    .Q(\cpu0.ir[5] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1462_ (.RESET_B(net137),
    .D(_0089_),
    .Q(\cpu0.ir[6] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1463_ (.RESET_B(net135),
    .D(net449),
    .Q(\cpu0.ir[7] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1464_ (.RESET_B(net133),
    .D(_0091_),
    .Q(uo_out[0]),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1465_ (.RESET_B(net131),
    .D(net323),
    .Q(uo_out[1]),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1466_ (.RESET_B(net129),
    .D(net302),
    .Q(uo_out[2]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1467_ (.RESET_B(net127),
    .D(net290),
    .Q(uo_out[3]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1468_ (.RESET_B(net125),
    .D(net306),
    .Q(uo_out[4]),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net123),
    .D(_0096_),
    .Q(uo_out[5]),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1470_ (.RESET_B(net121),
    .D(net292),
    .Q(uo_out[6]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1471_ (.RESET_B(net119),
    .D(net294),
    .Q(uo_out[7]),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1472_ (.RESET_B(net117),
    .D(_0099_),
    .Q(\cpu0.a_reg[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1473_ (.RESET_B(net115),
    .D(net454),
    .Q(\cpu0.a_reg[1] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1474_ (.RESET_B(net113),
    .D(_0101_),
    .Q(\cpu0.a_reg[2] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1475_ (.RESET_B(net111),
    .D(_0102_),
    .Q(\cpu0.a_reg[3] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1476_ (.RESET_B(net109),
    .D(_0103_),
    .Q(\cpu0.a_reg[4] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1477_ (.RESET_B(net107),
    .D(_0104_),
    .Q(\cpu0.a_reg[5] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1478_ (.RESET_B(net105),
    .D(_0105_),
    .Q(\cpu0.a_reg[6] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1479_ (.RESET_B(net103),
    .D(_0106_),
    .Q(\cpu0.a_reg[7] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1480_ (.RESET_B(net101),
    .D(net438),
    .Q(\cpu0.b_reg[0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1481_ (.RESET_B(net99),
    .D(net372),
    .Q(\cpu0.b_reg[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net97),
    .D(net300),
    .Q(\cpu0.b_reg[2] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1483_ (.RESET_B(net95),
    .D(net358),
    .Q(\cpu0.b_reg[3] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net93),
    .D(_0111_),
    .Q(\cpu0.b_reg[4] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1485_ (.RESET_B(net91),
    .D(_0112_),
    .Q(\cpu0.b_reg[5] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1486_ (.RESET_B(net89),
    .D(_0113_),
    .Q(\cpu0.b_reg[6] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1487_ (.RESET_B(net87),
    .D(net296),
    .Q(\cpu0.b_reg[7] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1488_ (.RESET_B(net85),
    .D(_0115_),
    .Q(\cpu0.ram[6][0] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1489_ (.RESET_B(net84),
    .D(_0116_),
    .Q(\cpu0.ram[6][1] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net83),
    .D(_0117_),
    .Q(\cpu0.ram[6][2] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1491_ (.RESET_B(net82),
    .D(_0118_),
    .Q(\cpu0.ram[6][3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net81),
    .D(_0119_),
    .Q(\cpu0.ram[6][4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1493_ (.RESET_B(net80),
    .D(_0120_),
    .Q(\cpu0.ram[6][5] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net79),
    .D(_0121_),
    .Q(\cpu0.ram[6][6] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1495_ (.RESET_B(net78),
    .D(_0122_),
    .Q(\cpu0.ram[6][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1496_ (.RESET_B(net77),
    .D(_0123_),
    .Q(\cpu0.ram[10][0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1497_ (.RESET_B(net76),
    .D(_0124_),
    .Q(\cpu0.ram[10][1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net75),
    .D(_0125_),
    .Q(\cpu0.ram[10][2] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1499_ (.RESET_B(net74),
    .D(_0126_),
    .Q(\cpu0.ram[10][3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1500_ (.RESET_B(net73),
    .D(_0127_),
    .Q(\cpu0.ram[10][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1501_ (.RESET_B(net72),
    .D(_0128_),
    .Q(\cpu0.ram[10][5] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net71),
    .D(_0129_),
    .Q(\cpu0.ram[10][6] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1503_ (.RESET_B(net70),
    .D(_0130_),
    .Q(\cpu0.ram[10][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1504_ (.RESET_B(net69),
    .D(_0131_),
    .Q(\cpu0.ram[8][0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1505_ (.RESET_B(net68),
    .D(_0132_),
    .Q(\cpu0.ram[8][1] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net67),
    .D(_0133_),
    .Q(\cpu0.ram[8][2] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1507_ (.RESET_B(net66),
    .D(_0134_),
    .Q(\cpu0.ram[8][3] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net65),
    .D(_0135_),
    .Q(\cpu0.ram[8][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1509_ (.RESET_B(net64),
    .D(_0136_),
    .Q(\cpu0.ram[8][5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1510_ (.RESET_B(net63),
    .D(_0137_),
    .Q(\cpu0.ram[8][6] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1511_ (.RESET_B(net62),
    .D(_0138_),
    .Q(\cpu0.ram[8][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net61),
    .D(_0139_),
    .Q(\cpu0.ram[0][0] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1513_ (.RESET_B(net60),
    .D(_0140_),
    .Q(\cpu0.ram[0][1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1514_ (.RESET_B(net59),
    .D(_0141_),
    .Q(\cpu0.ram[0][2] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1515_ (.RESET_B(net58),
    .D(_0142_),
    .Q(\cpu0.ram[0][3] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1516_ (.RESET_B(net57),
    .D(_0143_),
    .Q(\cpu0.ram[0][4] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1517_ (.RESET_B(net56),
    .D(_0144_),
    .Q(\cpu0.ram[0][5] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1518_ (.RESET_B(net55),
    .D(_0145_),
    .Q(\cpu0.ram[0][6] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1519_ (.RESET_B(net54),
    .D(_0146_),
    .Q(\cpu0.ram[0][7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1520_ (.RESET_B(net53),
    .D(_0147_),
    .Q(\cpu0.ram[7][0] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1521_ (.RESET_B(net217),
    .D(_0148_),
    .Q(\cpu0.ram[7][1] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1522_ (.RESET_B(net215),
    .D(_0149_),
    .Q(\cpu0.ram[7][2] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1523_ (.RESET_B(net213),
    .D(_0150_),
    .Q(\cpu0.ram[7][3] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1524_ (.RESET_B(net211),
    .D(_0151_),
    .Q(\cpu0.ram[7][4] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1525_ (.RESET_B(net209),
    .D(_0152_),
    .Q(\cpu0.ram[7][5] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1526_ (.RESET_B(net138),
    .D(_0153_),
    .Q(\cpu0.ram[7][6] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1527_ (.RESET_B(net136),
    .D(_0154_),
    .Q(\cpu0.ram[7][7] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1528_ (.RESET_B(net134),
    .D(_0155_),
    .Q(\cpu0.ram[11][0] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1529_ (.RESET_B(net132),
    .D(_0156_),
    .Q(\cpu0.ram[11][1] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1530_ (.RESET_B(net130),
    .D(_0157_),
    .Q(\cpu0.ram[11][2] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1531_ (.RESET_B(net128),
    .D(_0158_),
    .Q(\cpu0.ram[11][3] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1532_ (.RESET_B(net126),
    .D(_0159_),
    .Q(\cpu0.ram[11][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1533_ (.RESET_B(net124),
    .D(_0160_),
    .Q(\cpu0.ram[11][5] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1534_ (.RESET_B(net122),
    .D(_0161_),
    .Q(\cpu0.ram[11][6] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1535_ (.RESET_B(net120),
    .D(_0162_),
    .Q(\cpu0.ram[11][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_2 _1536_ (.RESET_B(net118),
    .D(net443),
    .Q(\cpu0.pc[0] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1537_ (.RESET_B(net114),
    .D(_0164_),
    .Q(\cpu0.pc[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1538_ (.RESET_B(net110),
    .D(_0165_),
    .Q(\cpu0.pc[2] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1539_ (.RESET_B(net106),
    .D(_0166_),
    .Q(\cpu0.pc[3] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1540_ (.RESET_B(net102),
    .D(_0167_),
    .Q(\cpu0.ram[9][0] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1541_ (.RESET_B(net100),
    .D(_0168_),
    .Q(\cpu0.ram[9][1] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1542_ (.RESET_B(net98),
    .D(_0169_),
    .Q(\cpu0.ram[9][2] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1543_ (.RESET_B(net96),
    .D(net282),
    .Q(\cpu0.ram[9][3] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1544_ (.RESET_B(net94),
    .D(_0171_),
    .Q(\cpu0.ram[9][4] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1545_ (.RESET_B(net92),
    .D(_0172_),
    .Q(\cpu0.ram[9][5] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1546_ (.RESET_B(net90),
    .D(_0173_),
    .Q(\cpu0.ram[9][6] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1547_ (.RESET_B(net88),
    .D(_0174_),
    .Q(\cpu0.ram[9][7] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1548_ (.RESET_B(net86),
    .D(_0175_),
    .Q(\cpu0.mar[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1549_ (.RESET_B(net112),
    .D(_0176_),
    .Q(\cpu0.mar[1] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1550_ (.RESET_B(net104),
    .D(_0177_),
    .Q(\cpu0.mar[2] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1551_ (.RESET_B(net108),
    .D(_0178_),
    .Q(\cpu0.mar[3] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_tiehi _1399__31 (.L_HI(net31));
 sg13g2_tiehi _1398__32 (.L_HI(net32));
 sg13g2_tiehi _1397__33 (.L_HI(net33));
 sg13g2_tiehi _1396__34 (.L_HI(net34));
 sg13g2_tiehi _1395__35 (.L_HI(net35));
 sg13g2_tiehi _1394__36 (.L_HI(net36));
 sg13g2_tiehi _1393__37 (.L_HI(net37));
 sg13g2_tiehi _1392__38 (.L_HI(net38));
 sg13g2_tiehi _1391__39 (.L_HI(net39));
 sg13g2_tiehi _1390__40 (.L_HI(net40));
 sg13g2_tiehi _1389__41 (.L_HI(net41));
 sg13g2_tiehi _1388__42 (.L_HI(net42));
 sg13g2_tiehi _1387__43 (.L_HI(net43));
 sg13g2_tiehi _1386__44 (.L_HI(net44));
 sg13g2_tiehi _1385__45 (.L_HI(net45));
 sg13g2_tiehi _1384__46 (.L_HI(net46));
 sg13g2_tiehi _1383__47 (.L_HI(net47));
 sg13g2_tiehi _1382__48 (.L_HI(net48));
 sg13g2_tiehi _1381__49 (.L_HI(net49));
 sg13g2_tiehi _1380__50 (.L_HI(net50));
 sg13g2_tiehi _1379__51 (.L_HI(net51));
 sg13g2_tiehi _1378__52 (.L_HI(net52));
 sg13g2_tiehi _1520__53 (.L_HI(net53));
 sg13g2_tiehi _1519__54 (.L_HI(net54));
 sg13g2_tiehi _1518__55 (.L_HI(net55));
 sg13g2_tiehi _1517__56 (.L_HI(net56));
 sg13g2_tiehi _1516__57 (.L_HI(net57));
 sg13g2_tiehi _1515__58 (.L_HI(net58));
 sg13g2_tiehi _1514__59 (.L_HI(net59));
 sg13g2_tiehi _1513__60 (.L_HI(net60));
 sg13g2_tiehi _1512__61 (.L_HI(net61));
 sg13g2_tiehi _1511__62 (.L_HI(net62));
 sg13g2_tiehi _1510__63 (.L_HI(net63));
 sg13g2_tiehi _1509__64 (.L_HI(net64));
 sg13g2_tiehi _1508__65 (.L_HI(net65));
 sg13g2_tiehi _1507__66 (.L_HI(net66));
 sg13g2_tiehi _1506__67 (.L_HI(net67));
 sg13g2_tiehi _1505__68 (.L_HI(net68));
 sg13g2_tiehi _1504__69 (.L_HI(net69));
 sg13g2_tiehi _1503__70 (.L_HI(net70));
 sg13g2_tiehi _1502__71 (.L_HI(net71));
 sg13g2_tiehi _1501__72 (.L_HI(net72));
 sg13g2_tiehi _1500__73 (.L_HI(net73));
 sg13g2_tiehi _1499__74 (.L_HI(net74));
 sg13g2_tiehi _1498__75 (.L_HI(net75));
 sg13g2_tiehi _1497__76 (.L_HI(net76));
 sg13g2_tiehi _1496__77 (.L_HI(net77));
 sg13g2_tiehi _1495__78 (.L_HI(net78));
 sg13g2_tiehi _1494__79 (.L_HI(net79));
 sg13g2_tiehi _1493__80 (.L_HI(net80));
 sg13g2_tiehi _1492__81 (.L_HI(net81));
 sg13g2_tiehi _1491__82 (.L_HI(net82));
 sg13g2_tiehi _1490__83 (.L_HI(net83));
 sg13g2_tiehi _1489__84 (.L_HI(net84));
 sg13g2_tiehi _1488__85 (.L_HI(net85));
 sg13g2_tiehi _1548__86 (.L_HI(net86));
 sg13g2_tiehi _1487__87 (.L_HI(net87));
 sg13g2_tiehi _1547__88 (.L_HI(net88));
 sg13g2_tiehi _1486__89 (.L_HI(net89));
 sg13g2_tiehi _1546__90 (.L_HI(net90));
 sg13g2_tiehi _1485__91 (.L_HI(net91));
 sg13g2_tiehi _1545__92 (.L_HI(net92));
 sg13g2_tiehi _1484__93 (.L_HI(net93));
 sg13g2_tiehi _1544__94 (.L_HI(net94));
 sg13g2_tiehi _1483__95 (.L_HI(net95));
 sg13g2_tiehi _1543__96 (.L_HI(net96));
 sg13g2_tiehi _1482__97 (.L_HI(net97));
 sg13g2_tiehi _1542__98 (.L_HI(net98));
 sg13g2_tiehi _1481__99 (.L_HI(net99));
 sg13g2_tiehi _1541__100 (.L_HI(net100));
 sg13g2_tiehi _1480__101 (.L_HI(net101));
 sg13g2_tiehi _1540__102 (.L_HI(net102));
 sg13g2_tiehi _1479__103 (.L_HI(net103));
 sg13g2_tiehi _1550__104 (.L_HI(net104));
 sg13g2_tiehi _1478__105 (.L_HI(net105));
 sg13g2_tiehi _1539__106 (.L_HI(net106));
 sg13g2_tiehi _1477__107 (.L_HI(net107));
 sg13g2_tiehi _1551__108 (.L_HI(net108));
 sg13g2_tiehi _1476__109 (.L_HI(net109));
 sg13g2_tiehi _1538__110 (.L_HI(net110));
 sg13g2_tiehi _1475__111 (.L_HI(net111));
 sg13g2_tiehi _1549__112 (.L_HI(net112));
 sg13g2_tiehi _1474__113 (.L_HI(net113));
 sg13g2_tiehi _1537__114 (.L_HI(net114));
 sg13g2_tiehi _1473__115 (.L_HI(net115));
 sg13g2_tiehi _1377__116 (.L_HI(net116));
 sg13g2_tiehi _1472__117 (.L_HI(net117));
 sg13g2_tiehi _1536__118 (.L_HI(net118));
 sg13g2_tiehi _1471__119 (.L_HI(net119));
 sg13g2_tiehi _1535__120 (.L_HI(net120));
 sg13g2_tiehi _1470__121 (.L_HI(net121));
 sg13g2_tiehi _1534__122 (.L_HI(net122));
 sg13g2_tiehi _1469__123 (.L_HI(net123));
 sg13g2_tiehi _1533__124 (.L_HI(net124));
 sg13g2_tiehi _1468__125 (.L_HI(net125));
 sg13g2_tiehi _1532__126 (.L_HI(net126));
 sg13g2_tiehi _1467__127 (.L_HI(net127));
 sg13g2_tiehi _1531__128 (.L_HI(net128));
 sg13g2_tiehi _1466__129 (.L_HI(net129));
 sg13g2_tiehi _1530__130 (.L_HI(net130));
 sg13g2_tiehi _1465__131 (.L_HI(net131));
 sg13g2_tiehi _1529__132 (.L_HI(net132));
 sg13g2_tiehi _1464__133 (.L_HI(net133));
 sg13g2_tiehi _1528__134 (.L_HI(net134));
 sg13g2_tiehi _1463__135 (.L_HI(net135));
 sg13g2_tiehi _1527__136 (.L_HI(net136));
 sg13g2_tiehi _1462__137 (.L_HI(net137));
 sg13g2_tiehi _1526__138 (.L_HI(net138));
 sg13g2_tiehi _1461__139 (.L_HI(net208));
 sg13g2_tiehi _1525__140 (.L_HI(net209));
 sg13g2_tiehi _1460__141 (.L_HI(net210));
 sg13g2_tiehi _1524__142 (.L_HI(net211));
 sg13g2_tiehi _1459__143 (.L_HI(net212));
 sg13g2_tiehi _1523__144 (.L_HI(net213));
 sg13g2_tiehi _1458__145 (.L_HI(net214));
 sg13g2_tiehi _1522__146 (.L_HI(net215));
 sg13g2_tiehi _1457__147 (.L_HI(net216));
 sg13g2_tiehi _1521__148 (.L_HI(net217));
 sg13g2_tiehi _1456__149 (.L_HI(net218));
 sg13g2_tiehi _1455__150 (.L_HI(net219));
 sg13g2_tiehi _1454__151 (.L_HI(net220));
 sg13g2_tiehi _1453__152 (.L_HI(net221));
 sg13g2_tiehi _1452__153 (.L_HI(net222));
 sg13g2_tiehi _1451__154 (.L_HI(net223));
 sg13g2_tiehi _1450__155 (.L_HI(net224));
 sg13g2_tiehi _1449__156 (.L_HI(net225));
 sg13g2_tiehi _1448__157 (.L_HI(net226));
 sg13g2_tiehi _1447__158 (.L_HI(net227));
 sg13g2_tiehi _1446__159 (.L_HI(net228));
 sg13g2_tiehi _1445__160 (.L_HI(net229));
 sg13g2_tiehi _1444__161 (.L_HI(net230));
 sg13g2_tiehi _1443__162 (.L_HI(net231));
 sg13g2_tiehi _1442__163 (.L_HI(net232));
 sg13g2_tiehi _1441__164 (.L_HI(net233));
 sg13g2_tiehi _1440__165 (.L_HI(net234));
 sg13g2_tiehi _1439__166 (.L_HI(net235));
 sg13g2_tiehi _1438__167 (.L_HI(net236));
 sg13g2_tiehi _1437__168 (.L_HI(net237));
 sg13g2_tiehi _1436__169 (.L_HI(net238));
 sg13g2_tiehi _1435__170 (.L_HI(net239));
 sg13g2_tiehi _1434__171 (.L_HI(net240));
 sg13g2_tiehi _1433__172 (.L_HI(net241));
 sg13g2_tiehi _1432__173 (.L_HI(net242));
 sg13g2_tiehi _1431__174 (.L_HI(net243));
 sg13g2_tiehi _1430__175 (.L_HI(net244));
 sg13g2_tiehi _1429__176 (.L_HI(net245));
 sg13g2_tiehi _1428__177 (.L_HI(net246));
 sg13g2_tiehi _1427__178 (.L_HI(net247));
 sg13g2_tiehi _1426__179 (.L_HI(net248));
 sg13g2_tiehi _1425__180 (.L_HI(net249));
 sg13g2_tiehi _1424__181 (.L_HI(net250));
 sg13g2_tiehi _1423__182 (.L_HI(net251));
 sg13g2_tiehi _1422__183 (.L_HI(net252));
 sg13g2_tiehi _1421__184 (.L_HI(net253));
 sg13g2_tiehi _1420__185 (.L_HI(net254));
 sg13g2_tiehi _1419__186 (.L_HI(net255));
 sg13g2_tiehi _1418__187 (.L_HI(net256));
 sg13g2_tiehi _1417__188 (.L_HI(net257));
 sg13g2_tiehi _1416__189 (.L_HI(net258));
 sg13g2_tiehi _1415__190 (.L_HI(net259));
 sg13g2_tiehi _1414__191 (.L_HI(net260));
 sg13g2_tiehi _1413__192 (.L_HI(net261));
 sg13g2_tiehi _1412__193 (.L_HI(net262));
 sg13g2_tiehi _1411__194 (.L_HI(net263));
 sg13g2_tiehi _1410__195 (.L_HI(net264));
 sg13g2_tiehi _1409__196 (.L_HI(net265));
 sg13g2_tiehi _1408__197 (.L_HI(net266));
 sg13g2_tiehi _1407__198 (.L_HI(net267));
 sg13g2_tiehi _1406__199 (.L_HI(net268));
 sg13g2_tiehi _1405__200 (.L_HI(net269));
 sg13g2_tiehi _1404__201 (.L_HI(net270));
 sg13g2_tiehi _1403__202 (.L_HI(net271));
 sg13g2_tiehi _1402__203 (.L_HI(net272));
 sg13g2_tiehi _1401__204 (.L_HI(net273));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_dranoel06_SAP1_15 (.L_LO(net15));
 sg13g2_tielo tt_um_dranoel06_SAP1_16 (.L_LO(net16));
 sg13g2_tielo tt_um_dranoel06_SAP1_17 (.L_LO(net17));
 sg13g2_tielo tt_um_dranoel06_SAP1_18 (.L_LO(net18));
 sg13g2_tielo tt_um_dranoel06_SAP1_19 (.L_LO(net19));
 sg13g2_tielo tt_um_dranoel06_SAP1_20 (.L_LO(net20));
 sg13g2_tielo tt_um_dranoel06_SAP1_21 (.L_LO(net21));
 sg13g2_tielo tt_um_dranoel06_SAP1_22 (.L_LO(net22));
 sg13g2_tielo tt_um_dranoel06_SAP1_23 (.L_LO(net23));
 sg13g2_tielo tt_um_dranoel06_SAP1_24 (.L_LO(net24));
 sg13g2_tielo tt_um_dranoel06_SAP1_25 (.L_LO(net25));
 sg13g2_tielo tt_um_dranoel06_SAP1_26 (.L_LO(net26));
 sg13g2_tielo tt_um_dranoel06_SAP1_27 (.L_LO(net27));
 sg13g2_tielo tt_um_dranoel06_SAP1_28 (.L_LO(net28));
 sg13g2_tielo tt_um_dranoel06_SAP1_29 (.L_LO(net29));
 sg13g2_tiehi _1400__30 (.L_HI(net30));
 sg13g2_buf_8 fanout139 (.A(_0504_),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(_0504_),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(_0475_),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(_0475_),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(_0442_),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0442_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0413_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(_0413_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(_0383_),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(_0278_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(_0348_),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(_0312_),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(_0578_),
    .X(net155));
 sg13g2_buf_8 fanout156 (.A(_0524_),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(_0528_),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(_0519_),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(_0216_),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(_0601_),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(_0254_),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(_0506_),
    .X(net162));
 sg13g2_buf_1 fanout163 (.A(_0506_),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(net165),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_1 fanout166 (.A(_0248_),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(_0246_),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net170),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(_0206_),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(_0251_),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(_0219_),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(_0183_),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(_0003_),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(net181),
    .X(net177));
 sg13g2_buf_1 fanout178 (.A(net181),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(net181),
    .X(net179));
 sg13g2_buf_1 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_8 fanout182 (.A(_0002_),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(net186),
    .X(net183));
 sg13g2_buf_1 fanout184 (.A(net186),
    .X(net184));
 sg13g2_buf_8 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_0001_),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(_0001_),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(net191),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_8 fanout191 (.A(net193),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_8 fanout193 (.A(_0000_),
    .X(net193));
 sg13g2_buf_8 fanout194 (.A(net196),
    .X(net194));
 sg13g2_buf_8 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(net199),
    .X(net196));
 sg13g2_buf_8 fanout197 (.A(net198),
    .X(net197));
 sg13g2_buf_8 fanout198 (.A(net199),
    .X(net198));
 sg13g2_buf_8 fanout199 (.A(net201),
    .X(net199));
 sg13g2_buf_8 fanout200 (.A(net201),
    .X(net200));
 sg13g2_buf_8 fanout201 (.A(_0000_),
    .X(net201));
 sg13g2_buf_8 fanout202 (.A(net203),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_0182_),
    .X(net203));
 sg13g2_buf_8 fanout204 (.A(net206),
    .X(net204));
 sg13g2_buf_8 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_8 fanout206 (.A(rst_n),
    .X(net206));
 sg13g2_buf_8 fanout207 (.A(rst_n),
    .X(net207));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_dranoel06_SAP1_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkload15 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cpu0.ir[2] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0085_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold3 (.A(\cpu0.ir[1] ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0084_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold5 (.A(\cpu0.ir[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0086_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold7 (.A(\cpu0.ram[11][3] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold8 (.A(\cpu0.ram[9][3] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0170_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cpu0.ram[11][1] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold11 (.A(\cpu0.ram[13][3] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold12 (.A(\cpu0.ram[5][2] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold13 (.A(\cpu0.ram[3][2] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0053_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cpu0.ram[15][1] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold16 (.A(uo_out[3]),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0094_),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold18 (.A(uo_out[6]),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0097_),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold20 (.A(uo_out[7]),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0098_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold22 (.A(\cpu0.b_reg[7] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0114_),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cpu0.ir[0] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0531_),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold26 (.A(\cpu0.b_reg[2] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0109_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold28 (.A(uo_out[2]),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0093_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold30 (.A(\cpu0.ram[4][7] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold31 (.A(\cpu0.ram[13][1] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold32 (.A(uo_out[4]),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0095_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cpu0.ram[13][4] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold35 (.A(\cpu0.ram[4][0] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cpu0.b_reg[6] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold37 (.A(\cpu0.ram[8][7] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold38 (.A(\cpu0.ram[5][4] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold39 (.A(\cpu0.ram[0][4] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold40 (.A(\cpu0.ram[9][1] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold41 (.A(\cpu0.ram[15][7] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold42 (.A(\cpu0.ram[11][2] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cpu0.ram[13][0] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cpu0.ram[5][6] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold45 (.A(\cpu0.ram[1][5] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold46 (.A(\cpu0.ram[1][2] ),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold47 (.A(\cpu0.ram[1][1] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold48 (.A(\cpu0.ram[11][6] ),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold49 (.A(uo_out[1]),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0092_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold51 (.A(\cpu0.ram[13][2] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold52 (.A(\cpu0.ram[7][5] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold53 (.A(\cpu0.ram[12][6] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold54 (.A(\cpu0.ram[0][0] ),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold55 (.A(\cpu0.ram[12][1] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold56 (.A(\cpu0.ram[1][4] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold57 (.A(\cpu0.ram[14][6] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold58 (.A(\cpu0.ram[14][3] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold59 (.A(\cpu0.ram[4][2] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold60 (.A(\cpu0.ram[5][3] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold61 (.A(\cpu0.ram[14][0] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold62 (.A(\cpu0.ram[3][7] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold63 (.A(\cpu0.ram[3][0] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold64 (.A(\cpu0.ram[6][2] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold65 (.A(\cpu0.ram[8][2] ),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold66 (.A(\cpu0.ram[15][4] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold67 (.A(\cpu0.ram[8][1] ),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold68 (.A(\cpu0.ram[11][4] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold69 (.A(\cpu0.ram[7][3] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold70 (.A(\cpu0.ram[9][2] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold71 (.A(\cpu0.ram[13][5] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold72 (.A(\cpu0.ram[6][4] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold73 (.A(\cpu0.ram[11][5] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold74 (.A(\cpu0.ram[2][4] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold75 (.A(\cpu0.ram[3][1] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold76 (.A(\cpu0.ram[12][5] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold77 (.A(\cpu0.ram[0][5] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold78 (.A(\cpu0.ram[7][6] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold79 (.A(\cpu0.ram[12][3] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold80 (.A(\cpu0.ram[5][7] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold81 (.A(\cpu0.ram[10][5] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold82 (.A(\cpu0.ram[10][3] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold83 (.A(\cpu0.ram[10][0] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold84 (.A(\cpu0.b_reg[3] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0110_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold86 (.A(\cpu0.ram[11][0] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold87 (.A(\cpu0.ram[12][0] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold88 (.A(\cpu0.ram[4][3] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold89 (.A(\cpu0.ram[12][2] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold90 (.A(\cpu0.ram[3][6] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold91 (.A(\cpu0.ram[6][0] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold92 (.A(\cpu0.ram[3][3] ),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold93 (.A(\cpu0.ram[5][5] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold94 (.A(\cpu0.ram[13][6] ),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold95 (.A(\cpu0.ram[6][3] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cpu0.ram[15][5] ),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold97 (.A(\cpu0.ram[2][3] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold98 (.A(\cpu0.b_reg[1] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0108_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold100 (.A(\cpu0.ram[7][7] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold101 (.A(\cpu0.ram[4][6] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold102 (.A(\cpu0.ram[7][4] ),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cpu0.ram[14][7] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold104 (.A(\cpu0.ram[5][0] ),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold105 (.A(\cpu0.ram[10][1] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold106 (.A(\cpu0.ram[9][5] ),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cpu0.ram[6][7] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold108 (.A(\cpu0.ram[15][3] ),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold109 (.A(\cpu0.ram[14][5] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold110 (.A(\cpu0.ram[6][1] ),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold111 (.A(\cpu0.ram[6][5] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold112 (.A(\cpu0.ram[14][1] ),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold113 (.A(\cpu0.ram[2][0] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold114 (.A(\cpu0.ram[12][7] ),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold115 (.A(\cpu0.ram[1][7] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold116 (.A(\cpu0.ram[13][7] ),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold117 (.A(\cpu0.ram[8][6] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold118 (.A(\cpu0.ram[4][1] ),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold119 (.A(\cpu0.ram[14][4] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold120 (.A(\cpu0.ram[15][6] ),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold121 (.A(\cpu0.ram[2][2] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold122 (.A(\cpu0.ram[2][5] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold123 (.A(\cpu0.ram[9][0] ),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold124 (.A(\cpu0.ram[2][1] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold125 (.A(\cpu0.ram[10][2] ),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold126 (.A(\cpu0.ram[3][5] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold127 (.A(\cpu0.b_reg[4] ),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold128 (.A(\cpu0.ram[9][6] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold129 (.A(\cpu0.ram[15][0] ),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold130 (.A(\cpu0.ram[11][7] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold131 (.A(\cpu0.ram[8][4] ),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold132 (.A(\cpu0.ram[12][4] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold133 (.A(\cpu0.ram[8][0] ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold134 (.A(\cpu0.ram[10][6] ),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold135 (.A(\cpu0.ram[2][6] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold136 (.A(\cpu0.ram[9][7] ),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold137 (.A(\cpu0.ram[14][2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold138 (.A(\cpu0.ram[8][5] ),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold139 (.A(\cpu0.ram[0][6] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold140 (.A(\cpu0.ram[1][0] ),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold141 (.A(\cpu0.ram[3][4] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold142 (.A(\cpu0.ram[8][3] ),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold143 (.A(\cpu0.ram[5][1] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold144 (.A(\cpu0.ram[6][6] ),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold145 (.A(\cpu0.ram[9][4] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold146 (.A(\cpu0.ram[2][7] ),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold147 (.A(uo_out[5]),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold148 (.A(_0545_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold149 (.A(\cpu0.ram[10][7] ),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold150 (.A(\cpu0.ram[0][7] ),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold151 (.A(\cpu0.ram[1][3] ),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold152 (.A(\cpu0.ram[1][6] ),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold153 (.A(\cpu0.ram[7][1] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold154 (.A(\cpu0.ram[0][1] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold155 (.A(\cpu0.ram[0][2] ),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold156 (.A(\cpu0.ram[10][4] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold157 (.A(\cpu0.ram[4][5] ),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold158 (.A(\cpu0.ram[4][4] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold159 (.A(\cpu0.ram[0][3] ),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold160 (.A(\cpu0.ram[7][0] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold161 (.A(uo_out[0]),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0540_),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold163 (.A(\cpu0.ram[15][2] ),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold164 (.A(\cpu0.b_reg[0] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold165 (.A(_0107_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold166 (.A(\cpu0.ram[7][2] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold167 (.A(\cpu0.ir[4] ),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold168 (.A(\cpu0.a_reg[5] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold169 (.A(\cpu0.pc[0] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0163_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold171 (.A(\cpu0.ir[5] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0536_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold173 (.A(\cpu0.ir[6] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold174 (.A(\cpu0.a_reg[4] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold175 (.A(\cpu0.ir[7] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0090_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold177 (.A(\cpu0.step[0] ),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0218_),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold179 (.A(_0024_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold180 (.A(\cpu0.a_reg[1] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0100_),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold182 (.A(\cpu0.b_reg[5] ),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0569_),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold184 (.A(\cpu0.pc[1] ),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0590_),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold186 (.A(\cpu0.pc[2] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0596_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold188 (.A(\cpu0.pc[3] ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold189 (.A(\cpu0.a_reg[3] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold190 (.A(\cpu0.mar[3] ),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold191 (.A(\cpu0.mar[2] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold192 (.A(\cpu0.a_reg[0] ),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold193 (.A(\cpu0.a_reg[2] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold194 (.A(\cpu0.mar[0] ),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold195 (.A(\cpu0.step[2] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold196 (.A(\cpu0.mar[1] ),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold197 (.A(\cpu0.a_reg[7] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold198 (.A(\cpu0.a_reg[6] ),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold199 (.A(\cpu0.step[1] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold200 (.A(\cpu0.step[2] ),
    .X(net473));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_4 FILLER_0_105 ();
 sg13g2_fill_1 FILLER_0_109 ();
 sg13g2_decap_8 FILLER_0_114 ();
 sg13g2_decap_8 FILLER_0_121 ();
 sg13g2_decap_8 FILLER_0_128 ();
 sg13g2_decap_8 FILLER_0_135 ();
 sg13g2_decap_8 FILLER_0_142 ();
 sg13g2_decap_4 FILLER_0_149 ();
 sg13g2_fill_2 FILLER_0_167 ();
 sg13g2_fill_1 FILLER_0_169 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_4 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_fill_2 FILLER_0_249 ();
 sg13g2_fill_1 FILLER_0_251 ();
 sg13g2_decap_4 FILLER_0_256 ();
 sg13g2_fill_1 FILLER_0_260 ();
 sg13g2_decap_8 FILLER_0_288 ();
 sg13g2_decap_4 FILLER_0_295 ();
 sg13g2_decap_4 FILLER_0_309 ();
 sg13g2_fill_2 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_fill_2 FILLER_0_345 ();
 sg13g2_fill_2 FILLER_0_356 ();
 sg13g2_fill_1 FILLER_0_358 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_fill_2 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_4 FILLER_1_91 ();
 sg13g2_fill_1 FILLER_1_95 ();
 sg13g2_decap_8 FILLER_1_132 ();
 sg13g2_decap_4 FILLER_1_139 ();
 sg13g2_decap_8 FILLER_1_183 ();
 sg13g2_fill_1 FILLER_1_190 ();
 sg13g2_fill_2 FILLER_1_201 ();
 sg13g2_fill_1 FILLER_1_203 ();
 sg13g2_decap_4 FILLER_1_241 ();
 sg13g2_fill_2 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_292 ();
 sg13g2_fill_1 FILLER_1_299 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_fill_2 FILLER_1_334 ();
 sg13g2_fill_1 FILLER_1_336 ();
 sg13g2_fill_2 FILLER_1_364 ();
 sg13g2_fill_1 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_4 FILLER_2_77 ();
 sg13g2_fill_1 FILLER_2_81 ();
 sg13g2_fill_1 FILLER_2_109 ();
 sg13g2_fill_1 FILLER_2_137 ();
 sg13g2_fill_1 FILLER_2_175 ();
 sg13g2_fill_2 FILLER_2_186 ();
 sg13g2_fill_1 FILLER_2_239 ();
 sg13g2_decap_4 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_30 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_fill_2 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_44 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_4 FILLER_3_77 ();
 sg13g2_fill_1 FILLER_3_81 ();
 sg13g2_fill_2 FILLER_3_96 ();
 sg13g2_decap_8 FILLER_3_131 ();
 sg13g2_fill_1 FILLER_3_138 ();
 sg13g2_fill_2 FILLER_3_166 ();
 sg13g2_fill_1 FILLER_3_215 ();
 sg13g2_fill_2 FILLER_3_244 ();
 sg13g2_fill_1 FILLER_3_266 ();
 sg13g2_decap_4 FILLER_3_294 ();
 sg13g2_fill_1 FILLER_3_325 ();
 sg13g2_fill_2 FILLER_3_349 ();
 sg13g2_fill_1 FILLER_3_371 ();
 sg13g2_fill_2 FILLER_3_376 ();
 sg13g2_fill_1 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_4 FILLER_4_7 ();
 sg13g2_fill_2 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_4 FILLER_4_88 ();
 sg13g2_decap_4 FILLER_4_102 ();
 sg13g2_fill_1 FILLER_4_106 ();
 sg13g2_fill_1 FILLER_4_120 ();
 sg13g2_fill_1 FILLER_4_125 ();
 sg13g2_fill_1 FILLER_4_176 ();
 sg13g2_fill_1 FILLER_4_197 ();
 sg13g2_decap_4 FILLER_4_234 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_4 FILLER_4_298 ();
 sg13g2_decap_4 FILLER_4_329 ();
 sg13g2_fill_2 FILLER_4_333 ();
 sg13g2_decap_4 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_fill_2 FILLER_5_134 ();
 sg13g2_fill_2 FILLER_5_173 ();
 sg13g2_decap_4 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_204 ();
 sg13g2_fill_1 FILLER_5_211 ();
 sg13g2_fill_1 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_fill_1 FILLER_5_242 ();
 sg13g2_fill_2 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_4 FILLER_5_291 ();
 sg13g2_fill_1 FILLER_5_295 ();
 sg13g2_fill_2 FILLER_5_300 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_fill_1 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_5_405 ();
 sg13g2_fill_1 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_38 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_fill_1 FILLER_6_79 ();
 sg13g2_fill_2 FILLER_6_117 ();
 sg13g2_fill_1 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_145 ();
 sg13g2_decap_4 FILLER_6_174 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_decap_8 FILLER_6_199 ();
 sg13g2_fill_2 FILLER_6_206 ();
 sg13g2_fill_1 FILLER_6_208 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_fill_2 FILLER_6_221 ();
 sg13g2_fill_1 FILLER_6_223 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_decap_8 FILLER_6_236 ();
 sg13g2_decap_4 FILLER_6_243 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_decap_4 FILLER_6_285 ();
 sg13g2_fill_2 FILLER_6_289 ();
 sg13g2_decap_4 FILLER_6_333 ();
 sg13g2_decap_4 FILLER_6_404 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_66 ();
 sg13g2_fill_2 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_123 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_decap_4 FILLER_7_192 ();
 sg13g2_fill_1 FILLER_7_196 ();
 sg13g2_decap_4 FILLER_7_224 ();
 sg13g2_fill_2 FILLER_7_238 ();
 sg13g2_fill_2 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_4 FILLER_7_294 ();
 sg13g2_fill_2 FILLER_7_298 ();
 sg13g2_fill_2 FILLER_7_310 ();
 sg13g2_fill_2 FILLER_7_335 ();
 sg13g2_fill_1 FILLER_7_376 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_40 ();
 sg13g2_fill_1 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_68 ();
 sg13g2_decap_4 FILLER_8_75 ();
 sg13g2_fill_1 FILLER_8_79 ();
 sg13g2_fill_2 FILLER_8_107 ();
 sg13g2_fill_1 FILLER_8_109 ();
 sg13g2_fill_2 FILLER_8_131 ();
 sg13g2_fill_1 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_164 ();
 sg13g2_fill_2 FILLER_8_175 ();
 sg13g2_fill_1 FILLER_8_177 ();
 sg13g2_decap_4 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_186 ();
 sg13g2_fill_1 FILLER_8_264 ();
 sg13g2_fill_1 FILLER_8_300 ();
 sg13g2_fill_1 FILLER_8_341 ();
 sg13g2_fill_2 FILLER_8_360 ();
 sg13g2_fill_1 FILLER_8_362 ();
 sg13g2_decap_4 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_4 ();
 sg13g2_decap_4 FILLER_9_86 ();
 sg13g2_decap_8 FILLER_9_115 ();
 sg13g2_fill_1 FILLER_9_122 ();
 sg13g2_fill_2 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_171 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_fill_2 FILLER_9_190 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_1 FILLER_9_289 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_332 ();
 sg13g2_decap_4 FILLER_9_339 ();
 sg13g2_fill_2 FILLER_9_356 ();
 sg13g2_fill_1 FILLER_9_358 ();
 sg13g2_fill_2 FILLER_9_367 ();
 sg13g2_fill_1 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_4 FILLER_9_403 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_decap_8 FILLER_10_79 ();
 sg13g2_decap_4 FILLER_10_86 ();
 sg13g2_fill_2 FILLER_10_90 ();
 sg13g2_fill_1 FILLER_10_124 ();
 sg13g2_fill_2 FILLER_10_166 ();
 sg13g2_decap_4 FILLER_10_177 ();
 sg13g2_fill_2 FILLER_10_181 ();
 sg13g2_fill_2 FILLER_10_193 ();
 sg13g2_decap_4 FILLER_10_208 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_decap_4 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_237 ();
 sg13g2_decap_8 FILLER_10_285 ();
 sg13g2_fill_2 FILLER_10_292 ();
 sg13g2_fill_1 FILLER_10_294 ();
 sg13g2_fill_2 FILLER_10_331 ();
 sg13g2_fill_1 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_365 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_4 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_4 ();
 sg13g2_fill_1 FILLER_11_9 ();
 sg13g2_fill_2 FILLER_11_37 ();
 sg13g2_fill_1 FILLER_11_66 ();
 sg13g2_decap_4 FILLER_11_76 ();
 sg13g2_fill_1 FILLER_11_134 ();
 sg13g2_fill_1 FILLER_11_148 ();
 sg13g2_fill_2 FILLER_11_176 ();
 sg13g2_fill_1 FILLER_11_178 ();
 sg13g2_decap_4 FILLER_11_214 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_fill_1 FILLER_11_255 ();
 sg13g2_decap_4 FILLER_11_270 ();
 sg13g2_fill_2 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_285 ();
 sg13g2_fill_2 FILLER_11_297 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_decap_4 FILLER_11_304 ();
 sg13g2_fill_1 FILLER_11_308 ();
 sg13g2_fill_1 FILLER_11_314 ();
 sg13g2_fill_1 FILLER_11_328 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_117 ();
 sg13g2_fill_2 FILLER_12_124 ();
 sg13g2_fill_1 FILLER_12_135 ();
 sg13g2_fill_1 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_174 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_fill_2 FILLER_12_215 ();
 sg13g2_fill_2 FILLER_12_244 ();
 sg13g2_decap_4 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_306 ();
 sg13g2_fill_1 FILLER_12_313 ();
 sg13g2_fill_1 FILLER_12_350 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_fill_2 FILLER_13_29 ();
 sg13g2_fill_2 FILLER_13_40 ();
 sg13g2_fill_1 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_73 ();
 sg13g2_decap_8 FILLER_13_80 ();
 sg13g2_fill_2 FILLER_13_87 ();
 sg13g2_decap_4 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_decap_8 FILLER_13_124 ();
 sg13g2_fill_1 FILLER_13_136 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_4 FILLER_13_186 ();
 sg13g2_fill_2 FILLER_13_239 ();
 sg13g2_fill_2 FILLER_13_246 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_fill_2 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_280 ();
 sg13g2_fill_2 FILLER_13_318 ();
 sg13g2_fill_1 FILLER_13_366 ();
 sg13g2_decap_4 FILLER_13_404 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_4 FILLER_14_14 ();
 sg13g2_fill_1 FILLER_14_18 ();
 sg13g2_fill_1 FILLER_14_29 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_68 ();
 sg13g2_decap_4 FILLER_14_75 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_4 FILLER_14_177 ();
 sg13g2_fill_2 FILLER_14_212 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_4 FILLER_14_230 ();
 sg13g2_decap_4 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_247 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_decap_8 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_fill_2 FILLER_14_366 ();
 sg13g2_fill_1 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_4 FILLER_15_14 ();
 sg13g2_fill_1 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_50 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_59 ();
 sg13g2_decap_4 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_fill_2 FILLER_15_127 ();
 sg13g2_fill_1 FILLER_15_129 ();
 sg13g2_fill_1 FILLER_15_135 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_2 FILLER_15_202 ();
 sg13g2_fill_1 FILLER_15_226 ();
 sg13g2_fill_2 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_233 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_1 FILLER_15_282 ();
 sg13g2_decap_8 FILLER_15_297 ();
 sg13g2_fill_2 FILLER_15_304 ();
 sg13g2_fill_1 FILLER_15_306 ();
 sg13g2_decap_4 FILLER_15_311 ();
 sg13g2_fill_2 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_365 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_fill_2 FILLER_16_114 ();
 sg13g2_fill_1 FILLER_16_164 ();
 sg13g2_decap_8 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_196 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_decap_8 FILLER_16_212 ();
 sg13g2_decap_8 FILLER_16_219 ();
 sg13g2_decap_8 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_235 ();
 sg13g2_fill_1 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_249 ();
 sg13g2_fill_1 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_351 ();
 sg13g2_fill_2 FILLER_16_391 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_1 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_166 ();
 sg13g2_decap_4 FILLER_17_173 ();
 sg13g2_fill_1 FILLER_17_177 ();
 sg13g2_fill_2 FILLER_17_182 ();
 sg13g2_fill_1 FILLER_17_188 ();
 sg13g2_decap_4 FILLER_17_198 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_213 ();
 sg13g2_decap_8 FILLER_17_220 ();
 sg13g2_fill_1 FILLER_17_227 ();
 sg13g2_fill_1 FILLER_17_232 ();
 sg13g2_decap_4 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_260 ();
 sg13g2_fill_1 FILLER_17_262 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_345 ();
 sg13g2_fill_2 FILLER_17_352 ();
 sg13g2_fill_1 FILLER_17_354 ();
 sg13g2_fill_2 FILLER_17_375 ();
 sg13g2_decap_4 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_64 ();
 sg13g2_decap_8 FILLER_18_108 ();
 sg13g2_decap_8 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_1 FILLER_18_164 ();
 sg13g2_decap_4 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_174 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_fill_2 FILLER_18_227 ();
 sg13g2_fill_1 FILLER_18_229 ();
 sg13g2_fill_2 FILLER_18_272 ();
 sg13g2_fill_1 FILLER_18_274 ();
 sg13g2_fill_2 FILLER_18_283 ();
 sg13g2_fill_1 FILLER_18_285 ();
 sg13g2_fill_1 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_1 FILLER_18_345 ();
 sg13g2_fill_2 FILLER_18_350 ();
 sg13g2_fill_1 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_fill_2 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_fill_2 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_78 ();
 sg13g2_decap_8 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_decap_8 FILLER_19_149 ();
 sg13g2_fill_2 FILLER_19_156 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_decap_4 FILLER_19_196 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_293 ();
 sg13g2_decap_8 FILLER_19_300 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_fill_2 FILLER_19_329 ();
 sg13g2_fill_2 FILLER_19_368 ();
 sg13g2_fill_1 FILLER_19_370 ();
 sg13g2_fill_1 FILLER_19_384 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_decap_4 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_9 ();
 sg13g2_fill_2 FILLER_20_14 ();
 sg13g2_fill_1 FILLER_20_16 ();
 sg13g2_decap_8 FILLER_20_50 ();
 sg13g2_decap_8 FILLER_20_57 ();
 sg13g2_decap_4 FILLER_20_64 ();
 sg13g2_decap_4 FILLER_20_100 ();
 sg13g2_fill_2 FILLER_20_117 ();
 sg13g2_decap_4 FILLER_20_152 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_199 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_decap_4 FILLER_20_213 ();
 sg13g2_fill_2 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_223 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_decap_4 FILLER_20_307 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_75 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_4 FILLER_21_164 ();
 sg13g2_decap_8 FILLER_21_188 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_4 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_285 ();
 sg13g2_fill_1 FILLER_21_287 ();
 sg13g2_decap_4 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_300 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_fill_1 FILLER_21_355 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_decap_4 FILLER_22_58 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_fill_2 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_79 ();
 sg13g2_decap_4 FILLER_22_153 ();
 sg13g2_fill_2 FILLER_22_157 ();
 sg13g2_fill_1 FILLER_22_213 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_fill_2 FILLER_22_249 ();
 sg13g2_fill_1 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_316 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_1 FILLER_22_354 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_4 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_71 ();
 sg13g2_decap_4 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_2 FILLER_23_87 ();
 sg13g2_fill_2 FILLER_23_93 ();
 sg13g2_decap_4 FILLER_23_104 ();
 sg13g2_fill_2 FILLER_23_144 ();
 sg13g2_fill_1 FILLER_23_146 ();
 sg13g2_fill_2 FILLER_23_182 ();
 sg13g2_fill_1 FILLER_23_184 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_238 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_342 ();
 sg13g2_decap_4 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_375 ();
 sg13g2_decap_4 FILLER_23_405 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_9 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_67 ();
 sg13g2_fill_2 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_4 FILLER_24_152 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_4 FILLER_24_233 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_4 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_350 ();
 sg13g2_decap_4 FILLER_24_357 ();
 sg13g2_fill_1 FILLER_24_361 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_51 ();
 sg13g2_decap_8 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_65 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_193 ();
 sg13g2_decap_4 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_208 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_decap_4 FILLER_25_229 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_decap_4 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_281 ();
 sg13g2_decap_4 FILLER_25_288 ();
 sg13g2_fill_2 FILLER_25_320 ();
 sg13g2_decap_4 FILLER_25_331 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_353 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_64 ();
 sg13g2_fill_2 FILLER_26_85 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_fill_2 FILLER_26_222 ();
 sg13g2_fill_1 FILLER_26_224 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_8 FILLER_26_271 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_fill_1 FILLER_26_362 ();
 sg13g2_fill_2 FILLER_26_382 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_61 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_107 ();
 sg13g2_decap_8 FILLER_27_121 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_fill_2 FILLER_27_331 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_decap_4 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_fill_2 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_54 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_120 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_134 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_fill_2 FILLER_28_173 ();
 sg13g2_fill_2 FILLER_28_199 ();
 sg13g2_fill_2 FILLER_28_270 ();
 sg13g2_fill_2 FILLER_28_318 ();
 sg13g2_fill_1 FILLER_28_320 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_4 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_371 ();
 sg13g2_fill_1 FILLER_28_386 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_11 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_222 ();
 sg13g2_fill_2 FILLER_29_229 ();
 sg13g2_decap_4 FILLER_29_269 ();
 sg13g2_fill_2 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_302 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_decap_4 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_334 ();
 sg13g2_decap_4 FILLER_29_340 ();
 sg13g2_decap_4 FILLER_29_367 ();
 sg13g2_decap_4 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_111 ();
 sg13g2_decap_4 FILLER_30_118 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_fill_2 FILLER_30_231 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_fill_2 FILLER_30_248 ();
 sg13g2_decap_4 FILLER_30_268 ();
 sg13g2_decap_8 FILLER_30_285 ();
 sg13g2_fill_2 FILLER_30_299 ();
 sg13g2_decap_4 FILLER_30_306 ();
 sg13g2_decap_8 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_59 ();
 sg13g2_fill_2 FILLER_31_107 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_1 FILLER_31_146 ();
 sg13g2_fill_2 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_216 ();
 sg13g2_decap_4 FILLER_31_222 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_258 ();
 sg13g2_fill_1 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_297 ();
 sg13g2_fill_1 FILLER_31_299 ();
 sg13g2_fill_1 FILLER_31_335 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_58 ();
 sg13g2_decap_8 FILLER_32_65 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_103 ();
 sg13g2_fill_2 FILLER_32_194 ();
 sg13g2_decap_8 FILLER_32_211 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_4 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_2 FILLER_32_324 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_decap_4 FILLER_32_344 ();
 sg13g2_fill_2 FILLER_32_348 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_373 ();
 sg13g2_fill_2 FILLER_32_392 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_10 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_fill_1 FILLER_33_34 ();
 sg13g2_decap_4 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_fill_2 FILLER_33_74 ();
 sg13g2_fill_1 FILLER_33_124 ();
 sg13g2_fill_1 FILLER_33_202 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_fill_1 FILLER_33_220 ();
 sg13g2_fill_1 FILLER_33_236 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_fill_1 FILLER_33_310 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_fill_1 FILLER_33_341 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_fill_1 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_12 ();
 sg13g2_decap_8 FILLER_34_41 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_118 ();
 sg13g2_fill_2 FILLER_34_166 ();
 sg13g2_fill_2 FILLER_34_220 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_fill_2 FILLER_34_279 ();
 sg13g2_fill_1 FILLER_34_281 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_324 ();
 sg13g2_fill_2 FILLER_34_353 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_decap_8 FILLER_35_290 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_1 FILLER_35_376 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_4 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_18 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_fill_1 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_1 FILLER_36_101 ();
 sg13g2_fill_1 FILLER_36_138 ();
 sg13g2_fill_1 FILLER_36_148 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_306 ();
 sg13g2_fill_2 FILLER_36_341 ();
 sg13g2_fill_2 FILLER_36_357 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_79 ();
 sg13g2_fill_1 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_113 ();
 sg13g2_fill_2 FILLER_37_198 ();
 sg13g2_fill_2 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_239 ();
 sg13g2_decap_8 FILLER_37_292 ();
 sg13g2_decap_4 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_384 ();
 sg13g2_fill_1 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_59 ();
 sg13g2_fill_2 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_80 ();
 sg13g2_fill_1 FILLER_38_107 ();
 sg13g2_fill_1 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_4 FILLER_38_210 ();
 sg13g2_fill_2 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_fill_1 FILLER_38_229 ();
 sg13g2_decap_4 FILLER_38_239 ();
 sg13g2_fill_1 FILLER_38_243 ();
 sg13g2_fill_2 FILLER_38_265 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_345 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net14;
 assign uio_oe[1] = net15;
 assign uio_oe[2] = net16;
 assign uio_oe[3] = net17;
 assign uio_oe[4] = net18;
 assign uio_oe[5] = net19;
 assign uio_oe[6] = net20;
 assign uio_oe[7] = net21;
 assign uio_out[0] = net22;
 assign uio_out[1] = net23;
 assign uio_out[2] = net24;
 assign uio_out[3] = net25;
 assign uio_out[4] = net26;
 assign uio_out[5] = net27;
 assign uio_out[6] = net28;
 assign uio_out[7] = net29;
endmodule
