module tt_um_arthfink_ddmtd (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire clk_fb;
 wire clk_helper;
 wire \ctrl[0] ;
 wire \ctrl[10] ;
 wire \ctrl[11] ;
 wire \ctrl[12] ;
 wire \ctrl[13] ;
 wire \ctrl[14] ;
 wire \ctrl[15] ;
 wire \ctrl[16] ;
 wire \ctrl[17] ;
 wire \ctrl[18] ;
 wire \ctrl[19] ;
 wire \ctrl[1] ;
 wire \ctrl[20] ;
 wire \ctrl[21] ;
 wire \ctrl[22] ;
 wire \ctrl[23] ;
 wire \ctrl[2] ;
 wire \ctrl[3] ;
 wire \ctrl[8] ;
 wire \ctrl[9] ;
 wire fb_samp;
 wire helper_msb_d;
 wire \nco_phase_acc[0] ;
 wire \nco_phase_acc[10] ;
 wire \nco_phase_acc[11] ;
 wire \nco_phase_acc[12] ;
 wire \nco_phase_acc[13] ;
 wire \nco_phase_acc[14] ;
 wire \nco_phase_acc[15] ;
 wire \nco_phase_acc[16] ;
 wire \nco_phase_acc[17] ;
 wire \nco_phase_acc[18] ;
 wire \nco_phase_acc[19] ;
 wire \nco_phase_acc[1] ;
 wire \nco_phase_acc[20] ;
 wire \nco_phase_acc[21] ;
 wire \nco_phase_acc[22] ;
 wire \nco_phase_acc[2] ;
 wire \nco_phase_acc[3] ;
 wire \nco_phase_acc[4] ;
 wire \nco_phase_acc[5] ;
 wire \nco_phase_acc[6] ;
 wire \nco_phase_acc[7] ;
 wire \nco_phase_acc[8] ;
 wire \nco_phase_acc[9] ;
 wire \phase_err_beat[10] ;
 wire \phase_err_beat[11] ;
 wire \phase_err_beat[12] ;
 wire \phase_err_beat[13] ;
 wire \phase_err_beat[14] ;
 wire \phase_err_beat[15] ;
 wire \phase_err_beat[4] ;
 wire \phase_err_beat[5] ;
 wire \phase_err_beat[6] ;
 wire \phase_err_beat[7] ;
 wire \phase_err_beat[8] ;
 wire \phase_err_beat[9] ;
 wire phase_valid;
 wire ref_samp;
 wire \u_core.beat_cnt[0] ;
 wire \u_core.beat_cnt[10] ;
 wire \u_core.beat_cnt[11] ;
 wire \u_core.beat_cnt[12] ;
 wire \u_core.beat_cnt[13] ;
 wire \u_core.beat_cnt[14] ;
 wire \u_core.beat_cnt[15] ;
 wire \u_core.beat_cnt[1] ;
 wire \u_core.beat_cnt[2] ;
 wire \u_core.beat_cnt[3] ;
 wire \u_core.beat_cnt[4] ;
 wire \u_core.beat_cnt[5] ;
 wire \u_core.beat_cnt[6] ;
 wire \u_core.beat_cnt[7] ;
 wire \u_core.beat_cnt[8] ;
 wire \u_core.beat_cnt[9] ;
 wire \u_core.fb_samp_d ;
 wire \u_core.fb_sync[0] ;
 wire \u_core.fb_sync[1] ;
 wire \u_core.have_fb ;
 wire \u_core.have_ref ;
 wire \u_core.ref_samp_d ;
 wire \u_core.ref_sync[0] ;
 wire \u_core.ref_sync[1] ;
 wire \u_core.t_fb[0] ;
 wire \u_core.t_fb[10] ;
 wire \u_core.t_fb[11] ;
 wire \u_core.t_fb[12] ;
 wire \u_core.t_fb[13] ;
 wire \u_core.t_fb[14] ;
 wire \u_core.t_fb[15] ;
 wire \u_core.t_fb[1] ;
 wire \u_core.t_fb[2] ;
 wire \u_core.t_fb[3] ;
 wire \u_core.t_fb[4] ;
 wire \u_core.t_fb[5] ;
 wire \u_core.t_fb[6] ;
 wire \u_core.t_fb[7] ;
 wire \u_core.t_fb[8] ;
 wire \u_core.t_fb[9] ;
 wire \u_core.t_ref[0] ;
 wire \u_core.t_ref[10] ;
 wire \u_core.t_ref[11] ;
 wire \u_core.t_ref[12] ;
 wire \u_core.t_ref[13] ;
 wire \u_core.t_ref[14] ;
 wire \u_core.t_ref[15] ;
 wire \u_core.t_ref[1] ;
 wire \u_core.t_ref[2] ;
 wire \u_core.t_ref[3] ;
 wire \u_core.t_ref[4] ;
 wire \u_core.t_ref[5] ;
 wire \u_core.t_ref[6] ;
 wire \u_core.t_ref[7] ;
 wire \u_core.t_ref[8] ;
 wire \u_core.t_ref[9] ;
 wire \u_lf.i_acc[0] ;
 wire \u_lf.i_acc[10] ;
 wire \u_lf.i_acc[11] ;
 wire \u_lf.i_acc[12] ;
 wire \u_lf.i_acc[13] ;
 wire \u_lf.i_acc[14] ;
 wire \u_lf.i_acc[15] ;
 wire \u_lf.i_acc[16] ;
 wire \u_lf.i_acc[17] ;
 wire \u_lf.i_acc[18] ;
 wire \u_lf.i_acc[19] ;
 wire \u_lf.i_acc[1] ;
 wire \u_lf.i_acc[20] ;
 wire \u_lf.i_acc[21] ;
 wire \u_lf.i_acc[22] ;
 wire \u_lf.i_acc[23] ;
 wire \u_lf.i_acc[24] ;
 wire \u_lf.i_acc[25] ;
 wire \u_lf.i_acc[26] ;
 wire \u_lf.i_acc[27] ;
 wire \u_lf.i_acc[28] ;
 wire \u_lf.i_acc[29] ;
 wire \u_lf.i_acc[2] ;
 wire \u_lf.i_acc[3] ;
 wire \u_lf.i_acc[4] ;
 wire \u_lf.i_acc[5] ;
 wire \u_lf.i_acc[6] ;
 wire \u_lf.i_acc[7] ;
 wire \u_lf.i_acc[8] ;
 wire \u_lf.i_acc[9] ;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;

 sg13g2_inv_1 _0638_ (.Y(_0141_),
    .A(net210));
 sg13g2_inv_1 _0639_ (.Y(_0142_),
    .A(net57));
 sg13g2_inv_1 _0640_ (.Y(_0143_),
    .A(net107));
 sg13g2_inv_1 _0641_ (.Y(_0144_),
    .A(net41));
 sg13g2_inv_1 _0642_ (.Y(_0145_),
    .A(net45));
 sg13g2_inv_1 _0643_ (.Y(_0146_),
    .A(net63));
 sg13g2_inv_1 _0644_ (.Y(_0147_),
    .A(net56));
 sg13g2_inv_1 _0645_ (.Y(_0148_),
    .A(net293));
 sg13g2_inv_1 _0646_ (.Y(_0149_),
    .A(net274));
 sg13g2_inv_1 _0647_ (.Y(_0150_),
    .A(net243));
 sg13g2_inv_1 _0648_ (.Y(_0151_),
    .A(net270));
 sg13g2_inv_1 _0649_ (.Y(_0152_),
    .A(net114));
 sg13g2_inv_1 _0650_ (.Y(_0153_),
    .A(\u_core.t_ref[5] ));
 sg13g2_inv_1 _0651_ (.Y(_0154_),
    .A(net96));
 sg13g2_inv_1 _0652_ (.Y(_0155_),
    .A(net66));
 sg13g2_inv_1 _0653_ (.Y(_0156_),
    .A(\u_core.t_fb[13] ));
 sg13g2_inv_1 _0654_ (.Y(_0157_),
    .A(net91));
 sg13g2_inv_1 _0655_ (.Y(_0158_),
    .A(net27));
 sg13g2_inv_1 _0656_ (.Y(_0159_),
    .A(net23));
 sg13g2_inv_1 _0657_ (.Y(_0160_),
    .A(net25));
 sg13g2_inv_1 _0658_ (.Y(_0161_),
    .A(net128));
 sg13g2_inv_1 _0659_ (.Y(_0162_),
    .A(net67));
 sg13g2_inv_1 _0660_ (.Y(_0163_),
    .A(net102));
 sg13g2_inv_1 _0661_ (.Y(_0164_),
    .A(net48));
 sg13g2_inv_1 _0662_ (.Y(_0165_),
    .A(net104));
 sg13g2_inv_1 _0663_ (.Y(_0166_),
    .A(net83));
 sg13g2_inv_1 _0664_ (.Y(_0167_),
    .A(net222));
 sg13g2_inv_1 _0665_ (.Y(_0168_),
    .A(net93));
 sg13g2_inv_1 _0666_ (.Y(_0169_),
    .A(net119));
 sg13g2_inv_1 _0667_ (.Y(_0170_),
    .A(net136));
 sg13g2_inv_1 _0668_ (.Y(_0171_),
    .A(net140));
 sg13g2_inv_1 _0669_ (.Y(_0172_),
    .A(net70));
 sg13g2_inv_1 _0670_ (.Y(_0173_),
    .A(net95));
 sg13g2_inv_1 _0671_ (.Y(_0174_),
    .A(\nco_phase_acc[11] ));
 sg13g2_inv_1 _0672_ (.Y(_0175_),
    .A(net282));
 sg13g2_inv_1 _0673_ (.Y(_0176_),
    .A(net97));
 sg13g2_inv_1 _0674_ (.Y(_0177_),
    .A(net89));
 sg13g2_inv_1 _0675_ (.Y(_0178_),
    .A(net112));
 sg13g2_inv_1 _0676_ (.Y(_0179_),
    .A(net121));
 sg13g2_inv_1 _0677_ (.Y(_0180_),
    .A(net76));
 sg13g2_xor2_1 _0678_ (.B(helper_msb_d),
    .A(net22),
    .X(_0181_));
 sg13g2_and2_1 _0679_ (.A(net210),
    .B(_0181_),
    .X(_0182_));
 sg13g2_nand3_1 _0680_ (.B(net276),
    .C(_0182_),
    .A(net263),
    .Y(_0183_));
 sg13g2_inv_2 _0681_ (.Y(_0000_),
    .A(net156));
 sg13g2_nand2_1 _0682_ (.Y(_0184_),
    .A(net209),
    .B(phase_valid));
 sg13g2_inv_1 _0683_ (.Y(net164),
    .A(net169));
 sg13g2_mux2_1 _0684_ (.A0(net2),
    .A1(net22),
    .S(net3),
    .X(clk_fb));
 sg13g2_and2_1 _0685_ (.A(net210),
    .B(ref_samp),
    .X(uo_out[1]));
 sg13g2_and2_1 _0686_ (.A(net210),
    .B(fb_samp),
    .X(uo_out[2]));
 sg13g2_and2_1 _0687_ (.A(net210),
    .B(net3),
    .X(uo_out[3]));
 sg13g2_nor2_1 _0688_ (.A(net182),
    .B(_0144_),
    .Y(uo_out[4]));
 sg13g2_nor2_1 _0689_ (.A(net182),
    .B(_0145_),
    .Y(uo_out[5]));
 sg13g2_nor2_1 _0690_ (.A(net182),
    .B(_0146_),
    .Y(uo_out[6]));
 sg13g2_nor2_1 _0691_ (.A(net182),
    .B(_0147_),
    .Y(uo_out[7]));
 sg13g2_nand2_1 _0692_ (.Y(_0185_),
    .A(_0181_),
    .B(uo_out[1]));
 sg13g2_o21ai_1 _0693_ (.B1(_0185_),
    .Y(_0001_),
    .A1(_0143_),
    .A2(_0182_));
 sg13g2_xor2_1 _0694_ (.B(_0182_),
    .A(net42),
    .X(_0002_));
 sg13g2_nand3_1 _0695_ (.B(net308),
    .C(_0182_),
    .A(net42),
    .Y(_0186_));
 sg13g2_a21o_1 _0696_ (.A2(_0182_),
    .A1(net42),
    .B1(net308),
    .X(_0187_));
 sg13g2_and2_1 _0697_ (.A(_0186_),
    .B(_0187_),
    .X(_0003_));
 sg13g2_nor2_2 _0698_ (.A(_0158_),
    .B(_0186_),
    .Y(_0188_));
 sg13g2_xnor2_1 _0699_ (.Y(_0004_),
    .A(net27),
    .B(_0186_));
 sg13g2_xor2_1 _0700_ (.B(_0188_),
    .A(net54),
    .X(_0005_));
 sg13g2_nand3_1 _0701_ (.B(net280),
    .C(_0188_),
    .A(net54),
    .Y(_0189_));
 sg13g2_a21o_1 _0702_ (.A2(_0188_),
    .A1(net54),
    .B1(net280),
    .X(_0190_));
 sg13g2_and2_1 _0703_ (.A(_0189_),
    .B(_0190_),
    .X(_0006_));
 sg13g2_nor2_1 _0704_ (.A(_0159_),
    .B(_0189_),
    .Y(_0191_));
 sg13g2_xnor2_1 _0705_ (.Y(_0007_),
    .A(net23),
    .B(_0189_));
 sg13g2_xor2_1 _0706_ (.B(_0191_),
    .A(net52),
    .X(_0008_));
 sg13g2_nand3_1 _0707_ (.B(net311),
    .C(_0191_),
    .A(net52),
    .Y(_0192_));
 sg13g2_a21o_1 _0708_ (.A2(_0191_),
    .A1(net52),
    .B1(net311),
    .X(_0193_));
 sg13g2_and2_1 _0709_ (.A(_0192_),
    .B(_0193_),
    .X(_0009_));
 sg13g2_nor2_1 _0710_ (.A(_0160_),
    .B(_0192_),
    .Y(_0194_));
 sg13g2_xnor2_1 _0711_ (.Y(_0010_),
    .A(net25),
    .B(_0192_));
 sg13g2_and2_1 _0712_ (.A(net35),
    .B(_0194_),
    .X(_0195_));
 sg13g2_xor2_1 _0713_ (.B(_0194_),
    .A(net35),
    .X(_0011_));
 sg13g2_xor2_1 _0714_ (.B(_0195_),
    .A(net46),
    .X(_0012_));
 sg13g2_and3_2 _0715_ (.X(_0196_),
    .A(net46),
    .B(net69),
    .C(_0195_));
 sg13g2_a21oi_1 _0716_ (.A1(net46),
    .A2(_0195_),
    .Y(_0197_),
    .B1(net69));
 sg13g2_nor2_1 _0717_ (.A(_0196_),
    .B(_0197_),
    .Y(_0013_));
 sg13g2_xor2_1 _0718_ (.B(_0196_),
    .A(net59),
    .X(_0014_));
 sg13g2_nand3_1 _0719_ (.B(net85),
    .C(_0196_),
    .A(net59),
    .Y(_0198_));
 sg13g2_a21o_1 _0720_ (.A2(_0196_),
    .A1(net59),
    .B1(net85),
    .X(_0199_));
 sg13g2_and2_1 _0721_ (.A(_0198_),
    .B(_0199_),
    .X(_0015_));
 sg13g2_nand4_1 _0722_ (.B(\u_core.beat_cnt[13] ),
    .C(\u_core.beat_cnt[14] ),
    .A(\u_core.beat_cnt[12] ),
    .Y(_0200_),
    .D(_0196_));
 sg13g2_xnor2_1 _0723_ (.Y(_0016_),
    .A(net61),
    .B(_0198_));
 sg13g2_xnor2_1 _0724_ (.Y(_0017_),
    .A(net43),
    .B(_0200_));
 sg13g2_nor2b_1 _0725_ (.A(\u_core.t_ref[4] ),
    .B_N(\u_core.t_fb[4] ),
    .Y(_0201_));
 sg13g2_xnor2_1 _0726_ (.Y(_0202_),
    .A(\u_core.t_fb[4] ),
    .B(\u_core.t_ref[4] ));
 sg13g2_nor2b_1 _0727_ (.A(\u_core.t_ref[2] ),
    .B_N(\u_core.t_fb[2] ),
    .Y(_0203_));
 sg13g2_nor2b_1 _0728_ (.A(\u_core.t_ref[3] ),
    .B_N(\u_core.t_fb[3] ),
    .Y(_0204_));
 sg13g2_nor2b_1 _0729_ (.A(\u_core.t_fb[3] ),
    .B_N(\u_core.t_ref[3] ),
    .Y(_0205_));
 sg13g2_nand2b_1 _0730_ (.Y(_0206_),
    .B(\u_core.t_ref[3] ),
    .A_N(\u_core.t_fb[3] ));
 sg13g2_o21ai_1 _0731_ (.B1(_0206_),
    .Y(_0207_),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_nor2b_1 _0732_ (.A(\u_core.t_ref[1] ),
    .B_N(\u_core.t_fb[1] ),
    .Y(_0208_));
 sg13g2_nand2b_1 _0733_ (.Y(_0209_),
    .B(\u_core.t_ref[0] ),
    .A_N(\u_core.t_fb[0] ));
 sg13g2_nand2b_1 _0734_ (.Y(_0210_),
    .B(\u_core.t_ref[1] ),
    .A_N(\u_core.t_fb[1] ));
 sg13g2_a21oi_1 _0735_ (.A1(_0209_),
    .A2(_0210_),
    .Y(_0211_),
    .B1(_0208_));
 sg13g2_nor2b_1 _0736_ (.A(\u_core.t_fb[2] ),
    .B_N(\u_core.t_ref[2] ),
    .Y(_0212_));
 sg13g2_or4_1 _0737_ (.A(_0203_),
    .B(_0204_),
    .C(_0205_),
    .D(_0212_),
    .X(_0213_));
 sg13g2_o21ai_1 _0738_ (.B1(_0207_),
    .Y(_0214_),
    .A1(_0211_),
    .A2(_0213_));
 sg13g2_xnor2_1 _0739_ (.Y(_0215_),
    .A(_0202_),
    .B(_0214_));
 sg13g2_nand2_1 _0740_ (.Y(_0216_),
    .A(net37),
    .B(net156));
 sg13g2_o21ai_1 _0741_ (.B1(_0216_),
    .Y(_0018_),
    .A1(net156),
    .A2(_0215_));
 sg13g2_a21oi_1 _0742_ (.A1(_0202_),
    .A2(_0214_),
    .Y(_0217_),
    .B1(_0201_));
 sg13g2_nor2_1 _0743_ (.A(\u_core.t_fb[5] ),
    .B(_0153_),
    .Y(_0218_));
 sg13g2_xnor2_1 _0744_ (.Y(_0219_),
    .A(\u_core.t_fb[5] ),
    .B(\u_core.t_ref[5] ));
 sg13g2_xnor2_1 _0745_ (.Y(_0220_),
    .A(_0217_),
    .B(_0219_));
 sg13g2_mux2_1 _0746_ (.A0(net253),
    .A1(_0220_),
    .S(net146),
    .X(_0019_));
 sg13g2_nand2b_1 _0747_ (.Y(_0221_),
    .B(\u_core.t_fb[6] ),
    .A_N(\u_core.t_ref[6] ));
 sg13g2_xor2_1 _0748_ (.B(net314),
    .A(\u_core.t_fb[6] ),
    .X(_0222_));
 sg13g2_a221oi_1 _0749_ (.B2(_0214_),
    .C1(_0201_),
    .B1(_0202_),
    .A1(\u_core.t_fb[5] ),
    .Y(_0223_),
    .A2(_0153_));
 sg13g2_o21ai_1 _0750_ (.B1(_0222_),
    .Y(_0224_),
    .A1(_0218_),
    .A2(_0223_));
 sg13g2_or3_1 _0751_ (.A(_0218_),
    .B(_0222_),
    .C(_0223_),
    .X(_0225_));
 sg13g2_and2_1 _0752_ (.A(_0224_),
    .B(_0225_),
    .X(_0226_));
 sg13g2_mux2_1 _0753_ (.A0(net242),
    .A1(_0226_),
    .S(net146),
    .X(_0020_));
 sg13g2_nor2b_1 _0754_ (.A(\u_core.t_ref[7] ),
    .B_N(\u_core.t_fb[7] ),
    .Y(_0227_));
 sg13g2_xor2_1 _0755_ (.B(\u_core.t_ref[7] ),
    .A(\u_core.t_fb[7] ),
    .X(_0228_));
 sg13g2_nand3_1 _0756_ (.B(_0225_),
    .C(_0228_),
    .A(_0221_),
    .Y(_0229_));
 sg13g2_a21oi_1 _0757_ (.A1(_0221_),
    .A2(_0225_),
    .Y(_0230_),
    .B1(_0228_));
 sg13g2_nand3b_1 _0758_ (.B(net146),
    .C(_0229_),
    .Y(_0231_),
    .A_N(_0230_));
 sg13g2_o21ai_1 _0759_ (.B1(_0231_),
    .Y(_0021_),
    .A1(_0150_),
    .A2(_0000_));
 sg13g2_or2_1 _0760_ (.X(_0232_),
    .B(_0230_),
    .A(_0227_));
 sg13g2_nor2b_1 _0761_ (.A(\u_core.t_ref[8] ),
    .B_N(\u_core.t_fb[8] ),
    .Y(_0233_));
 sg13g2_xnor2_1 _0762_ (.Y(_0234_),
    .A(net231),
    .B(net235));
 sg13g2_o21ai_1 _0763_ (.B1(_0234_),
    .Y(_0235_),
    .A1(_0227_),
    .A2(_0230_));
 sg13g2_o21ai_1 _0764_ (.B1(_0000_),
    .Y(_0236_),
    .A1(_0232_),
    .A2(_0234_));
 sg13g2_nor2b_1 _0765_ (.A(_0236_),
    .B_N(_0235_),
    .Y(_0237_));
 sg13g2_a21o_1 _0766_ (.A2(net155),
    .A1(net240),
    .B1(_0237_),
    .X(_0022_));
 sg13g2_xor2_1 _0767_ (.B(net66),
    .A(net96),
    .X(_0238_));
 sg13g2_nand2b_1 _0768_ (.Y(_0239_),
    .B(_0235_),
    .A_N(_0233_));
 sg13g2_xnor2_1 _0769_ (.Y(_0240_),
    .A(_0238_),
    .B(_0239_));
 sg13g2_mux2_1 _0770_ (.A0(net260),
    .A1(_0240_),
    .S(net146),
    .X(_0023_));
 sg13g2_nor2b_1 _0771_ (.A(\u_core.t_ref[10] ),
    .B_N(\u_core.t_fb[10] ),
    .Y(_0241_));
 sg13g2_xnor2_1 _0772_ (.Y(_0242_),
    .A(\u_core.t_fb[10] ),
    .B(\u_core.t_ref[10] ));
 sg13g2_inv_1 _0773_ (.Y(_0243_),
    .A(_0242_));
 sg13g2_a21oi_1 _0774_ (.A1(\u_core.t_fb[9] ),
    .A2(_0155_),
    .Y(_0244_),
    .B1(_0233_));
 sg13g2_a22oi_1 _0775_ (.Y(_0245_),
    .B1(_0235_),
    .B2(_0244_),
    .A2(\u_core.t_ref[9] ),
    .A1(_0154_));
 sg13g2_xnor2_1 _0776_ (.Y(_0246_),
    .A(_0243_),
    .B(_0245_));
 sg13g2_mux2_1 _0777_ (.A0(net305),
    .A1(_0246_),
    .S(net146),
    .X(_0024_));
 sg13g2_nor2b_1 _0778_ (.A(net238),
    .B_N(\u_core.t_fb[11] ),
    .Y(_0247_));
 sg13g2_nand2b_1 _0779_ (.Y(_0248_),
    .B(\u_core.t_ref[11] ),
    .A_N(net220));
 sg13g2_nand2b_1 _0780_ (.Y(_0249_),
    .B(_0248_),
    .A_N(_0247_));
 sg13g2_a21oi_1 _0781_ (.A1(_0242_),
    .A2(_0245_),
    .Y(_0250_),
    .B1(_0241_));
 sg13g2_xnor2_1 _0782_ (.Y(_0251_),
    .A(_0249_),
    .B(_0250_));
 sg13g2_nand2_1 _0783_ (.Y(_0252_),
    .A(net224),
    .B(net155));
 sg13g2_o21ai_1 _0784_ (.B1(net225),
    .Y(_0025_),
    .A1(net155),
    .A2(_0251_));
 sg13g2_nor2_1 _0785_ (.A(_0243_),
    .B(_0249_),
    .Y(_0253_));
 sg13g2_a221oi_1 _0786_ (.B2(_0245_),
    .C1(_0247_),
    .B1(_0253_),
    .A1(_0241_),
    .Y(_0254_),
    .A2(_0248_));
 sg13g2_nand2b_1 _0787_ (.Y(_0255_),
    .B(\u_core.t_fb[12] ),
    .A_N(\u_core.t_ref[12] ));
 sg13g2_xor2_1 _0788_ (.B(net269),
    .A(\u_core.t_fb[12] ),
    .X(_0256_));
 sg13g2_a21oi_1 _0789_ (.A1(_0254_),
    .A2(_0256_),
    .Y(_0257_),
    .B1(net155));
 sg13g2_o21ai_1 _0790_ (.B1(_0257_),
    .Y(_0258_),
    .A1(_0254_),
    .A2(_0256_));
 sg13g2_o21ai_1 _0791_ (.B1(_0258_),
    .Y(_0026_),
    .A1(_0148_),
    .A2(net146));
 sg13g2_xor2_1 _0792_ (.B(net91),
    .A(\u_core.t_fb[13] ),
    .X(_0259_));
 sg13g2_o21ai_1 _0793_ (.B1(_0255_),
    .Y(_0260_),
    .A1(_0254_),
    .A2(_0256_));
 sg13g2_xor2_1 _0794_ (.B(_0260_),
    .A(_0259_),
    .X(_0261_));
 sg13g2_nand2_1 _0795_ (.Y(_0262_),
    .A(net131),
    .B(net155));
 sg13g2_o21ai_1 _0796_ (.B1(net132),
    .Y(_0027_),
    .A1(net155),
    .A2(_0261_));
 sg13g2_nor2b_1 _0797_ (.A(net249),
    .B_N(net234),
    .Y(_0263_));
 sg13g2_nand2b_1 _0798_ (.Y(_0264_),
    .B(net249),
    .A_N(net234));
 sg13g2_nand2b_1 _0799_ (.Y(_0265_),
    .B(_0264_),
    .A_N(_0263_));
 sg13g2_or2_1 _0800_ (.X(_0266_),
    .B(_0259_),
    .A(_0256_));
 sg13g2_a21oi_1 _0801_ (.A1(_0156_),
    .A2(\u_core.t_ref[13] ),
    .Y(_0267_),
    .B1(_0255_));
 sg13g2_a21oi_1 _0802_ (.A1(\u_core.t_fb[13] ),
    .A2(_0157_),
    .Y(_0268_),
    .B1(_0267_));
 sg13g2_o21ai_1 _0803_ (.B1(_0268_),
    .Y(_0269_),
    .A1(_0254_),
    .A2(_0266_));
 sg13g2_xnor2_1 _0804_ (.Y(_0270_),
    .A(_0265_),
    .B(_0269_));
 sg13g2_mux2_1 _0805_ (.A0(net307),
    .A1(_0270_),
    .S(net146),
    .X(_0028_));
 sg13g2_a21oi_1 _0806_ (.A1(_0264_),
    .A2(_0269_),
    .Y(_0271_),
    .B1(_0263_));
 sg13g2_xor2_1 _0807_ (.B(net221),
    .A(net265),
    .X(_0272_));
 sg13g2_xnor2_1 _0808_ (.Y(_0273_),
    .A(_0271_),
    .B(_0272_));
 sg13g2_nand2_1 _0809_ (.Y(_0274_),
    .A(net175),
    .B(net155));
 sg13g2_o21ai_1 _0810_ (.B1(_0274_),
    .Y(_0029_),
    .A1(net155),
    .A2(_0273_));
 sg13g2_nor2_1 _0811_ (.A(net107),
    .B(_0185_),
    .Y(_0275_));
 sg13g2_mux2_1 _0812_ (.A0(net116),
    .A1(net42),
    .S(net154),
    .X(_0030_));
 sg13g2_mux2_1 _0813_ (.A0(net245),
    .A1(\u_core.beat_cnt[1] ),
    .S(net154),
    .X(_0031_));
 sg13g2_nor2_1 _0814_ (.A(net111),
    .B(net153),
    .Y(_0276_));
 sg13g2_a21oi_1 _0815_ (.A1(_0158_),
    .A2(net153),
    .Y(_0032_),
    .B1(_0276_));
 sg13g2_mux2_1 _0816_ (.A0(net304),
    .A1(net54),
    .S(net153),
    .X(_0033_));
 sg13g2_mux2_1 _0817_ (.A0(net292),
    .A1(net280),
    .S(net153),
    .X(_0034_));
 sg13g2_nor2_1 _0818_ (.A(net256),
    .B(net153),
    .Y(_0277_));
 sg13g2_a21oi_1 _0819_ (.A1(_0159_),
    .A2(net153),
    .Y(_0035_),
    .B1(_0277_));
 sg13g2_mux2_1 _0820_ (.A0(net289),
    .A1(net52),
    .S(net153),
    .X(_0036_));
 sg13g2_mux2_1 _0821_ (.A0(net277),
    .A1(\u_core.beat_cnt[7] ),
    .S(net153),
    .X(_0037_));
 sg13g2_nor2_1 _0822_ (.A(net235),
    .B(net151),
    .Y(_0278_));
 sg13g2_a21oi_1 _0823_ (.A1(_0160_),
    .A2(net152),
    .Y(_0038_),
    .B1(_0278_));
 sg13g2_nand2_1 _0824_ (.Y(_0279_),
    .A(net35),
    .B(net151));
 sg13g2_o21ai_1 _0825_ (.B1(_0279_),
    .Y(_0039_),
    .A1(_0155_),
    .A2(net151));
 sg13g2_mux2_1 _0826_ (.A0(net284),
    .A1(net46),
    .S(net152),
    .X(_0040_));
 sg13g2_mux2_1 _0827_ (.A0(net238),
    .A1(net69),
    .S(net151),
    .X(_0041_));
 sg13g2_mux2_1 _0828_ (.A0(net269),
    .A1(net59),
    .S(net151),
    .X(_0042_));
 sg13g2_nand2_1 _0829_ (.Y(_0280_),
    .A(net85),
    .B(net151));
 sg13g2_o21ai_1 _0830_ (.B1(_0280_),
    .Y(_0043_),
    .A1(_0157_),
    .A2(net151));
 sg13g2_mux2_1 _0831_ (.A0(net249),
    .A1(net61),
    .S(net151),
    .X(_0044_));
 sg13g2_mux2_1 _0832_ (.A0(net221),
    .A1(net43),
    .S(net152),
    .X(_0045_));
 sg13g2_mux2_1 _0833_ (.A0(fb_samp),
    .A1(net74),
    .S(_0182_),
    .X(_0046_));
 sg13g2_nand2_1 _0834_ (.Y(_0281_),
    .A(_0181_),
    .B(uo_out[2]));
 sg13g2_nor2_1 _0835_ (.A(net57),
    .B(_0281_),
    .Y(_0282_));
 sg13g2_mux2_1 _0836_ (.A0(net135),
    .A1(net42),
    .S(net150),
    .X(_0047_));
 sg13g2_mux2_1 _0837_ (.A0(net142),
    .A1(\u_core.beat_cnt[1] ),
    .S(net150),
    .X(_0048_));
 sg13g2_nor2_1 _0838_ (.A(net101),
    .B(net149),
    .Y(_0283_));
 sg13g2_a21oi_1 _0839_ (.A1(_0158_),
    .A2(net149),
    .Y(_0049_),
    .B1(_0283_));
 sg13g2_mux2_1 _0840_ (.A0(net295),
    .A1(net54),
    .S(net149),
    .X(_0050_));
 sg13g2_mux2_1 _0841_ (.A0(\u_core.t_fb[4] ),
    .A1(net280),
    .S(net149),
    .X(_0051_));
 sg13g2_nor2_1 _0842_ (.A(net255),
    .B(net149),
    .Y(_0284_));
 sg13g2_a21oi_1 _0843_ (.A1(_0159_),
    .A2(net149),
    .Y(_0052_),
    .B1(_0284_));
 sg13g2_mux2_1 _0844_ (.A0(net288),
    .A1(net52),
    .S(net149),
    .X(_0053_));
 sg13g2_mux2_1 _0845_ (.A0(net285),
    .A1(\u_core.beat_cnt[7] ),
    .S(net149),
    .X(_0054_));
 sg13g2_nor2_1 _0846_ (.A(net231),
    .B(net147),
    .Y(_0285_));
 sg13g2_a21oi_1 _0847_ (.A1(_0160_),
    .A2(net147),
    .Y(_0055_),
    .B1(_0285_));
 sg13g2_nand2_1 _0848_ (.Y(_0286_),
    .A(net35),
    .B(net148));
 sg13g2_o21ai_1 _0849_ (.B1(_0286_),
    .Y(_0056_),
    .A1(_0154_),
    .A2(net148));
 sg13g2_mux2_1 _0850_ (.A0(net287),
    .A1(net46),
    .S(net147),
    .X(_0057_));
 sg13g2_mux2_1 _0851_ (.A0(net220),
    .A1(net69),
    .S(net147),
    .X(_0058_));
 sg13g2_mux2_1 _0852_ (.A0(net296),
    .A1(net59),
    .S(net147),
    .X(_0059_));
 sg13g2_nand2_1 _0853_ (.Y(_0287_),
    .A(net85),
    .B(net147));
 sg13g2_o21ai_1 _0854_ (.B1(_0287_),
    .Y(_0060_),
    .A1(_0156_),
    .A2(net147));
 sg13g2_mux2_1 _0855_ (.A0(net234),
    .A1(net61),
    .S(net147),
    .X(_0061_));
 sg13g2_mux2_1 _0856_ (.A0(net265),
    .A1(net43),
    .S(net148),
    .X(_0062_));
 sg13g2_mux2_1 _0857_ (.A0(ref_samp),
    .A1(net125),
    .S(_0182_),
    .X(_0063_));
 sg13g2_o21ai_1 _0858_ (.B1(_0281_),
    .Y(_0064_),
    .A1(_0142_),
    .A2(_0182_));
 sg13g2_o21ai_1 _0859_ (.B1(net156),
    .Y(_0288_),
    .A1(net276),
    .A2(net154));
 sg13g2_inv_1 _0860_ (.Y(_0065_),
    .A(_0288_));
 sg13g2_nand2_1 _0861_ (.Y(_0289_),
    .A(net211),
    .B(\ctrl[8] ));
 sg13g2_xnor2_1 _0862_ (.Y(_0066_),
    .A(net33),
    .B(_0289_));
 sg13g2_nor2_1 _0863_ (.A(net212),
    .B(net134),
    .Y(_0290_));
 sg13g2_and2_1 _0864_ (.A(net33),
    .B(net67),
    .X(_0291_));
 sg13g2_and2_1 _0865_ (.A(\nco_phase_acc[1] ),
    .B(\ctrl[9] ),
    .X(_0292_));
 sg13g2_xor2_1 _0866_ (.B(net128),
    .A(net134),
    .X(_0293_));
 sg13g2_xnor2_1 _0867_ (.Y(_0294_),
    .A(_0291_),
    .B(_0293_));
 sg13g2_a21oi_1 _0868_ (.A1(net212),
    .A2(_0294_),
    .Y(_0067_),
    .B1(_0290_));
 sg13g2_nor2_1 _0869_ (.A(net212),
    .B(net117),
    .Y(_0295_));
 sg13g2_a21oi_1 _0870_ (.A1(_0291_),
    .A2(_0293_),
    .Y(_0296_),
    .B1(_0292_));
 sg13g2_nand2_1 _0871_ (.Y(_0297_),
    .A(\nco_phase_acc[2] ),
    .B(\ctrl[10] ));
 sg13g2_nor2_1 _0872_ (.A(\nco_phase_acc[2] ),
    .B(\ctrl[10] ),
    .Y(_0298_));
 sg13g2_xnor2_1 _0873_ (.Y(_0299_),
    .A(net117),
    .B(net102));
 sg13g2_xnor2_1 _0874_ (.Y(_0300_),
    .A(_0296_),
    .B(_0299_));
 sg13g2_a21oi_1 _0875_ (.A1(net212),
    .A2(_0300_),
    .Y(_0068_),
    .B1(_0295_));
 sg13g2_o21ai_1 _0876_ (.B1(_0297_),
    .Y(_0301_),
    .A1(_0296_),
    .A2(_0298_));
 sg13g2_and2_1 _0877_ (.A(\nco_phase_acc[3] ),
    .B(net48),
    .X(_0302_));
 sg13g2_or2_1 _0878_ (.X(_0303_),
    .B(net48),
    .A(\nco_phase_acc[3] ));
 sg13g2_nand2b_1 _0879_ (.Y(_0304_),
    .B(_0303_),
    .A_N(_0302_));
 sg13g2_xnor2_1 _0880_ (.Y(_0305_),
    .A(_0301_),
    .B(_0304_));
 sg13g2_mux2_1 _0881_ (.A0(net229),
    .A1(_0305_),
    .S(net211),
    .X(_0069_));
 sg13g2_nand2_1 _0882_ (.Y(_0306_),
    .A(\nco_phase_acc[4] ),
    .B(net104));
 sg13g2_xnor2_1 _0883_ (.Y(_0307_),
    .A(net216),
    .B(net104));
 sg13g2_a21oi_2 _0884_ (.B1(_0302_),
    .Y(_0308_),
    .A2(_0303_),
    .A1(_0301_));
 sg13g2_xnor2_1 _0885_ (.Y(_0309_),
    .A(_0307_),
    .B(_0308_));
 sg13g2_nor2_1 _0886_ (.A(net212),
    .B(net216),
    .Y(_0310_));
 sg13g2_a21oi_1 _0887_ (.A1(net211),
    .A2(_0309_),
    .Y(_0070_),
    .B1(_0310_));
 sg13g2_nor2_1 _0888_ (.A(net213),
    .B(net109),
    .Y(_0311_));
 sg13g2_or2_1 _0889_ (.X(_0312_),
    .B(\ctrl[13] ),
    .A(\nco_phase_acc[5] ));
 sg13g2_xor2_1 _0890_ (.B(net83),
    .A(net109),
    .X(_0313_));
 sg13g2_o21ai_1 _0891_ (.B1(_0306_),
    .Y(_0314_),
    .A1(_0307_),
    .A2(_0308_));
 sg13g2_xnor2_1 _0892_ (.Y(_0315_),
    .A(_0313_),
    .B(_0314_));
 sg13g2_a21oi_1 _0893_ (.A1(net214),
    .A2(_0315_),
    .Y(_0071_),
    .B1(_0311_));
 sg13g2_nand2_1 _0894_ (.Y(_0316_),
    .A(\nco_phase_acc[6] ),
    .B(net93));
 sg13g2_xor2_1 _0895_ (.B(net93),
    .A(net222),
    .X(_0317_));
 sg13g2_a22oi_1 _0896_ (.Y(_0318_),
    .B1(\nco_phase_acc[5] ),
    .B2(\ctrl[13] ),
    .A2(\ctrl[12] ),
    .A1(\nco_phase_acc[4] ));
 sg13g2_o21ai_1 _0897_ (.B1(_0318_),
    .Y(_0319_),
    .A1(_0307_),
    .A2(_0308_));
 sg13g2_nand3_1 _0898_ (.B(_0317_),
    .C(_0319_),
    .A(_0312_),
    .Y(_0320_));
 sg13g2_a21o_1 _0899_ (.A2(_0319_),
    .A1(_0312_),
    .B1(_0317_),
    .X(_0321_));
 sg13g2_nand3_1 _0900_ (.B(_0320_),
    .C(_0321_),
    .A(net213),
    .Y(_0322_));
 sg13g2_o21ai_1 _0901_ (.B1(_0322_),
    .Y(_0072_),
    .A1(net213),
    .A2(_0167_));
 sg13g2_nand2_1 _0902_ (.Y(_0323_),
    .A(\nco_phase_acc[7] ),
    .B(\ctrl[15] ));
 sg13g2_xnor2_1 _0903_ (.Y(_0324_),
    .A(net119),
    .B(\ctrl[15] ));
 sg13g2_a21o_1 _0904_ (.A2(_0320_),
    .A1(_0316_),
    .B1(_0324_),
    .X(_0325_));
 sg13g2_nand3_1 _0905_ (.B(_0320_),
    .C(_0324_),
    .A(_0316_),
    .Y(_0326_));
 sg13g2_a21oi_1 _0906_ (.A1(_0325_),
    .A2(_0326_),
    .Y(_0327_),
    .B1(net182));
 sg13g2_a21oi_1 _0907_ (.A1(net182),
    .A2(_0169_),
    .Y(_0073_),
    .B1(_0327_));
 sg13g2_nand2_1 _0908_ (.Y(_0328_),
    .A(_0323_),
    .B(_0325_));
 sg13g2_nand2_1 _0909_ (.Y(_0329_),
    .A(\nco_phase_acc[8] ),
    .B(\ctrl[16] ));
 sg13g2_xor2_1 _0910_ (.B(net140),
    .A(net297),
    .X(_0330_));
 sg13g2_nand2_1 _0911_ (.Y(_0331_),
    .A(_0328_),
    .B(_0330_));
 sg13g2_o21ai_1 _0912_ (.B1(net210),
    .Y(_0332_),
    .A1(_0328_),
    .A2(_0330_));
 sg13g2_nor2b_1 _0913_ (.A(_0332_),
    .B_N(_0331_),
    .Y(_0333_));
 sg13g2_a21o_1 _0914_ (.A2(net297),
    .A1(net182),
    .B1(_0333_),
    .X(_0074_));
 sg13g2_nor2_1 _0915_ (.A(net81),
    .B(net70),
    .Y(_0334_));
 sg13g2_nand2_1 _0916_ (.Y(_0335_),
    .A(net81),
    .B(net70));
 sg13g2_nor2b_1 _0917_ (.A(_0334_),
    .B_N(_0335_),
    .Y(_0336_));
 sg13g2_nand2_1 _0918_ (.Y(_0337_),
    .A(_0329_),
    .B(_0331_));
 sg13g2_xnor2_1 _0919_ (.Y(_0338_),
    .A(_0336_),
    .B(_0337_));
 sg13g2_nor2_1 _0920_ (.A(net210),
    .B(net81),
    .Y(_0339_));
 sg13g2_a21oi_1 _0921_ (.A1(net210),
    .A2(_0338_),
    .Y(_0075_),
    .B1(_0339_));
 sg13g2_nor2_1 _0922_ (.A(net209),
    .B(net127),
    .Y(_0340_));
 sg13g2_nand2_1 _0923_ (.Y(_0341_),
    .A(\nco_phase_acc[10] ),
    .B(net95));
 sg13g2_xnor2_1 _0924_ (.Y(_0342_),
    .A(net127),
    .B(net95));
 sg13g2_o21ai_1 _0925_ (.B1(_0335_),
    .Y(_0343_),
    .A1(_0329_),
    .A2(_0334_));
 sg13g2_nand2_1 _0926_ (.Y(_0344_),
    .A(_0330_),
    .B(_0336_));
 sg13g2_inv_1 _0927_ (.Y(_0345_),
    .A(_0344_));
 sg13g2_a21oi_1 _0928_ (.A1(_0328_),
    .A2(_0345_),
    .Y(_0346_),
    .B1(_0343_));
 sg13g2_xnor2_1 _0929_ (.Y(_0347_),
    .A(_0342_),
    .B(_0346_));
 sg13g2_a21oi_1 _0930_ (.A1(net209),
    .A2(_0347_),
    .Y(_0076_),
    .B1(_0340_));
 sg13g2_o21ai_1 _0931_ (.B1(_0341_),
    .Y(_0348_),
    .A1(_0342_),
    .A2(_0346_));
 sg13g2_xor2_1 _0932_ (.B(\ctrl[19] ),
    .A(net123),
    .X(_0349_));
 sg13g2_xnor2_1 _0933_ (.Y(_0350_),
    .A(_0348_),
    .B(_0349_));
 sg13g2_nor2_1 _0934_ (.A(net209),
    .B(net123),
    .Y(_0351_));
 sg13g2_a21oi_1 _0935_ (.A1(net209),
    .A2(_0350_),
    .Y(_0077_),
    .B1(_0351_));
 sg13g2_nor2_1 _0936_ (.A(net209),
    .B(net130),
    .Y(_0352_));
 sg13g2_nor2b_1 _0937_ (.A(_0342_),
    .B_N(_0349_),
    .Y(_0353_));
 sg13g2_nand2_1 _0938_ (.Y(_0354_),
    .A(_0345_),
    .B(_0353_));
 sg13g2_a21o_1 _0939_ (.A2(_0325_),
    .A1(_0323_),
    .B1(_0354_),
    .X(_0355_));
 sg13g2_a21oi_1 _0940_ (.A1(_0174_),
    .A2(_0175_),
    .Y(_0356_),
    .B1(_0341_));
 sg13g2_a221oi_1 _0941_ (.B2(_0353_),
    .C1(_0356_),
    .B1(_0343_),
    .A1(\nco_phase_acc[11] ),
    .Y(_0357_),
    .A2(\ctrl[19] ));
 sg13g2_and2_1 _0942_ (.A(_0355_),
    .B(_0357_),
    .X(_0358_));
 sg13g2_nand2_1 _0943_ (.Y(_0359_),
    .A(\nco_phase_acc[12] ),
    .B(net97));
 sg13g2_xnor2_1 _0944_ (.Y(_0360_),
    .A(net130),
    .B(net97));
 sg13g2_xnor2_1 _0945_ (.Y(_0361_),
    .A(_0358_),
    .B(_0360_));
 sg13g2_a21oi_1 _0946_ (.A1(net209),
    .A2(_0361_),
    .Y(_0078_),
    .B1(_0352_));
 sg13g2_nor2_1 _0947_ (.A(net99),
    .B(net89),
    .Y(_0362_));
 sg13g2_nand2_1 _0948_ (.Y(_0363_),
    .A(net99),
    .B(net89));
 sg13g2_nand2b_1 _0949_ (.Y(_0364_),
    .B(_0363_),
    .A_N(_0362_));
 sg13g2_o21ai_1 _0950_ (.B1(_0359_),
    .Y(_0365_),
    .A1(_0358_),
    .A2(_0360_));
 sg13g2_xor2_1 _0951_ (.B(_0365_),
    .A(_0364_),
    .X(_0366_));
 sg13g2_nor2_1 _0952_ (.A(net211),
    .B(net99),
    .Y(_0367_));
 sg13g2_a21oi_1 _0953_ (.A1(net209),
    .A2(_0366_),
    .Y(_0079_),
    .B1(_0367_));
 sg13g2_nand2_1 _0954_ (.Y(_0368_),
    .A(net112),
    .B(net121));
 sg13g2_xor2_1 _0955_ (.B(\ctrl[22] ),
    .A(\nco_phase_acc[14] ),
    .X(_0369_));
 sg13g2_or2_1 _0956_ (.X(_0370_),
    .B(_0364_),
    .A(_0360_));
 sg13g2_a21oi_1 _0957_ (.A1(_0355_),
    .A2(_0357_),
    .Y(_0371_),
    .B1(_0370_));
 sg13g2_o21ai_1 _0958_ (.B1(_0363_),
    .Y(_0372_),
    .A1(_0359_),
    .A2(_0362_));
 sg13g2_o21ai_1 _0959_ (.B1(_0369_),
    .Y(_0373_),
    .A1(_0371_),
    .A2(_0372_));
 sg13g2_or3_1 _0960_ (.A(_0369_),
    .B(_0371_),
    .C(_0372_),
    .X(_0374_));
 sg13g2_nand3_1 _0961_ (.B(_0373_),
    .C(_0374_),
    .A(net211),
    .Y(_0375_));
 sg13g2_o21ai_1 _0962_ (.B1(_0375_),
    .Y(_0080_),
    .A1(net211),
    .A2(_0178_));
 sg13g2_nor2_1 _0963_ (.A(\nco_phase_acc[15] ),
    .B(\ctrl[23] ),
    .Y(_0376_));
 sg13g2_xor2_1 _0964_ (.B(\ctrl[23] ),
    .A(net247),
    .X(_0377_));
 sg13g2_nand2_1 _0965_ (.Y(_0378_),
    .A(_0368_),
    .B(_0373_));
 sg13g2_xnor2_1 _0966_ (.Y(_0379_),
    .A(_0377_),
    .B(_0378_));
 sg13g2_nor2_1 _0967_ (.A(net211),
    .B(net247),
    .Y(_0380_));
 sg13g2_a21oi_1 _0968_ (.A1(net211),
    .A2(_0379_),
    .Y(_0081_),
    .B1(_0380_));
 sg13g2_and2_1 _0969_ (.A(_0369_),
    .B(_0377_),
    .X(_0381_));
 sg13g2_nand2b_1 _0970_ (.Y(_0382_),
    .B(_0381_),
    .A_N(_0370_));
 sg13g2_a21oi_1 _0971_ (.A1(_0355_),
    .A2(_0357_),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_nor2_1 _0972_ (.A(_0368_),
    .B(_0376_),
    .Y(_0384_));
 sg13g2_a221oi_1 _0973_ (.B2(_0381_),
    .C1(_0384_),
    .B1(_0372_),
    .A1(net309),
    .Y(_0385_),
    .A2(\ctrl[23] ));
 sg13g2_inv_1 _0974_ (.Y(_0386_),
    .A(_0385_));
 sg13g2_nand2b_1 _0975_ (.Y(_0387_),
    .B(net310),
    .A_N(_0383_));
 sg13g2_o21ai_1 _0976_ (.B1(net79),
    .Y(_0388_),
    .A1(_0141_),
    .A2(_0387_));
 sg13g2_nor3_1 _0977_ (.A(net79),
    .B(_0383_),
    .C(_0386_),
    .Y(_0389_));
 sg13g2_or2_1 _0978_ (.X(_0390_),
    .B(_0387_),
    .A(net79));
 sg13g2_o21ai_1 _0979_ (.B1(net80),
    .Y(_0082_),
    .A1(net182),
    .A2(_0390_));
 sg13g2_nand3_1 _0980_ (.B(net92),
    .C(_0390_),
    .A(net213),
    .Y(_0391_));
 sg13g2_a21o_1 _0981_ (.A2(_0390_),
    .A1(net213),
    .B1(net92),
    .X(_0392_));
 sg13g2_and2_1 _0982_ (.A(_0391_),
    .B(_0392_),
    .X(_0083_));
 sg13g2_nand3_1 _0983_ (.B(net92),
    .C(net31),
    .A(net213),
    .Y(_0393_));
 sg13g2_or2_1 _0984_ (.X(_0394_),
    .B(_0393_),
    .A(_0389_));
 sg13g2_xnor2_1 _0985_ (.Y(_0084_),
    .A(net31),
    .B(_0391_));
 sg13g2_nor3_2 _0986_ (.A(_0180_),
    .B(_0389_),
    .C(_0393_),
    .Y(_0395_));
 sg13g2_a21oi_1 _0987_ (.A1(_0180_),
    .A2(_0394_),
    .Y(_0085_),
    .B1(net77));
 sg13g2_xor2_1 _0988_ (.B(_0395_),
    .A(net39),
    .X(_0086_));
 sg13g2_a21oi_1 _0989_ (.A1(net39),
    .A2(net77),
    .Y(_0396_),
    .B1(net64));
 sg13g2_nand3_1 _0990_ (.B(net64),
    .C(_0395_),
    .A(net39),
    .Y(_0397_));
 sg13g2_nor2b_1 _0991_ (.A(_0396_),
    .B_N(_0397_),
    .Y(_0087_));
 sg13g2_nand4_1 _0992_ (.B(net64),
    .C(net29),
    .A(net39),
    .Y(_0398_),
    .D(_0395_));
 sg13g2_xnor2_1 _0993_ (.Y(_0088_),
    .A(net29),
    .B(_0397_));
 sg13g2_xnor2_1 _0994_ (.Y(_0089_),
    .A(net22),
    .B(net65));
 sg13g2_xor2_1 _0995_ (.B(net236),
    .A(net176),
    .X(_0399_));
 sg13g2_nand2_1 _0996_ (.Y(_0400_),
    .A(net176),
    .B(\u_lf.i_acc[26] ));
 sg13g2_nor2_1 _0997_ (.A(net176),
    .B(\u_lf.i_acc[26] ),
    .Y(_0401_));
 sg13g2_xor2_1 _0998_ (.B(net252),
    .A(net176),
    .X(_0402_));
 sg13g2_nand2_1 _0999_ (.Y(_0403_),
    .A(net181),
    .B(\u_lf.i_acc[25] ));
 sg13g2_nand2_1 _1000_ (.Y(_0404_),
    .A(net181),
    .B(net267));
 sg13g2_o21ai_1 _1001_ (.B1(net181),
    .Y(_0405_),
    .A1(\u_lf.i_acc[25] ),
    .A2(\u_lf.i_acc[24] ));
 sg13g2_nand2_1 _1002_ (.Y(_0406_),
    .A(_0403_),
    .B(_0404_));
 sg13g2_and2_1 _1003_ (.A(net178),
    .B(net87),
    .X(_0407_));
 sg13g2_o21ai_1 _1004_ (.B1(net178),
    .Y(_0408_),
    .A1(\u_lf.i_acc[17] ),
    .A2(\u_lf.i_acc[16] ));
 sg13g2_o21ai_1 _1005_ (.B1(net179),
    .Y(_0409_),
    .A1(\u_lf.i_acc[19] ),
    .A2(\u_lf.i_acc[18] ));
 sg13g2_nand2_1 _1006_ (.Y(_0410_),
    .A(_0408_),
    .B(_0409_));
 sg13g2_nand2_1 _1007_ (.Y(_0411_),
    .A(net177),
    .B(\u_lf.i_acc[22] ));
 sg13g2_nand2_1 _1008_ (.Y(_0412_),
    .A(net178),
    .B(\u_lf.i_acc[20] ));
 sg13g2_o21ai_1 _1009_ (.B1(net179),
    .Y(_0413_),
    .A1(\u_lf.i_acc[21] ),
    .A2(\u_lf.i_acc[20] ));
 sg13g2_inv_1 _1010_ (.Y(_0414_),
    .A(_0413_));
 sg13g2_and2_1 _1011_ (.A(_0411_),
    .B(_0413_),
    .X(_0415_));
 sg13g2_a21oi_1 _1012_ (.A1(net176),
    .A2(\u_lf.i_acc[23] ),
    .Y(_0416_),
    .B1(_0410_));
 sg13g2_and2_1 _1013_ (.A(_0415_),
    .B(_0416_),
    .X(_0417_));
 sg13g2_nand2_1 _1014_ (.Y(_0418_),
    .A(net171),
    .B(net313));
 sg13g2_nand2_1 _1015_ (.Y(_0419_),
    .A(net172),
    .B(net106));
 sg13g2_nand2_1 _1016_ (.Y(_0420_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_and2_1 _1017_ (.A(net171),
    .B(net259),
    .X(_0421_));
 sg13g2_o21ai_1 _1018_ (.B1(net171),
    .Y(_0422_),
    .A1(\u_lf.i_acc[15] ),
    .A2(\u_lf.i_acc[14] ));
 sg13g2_nand3_1 _1019_ (.B(_0419_),
    .C(_0422_),
    .A(_0418_),
    .Y(_0423_));
 sg13g2_xnor2_1 _1020_ (.Y(_0424_),
    .A(net172),
    .B(net106));
 sg13g2_or2_1 _1021_ (.X(_0425_),
    .B(net259),
    .A(net171));
 sg13g2_xnor2_1 _1022_ (.Y(_0426_),
    .A(net171),
    .B(net259));
 sg13g2_nor2_1 _1023_ (.A(_0424_),
    .B(_0426_),
    .Y(_0427_));
 sg13g2_xor2_1 _1024_ (.B(net262),
    .A(net171),
    .X(_0428_));
 sg13g2_xor2_1 _1025_ (.B(net266),
    .A(net171),
    .X(_0429_));
 sg13g2_nand3_1 _1026_ (.B(_0428_),
    .C(_0429_),
    .A(_0427_),
    .Y(_0430_));
 sg13g2_inv_1 _1027_ (.Y(_0431_),
    .A(_0430_));
 sg13g2_nor2_1 _1028_ (.A(net173),
    .B(\u_lf.i_acc[11] ),
    .Y(_0432_));
 sg13g2_a22oi_1 _1029_ (.Y(_0433_),
    .B1(\u_lf.i_acc[10] ),
    .B2(\phase_err_beat[14] ),
    .A2(\u_lf.i_acc[11] ),
    .A1(net173));
 sg13g2_xnor2_1 _1030_ (.Y(_0434_),
    .A(net172),
    .B(net279));
 sg13g2_xnor2_1 _1031_ (.Y(_0435_),
    .A(\u_lf.i_acc[10] ),
    .B(\phase_err_beat[14] ));
 sg13g2_nor2_1 _1032_ (.A(_0434_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_a22oi_1 _1033_ (.Y(_0437_),
    .B1(\u_lf.i_acc[8] ),
    .B2(\phase_err_beat[12] ),
    .A2(\phase_err_beat[13] ),
    .A1(\u_lf.i_acc[9] ));
 sg13g2_or2_1 _1034_ (.X(_0438_),
    .B(\phase_err_beat[13] ),
    .A(\u_lf.i_acc[9] ));
 sg13g2_nand3b_1 _1035_ (.B(_0438_),
    .C(_0436_),
    .Y(_0439_),
    .A_N(_0437_));
 sg13g2_o21ai_1 _1036_ (.B1(_0439_),
    .Y(_0440_),
    .A1(_0432_),
    .A2(_0433_));
 sg13g2_a22oi_1 _1037_ (.Y(_0441_),
    .B1(\u_lf.i_acc[6] ),
    .B2(\phase_err_beat[10] ),
    .A2(\phase_err_beat[11] ),
    .A1(\u_lf.i_acc[7] ));
 sg13g2_nand2_1 _1038_ (.Y(_0442_),
    .A(\phase_err_beat[8] ),
    .B(\u_lf.i_acc[4] ));
 sg13g2_nand2_1 _1039_ (.Y(_0443_),
    .A(\phase_err_beat[9] ),
    .B(\u_lf.i_acc[5] ));
 sg13g2_and2_1 _1040_ (.A(_0442_),
    .B(_0443_),
    .X(_0444_));
 sg13g2_and2_1 _1041_ (.A(\phase_err_beat[6] ),
    .B(\u_lf.i_acc[2] ),
    .X(_0445_));
 sg13g2_nand2_1 _1042_ (.Y(_0446_),
    .A(\phase_err_beat[5] ),
    .B(\u_lf.i_acc[1] ));
 sg13g2_nand2_1 _1043_ (.Y(_0447_),
    .A(\phase_err_beat[4] ),
    .B(\u_lf.i_acc[0] ));
 sg13g2_nor2_1 _1044_ (.A(\phase_err_beat[5] ),
    .B(\u_lf.i_acc[1] ),
    .Y(_0448_));
 sg13g2_o21ai_1 _1045_ (.B1(_0446_),
    .Y(_0449_),
    .A1(_0447_),
    .A2(_0448_));
 sg13g2_or2_1 _1046_ (.X(_0450_),
    .B(\u_lf.i_acc[2] ),
    .A(\phase_err_beat[6] ));
 sg13g2_a221oi_1 _1047_ (.B2(_0450_),
    .C1(_0445_),
    .B1(_0449_),
    .A1(\phase_err_beat[7] ),
    .Y(_0451_),
    .A2(\u_lf.i_acc[3] ));
 sg13g2_or2_1 _1048_ (.X(_0452_),
    .B(\u_lf.i_acc[4] ),
    .A(\phase_err_beat[8] ));
 sg13g2_or2_1 _1049_ (.X(_0453_),
    .B(\phase_err_beat[10] ),
    .A(\u_lf.i_acc[6] ));
 sg13g2_nor2_1 _1050_ (.A(\phase_err_beat[9] ),
    .B(\u_lf.i_acc[5] ),
    .Y(_0454_));
 sg13g2_or2_1 _1051_ (.X(_0455_),
    .B(\phase_err_beat[12] ),
    .A(\u_lf.i_acc[8] ));
 sg13g2_or2_1 _1052_ (.X(_0456_),
    .B(\phase_err_beat[11] ),
    .A(\u_lf.i_acc[7] ));
 sg13g2_nor2b_1 _1053_ (.A(_0441_),
    .B_N(_0456_),
    .Y(_0457_));
 sg13g2_and3_1 _1054_ (.X(_0458_),
    .A(_0441_),
    .B(_0453_),
    .C(_0456_));
 sg13g2_a21oi_1 _1055_ (.A1(_0150_),
    .A2(_0151_),
    .Y(_0459_),
    .B1(_0454_));
 sg13g2_nand4_1 _1056_ (.B(_0452_),
    .C(_0458_),
    .A(_0444_),
    .Y(_0460_),
    .D(_0459_));
 sg13g2_o21ai_1 _1057_ (.B1(_0443_),
    .Y(_0461_),
    .A1(_0442_),
    .A2(_0454_));
 sg13g2_a21oi_1 _1058_ (.A1(_0458_),
    .A2(_0461_),
    .Y(_0462_),
    .B1(_0457_));
 sg13g2_o21ai_1 _1059_ (.B1(_0462_),
    .Y(_0463_),
    .A1(_0451_),
    .A2(_0460_));
 sg13g2_nand4_1 _1060_ (.B(_0437_),
    .C(_0438_),
    .A(_0436_),
    .Y(_0464_),
    .D(_0455_));
 sg13g2_nor2_1 _1061_ (.A(_0430_),
    .B(_0464_),
    .Y(_0465_));
 sg13g2_a221oi_1 _1062_ (.B2(_0465_),
    .C1(_0423_),
    .B1(_0463_),
    .A1(_0431_),
    .Y(_0466_),
    .A2(_0440_));
 sg13g2_xnor2_1 _1063_ (.Y(_0467_),
    .A(net178),
    .B(net264));
 sg13g2_xor2_1 _1064_ (.B(net230),
    .A(net178),
    .X(_0468_));
 sg13g2_xor2_1 _1065_ (.B(net87),
    .A(net178),
    .X(_0469_));
 sg13g2_xnor2_1 _1066_ (.Y(_0470_),
    .A(net178),
    .B(net72));
 sg13g2_inv_1 _1067_ (.Y(_0471_),
    .A(_0470_));
 sg13g2_nand3_1 _1068_ (.B(_0469_),
    .C(_0471_),
    .A(_0468_),
    .Y(_0472_));
 sg13g2_nor2_1 _1069_ (.A(_0467_),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_xnor2_1 _1070_ (.Y(_0474_),
    .A(net179),
    .B(net218));
 sg13g2_xnor2_1 _1071_ (.Y(_0475_),
    .A(net179),
    .B(net273));
 sg13g2_nor2_1 _1072_ (.A(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sg13g2_xor2_1 _1073_ (.B(net232),
    .A(net176),
    .X(_0477_));
 sg13g2_nor2_1 _1074_ (.A(net177),
    .B(\u_lf.i_acc[22] ),
    .Y(_0478_));
 sg13g2_xor2_1 _1075_ (.B(net283),
    .A(net176),
    .X(_0479_));
 sg13g2_nand4_1 _1076_ (.B(_0476_),
    .C(_0477_),
    .A(_0473_),
    .Y(_0480_),
    .D(_0479_));
 sg13g2_o21ai_1 _1077_ (.B1(_0417_),
    .Y(_0481_),
    .A1(_0466_),
    .A2(_0480_));
 sg13g2_o21ai_1 _1078_ (.B1(_0405_),
    .Y(_0482_),
    .A1(net181),
    .A2(\u_lf.i_acc[25] ));
 sg13g2_xnor2_1 _1079_ (.Y(_0483_),
    .A(net181),
    .B(\u_lf.i_acc[24] ));
 sg13g2_xor2_1 _1080_ (.B(net303),
    .A(net181),
    .X(_0484_));
 sg13g2_nor2b_1 _1081_ (.A(_0483_),
    .B_N(_0484_),
    .Y(_0485_));
 sg13g2_and2_1 _1082_ (.A(_0481_),
    .B(_0485_),
    .X(_0486_));
 sg13g2_o21ai_1 _1083_ (.B1(_0402_),
    .Y(_0487_),
    .A1(_0406_),
    .A2(_0486_));
 sg13g2_nand2_1 _1084_ (.Y(_0488_),
    .A(_0400_),
    .B(_0487_));
 sg13g2_xnor2_1 _1085_ (.Y(_0489_),
    .A(_0399_),
    .B(_0488_));
 sg13g2_nor2b_1 _1086_ (.A(_0466_),
    .B_N(_0473_),
    .Y(_0490_));
 sg13g2_o21ai_1 _1087_ (.B1(_0476_),
    .Y(_0491_),
    .A1(_0410_),
    .A2(_0490_));
 sg13g2_a21oi_1 _1088_ (.A1(_0415_),
    .A2(_0491_),
    .Y(_0492_),
    .B1(_0478_));
 sg13g2_xor2_1 _1089_ (.B(_0492_),
    .A(_0477_),
    .X(_0493_));
 sg13g2_or3_1 _1090_ (.A(_0402_),
    .B(_0406_),
    .C(_0486_),
    .X(_0494_));
 sg13g2_xor2_1 _1091_ (.B(_0483_),
    .A(_0481_),
    .X(_0495_));
 sg13g2_nand3_1 _1092_ (.B(\u_lf.i_acc[25] ),
    .C(\u_lf.i_acc[24] ),
    .A(net181),
    .Y(_0496_));
 sg13g2_a21oi_1 _1093_ (.A1(_0482_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(_0495_));
 sg13g2_nand3_1 _1094_ (.B(_0494_),
    .C(_0497_),
    .A(_0487_),
    .Y(_0498_));
 sg13g2_o21ai_1 _1095_ (.B1(net176),
    .Y(_0499_),
    .A1(\u_lf.i_acc[27] ),
    .A2(net252));
 sg13g2_nand2_1 _1096_ (.Y(_0500_),
    .A(_0405_),
    .B(_0499_));
 sg13g2_and3_1 _1097_ (.X(_0501_),
    .A(_0399_),
    .B(_0402_),
    .C(_0485_));
 sg13g2_a21oi_1 _1098_ (.A1(_0481_),
    .A2(_0501_),
    .Y(_0502_),
    .B1(_0500_));
 sg13g2_nand2_1 _1099_ (.Y(_0503_),
    .A(net177),
    .B(\u_lf.i_acc[28] ));
 sg13g2_xnor2_1 _1100_ (.Y(_0504_),
    .A(net177),
    .B(net257));
 sg13g2_xnor2_1 _1101_ (.Y(_0505_),
    .A(_0502_),
    .B(_0504_));
 sg13g2_nor3_1 _1102_ (.A(_0489_),
    .B(_0498_),
    .C(_0505_),
    .Y(_0506_));
 sg13g2_o21ai_1 _1103_ (.B1(_0503_),
    .Y(_0507_),
    .A1(_0502_),
    .A2(_0504_));
 sg13g2_xor2_1 _1104_ (.B(net177),
    .A(net138),
    .X(_0508_));
 sg13g2_o21ai_1 _1105_ (.B1(net160),
    .Y(_0509_),
    .A1(_0507_),
    .A2(_0508_));
 sg13g2_a221oi_1 _1106_ (.B2(_0508_),
    .C1(_0509_),
    .B1(_0507_),
    .A1(_0493_),
    .Y(_0510_),
    .A2(_0506_));
 sg13g2_a21oi_1 _1107_ (.A1(_0144_),
    .A2(net168),
    .Y(_0090_),
    .B1(net143));
 sg13g2_a21oi_1 _1108_ (.A1(_0145_),
    .A2(net168),
    .Y(_0091_),
    .B1(net143));
 sg13g2_a21oi_1 _1109_ (.A1(_0146_),
    .A2(net168),
    .Y(_0092_),
    .B1(net143));
 sg13g2_a21oi_1 _1110_ (.A1(_0147_),
    .A2(net168),
    .Y(_0093_),
    .B1(net143));
 sg13g2_a21oi_1 _1111_ (.A1(_0162_),
    .A2(net166),
    .Y(_0094_),
    .B1(net144));
 sg13g2_a21oi_1 _1112_ (.A1(_0161_),
    .A2(net166),
    .Y(_0095_),
    .B1(net144));
 sg13g2_a21oi_1 _1113_ (.A1(_0163_),
    .A2(net166),
    .Y(_0096_),
    .B1(net144));
 sg13g2_a21oi_1 _1114_ (.A1(_0164_),
    .A2(net169),
    .Y(_0097_),
    .B1(net144));
 sg13g2_a21oi_1 _1115_ (.A1(_0165_),
    .A2(net169),
    .Y(_0098_),
    .B1(net144));
 sg13g2_a21oi_1 _1116_ (.A1(_0166_),
    .A2(net169),
    .Y(_0099_),
    .B1(net145));
 sg13g2_a21oi_1 _1117_ (.A1(_0168_),
    .A2(net169),
    .Y(_0100_),
    .B1(net144));
 sg13g2_a21oi_1 _1118_ (.A1(_0170_),
    .A2(net170),
    .Y(_0101_),
    .B1(net145));
 sg13g2_a21oi_1 _1119_ (.A1(_0171_),
    .A2(net169),
    .Y(_0102_),
    .B1(net143));
 sg13g2_a21oi_1 _1120_ (.A1(_0172_),
    .A2(net169),
    .Y(_0103_),
    .B1(net143));
 sg13g2_a21oi_1 _1121_ (.A1(_0173_),
    .A2(net168),
    .Y(_0104_),
    .B1(net145));
 sg13g2_a21oi_1 _1122_ (.A1(_0175_),
    .A2(net168),
    .Y(_0105_),
    .B1(net143));
 sg13g2_a21oi_1 _1123_ (.A1(_0176_),
    .A2(net167),
    .Y(_0106_),
    .B1(net143));
 sg13g2_a21oi_1 _1124_ (.A1(_0177_),
    .A2(net166),
    .Y(_0107_),
    .B1(net144));
 sg13g2_a21oi_1 _1125_ (.A1(_0179_),
    .A2(net170),
    .Y(_0108_),
    .B1(net144));
 sg13g2_a21o_1 _1126_ (.A2(net170),
    .A1(net250),
    .B1(net145),
    .X(_0109_));
 sg13g2_o21ai_1 _1127_ (.B1(net156),
    .Y(_0511_),
    .A1(net263),
    .A2(net150));
 sg13g2_inv_1 _1128_ (.Y(_0110_),
    .A(_0511_));
 sg13g2_nand2_1 _1129_ (.Y(_0512_),
    .A(\phase_err_beat[10] ),
    .B(uo_out[0]));
 sg13g2_xnor2_1 _1130_ (.Y(_0111_),
    .A(net50),
    .B(_0512_));
 sg13g2_nand2_1 _1131_ (.Y(_0513_),
    .A(\phase_err_beat[11] ),
    .B(\u_lf.i_acc[1] ));
 sg13g2_xor2_1 _1132_ (.B(net301),
    .A(net224),
    .X(_0514_));
 sg13g2_a21oi_1 _1133_ (.A1(\phase_err_beat[10] ),
    .A2(net50),
    .Y(_0515_),
    .B1(_0514_));
 sg13g2_nand3_1 _1134_ (.B(net50),
    .C(_0514_),
    .A(\phase_err_beat[10] ),
    .Y(_0516_));
 sg13g2_nor2_1 _1135_ (.A(net168),
    .B(_0515_),
    .Y(_0517_));
 sg13g2_a22oi_1 _1136_ (.Y(_0518_),
    .B1(_0516_),
    .B2(_0517_),
    .A2(net168),
    .A1(net301));
 sg13g2_inv_1 _1137_ (.Y(_0112_),
    .A(net302));
 sg13g2_nand2_1 _1138_ (.Y(_0519_),
    .A(\phase_err_beat[12] ),
    .B(net114));
 sg13g2_xnor2_1 _1139_ (.Y(_0520_),
    .A(\phase_err_beat[12] ),
    .B(net114));
 sg13g2_nand3_1 _1140_ (.B(_0516_),
    .C(_0520_),
    .A(_0513_),
    .Y(_0521_));
 sg13g2_a21o_1 _1141_ (.A2(_0516_),
    .A1(_0513_),
    .B1(_0520_),
    .X(_0522_));
 sg13g2_a21oi_1 _1142_ (.A1(_0521_),
    .A2(_0522_),
    .Y(_0523_),
    .B1(net165));
 sg13g2_a21oi_1 _1143_ (.A1(_0152_),
    .A2(net165),
    .Y(_0113_),
    .B1(_0523_));
 sg13g2_nand2_1 _1144_ (.Y(_0524_),
    .A(net131),
    .B(net270));
 sg13g2_xnor2_1 _1145_ (.Y(_0525_),
    .A(net131),
    .B(net270));
 sg13g2_nand3_1 _1146_ (.B(_0522_),
    .C(_0525_),
    .A(_0519_),
    .Y(_0526_));
 sg13g2_a21o_1 _1147_ (.A2(_0522_),
    .A1(_0519_),
    .B1(_0525_),
    .X(_0527_));
 sg13g2_a21oi_1 _1148_ (.A1(_0526_),
    .A2(_0527_),
    .Y(_0528_),
    .B1(net165));
 sg13g2_a21oi_1 _1149_ (.A1(_0151_),
    .A2(net165),
    .Y(_0114_),
    .B1(_0528_));
 sg13g2_xnor2_1 _1150_ (.Y(_0529_),
    .A(\phase_err_beat[14] ),
    .B(net274));
 sg13g2_a21o_2 _1151_ (.A2(_0527_),
    .A1(_0524_),
    .B1(_0529_),
    .X(_0530_));
 sg13g2_inv_1 _1152_ (.Y(_0531_),
    .A(_0530_));
 sg13g2_nand3_1 _1153_ (.B(_0527_),
    .C(_0529_),
    .A(_0524_),
    .Y(_0532_));
 sg13g2_a21oi_1 _1154_ (.A1(_0530_),
    .A2(_0532_),
    .Y(_0533_),
    .B1(net166));
 sg13g2_a21oi_1 _1155_ (.A1(_0149_),
    .A2(net166),
    .Y(_0115_),
    .B1(_0533_));
 sg13g2_nor2_1 _1156_ (.A(net290),
    .B(net159),
    .Y(_0534_));
 sg13g2_nor2_1 _1157_ (.A(net175),
    .B(net290),
    .Y(_0535_));
 sg13g2_xnor2_1 _1158_ (.Y(_0536_),
    .A(net175),
    .B(net290));
 sg13g2_a21oi_1 _1159_ (.A1(\phase_err_beat[14] ),
    .A2(net274),
    .Y(_0537_),
    .B1(_0531_));
 sg13g2_xnor2_1 _1160_ (.Y(_0538_),
    .A(_0536_),
    .B(_0537_));
 sg13g2_a21oi_1 _1161_ (.A1(net159),
    .A2(_0538_),
    .Y(_0116_),
    .B1(_0534_));
 sg13g2_a22oi_1 _1162_ (.Y(_0539_),
    .B1(\u_lf.i_acc[4] ),
    .B2(\phase_err_beat[14] ),
    .A2(\u_lf.i_acc[5] ),
    .A1(net175));
 sg13g2_a21oi_2 _1163_ (.B1(_0535_),
    .Y(_0540_),
    .A2(_0539_),
    .A1(_0530_));
 sg13g2_and2_1 _1164_ (.A(net173),
    .B(\u_lf.i_acc[6] ),
    .X(_0541_));
 sg13g2_xor2_1 _1165_ (.B(net300),
    .A(net173),
    .X(_0542_));
 sg13g2_inv_1 _1166_ (.Y(_0543_),
    .A(_0542_));
 sg13g2_o21ai_1 _1167_ (.B1(net159),
    .Y(_0544_),
    .A1(_0540_),
    .A2(_0542_));
 sg13g2_a21oi_1 _1168_ (.A1(_0540_),
    .A2(_0542_),
    .Y(_0545_),
    .B1(_0544_));
 sg13g2_a21o_1 _1169_ (.A2(net166),
    .A1(net300),
    .B1(_0545_),
    .X(_0117_));
 sg13g2_nor2_1 _1170_ (.A(net298),
    .B(net159),
    .Y(_0546_));
 sg13g2_xnor2_1 _1171_ (.Y(_0547_),
    .A(net173),
    .B(net298));
 sg13g2_a21oi_1 _1172_ (.A1(_0540_),
    .A2(_0542_),
    .Y(_0548_),
    .B1(_0541_));
 sg13g2_xnor2_1 _1173_ (.Y(_0549_),
    .A(_0547_),
    .B(_0548_));
 sg13g2_a21oi_1 _1174_ (.A1(net159),
    .A2(_0549_),
    .Y(_0118_),
    .B1(_0546_));
 sg13g2_nor2_1 _1175_ (.A(_0543_),
    .B(_0547_),
    .Y(_0550_));
 sg13g2_o21ai_1 _1176_ (.B1(net174),
    .Y(_0551_),
    .A1(\u_lf.i_acc[7] ),
    .A2(\u_lf.i_acc[6] ));
 sg13g2_inv_1 _1177_ (.Y(_0552_),
    .A(_0551_));
 sg13g2_a21o_2 _1178_ (.A2(_0550_),
    .A1(_0540_),
    .B1(_0552_),
    .X(_0553_));
 sg13g2_xor2_1 _1179_ (.B(net239),
    .A(net174),
    .X(_0554_));
 sg13g2_and2_1 _1180_ (.A(_0553_),
    .B(_0554_),
    .X(_0555_));
 sg13g2_nand2_1 _1181_ (.Y(_0556_),
    .A(net239),
    .B(net165));
 sg13g2_o21ai_1 _1182_ (.B1(net158),
    .Y(_0557_),
    .A1(_0553_),
    .A2(_0554_));
 sg13g2_o21ai_1 _1183_ (.B1(_0556_),
    .Y(_0119_),
    .A1(_0555_),
    .A2(_0557_));
 sg13g2_nor2_1 _1184_ (.A(net272),
    .B(net157),
    .Y(_0558_));
 sg13g2_xor2_1 _1185_ (.B(net272),
    .A(net173),
    .X(_0559_));
 sg13g2_a21oi_1 _1186_ (.A1(net173),
    .A2(net239),
    .Y(_0560_),
    .B1(_0555_));
 sg13g2_xor2_1 _1187_ (.B(_0560_),
    .A(_0559_),
    .X(_0561_));
 sg13g2_a21oi_1 _1188_ (.A1(net157),
    .A2(_0561_),
    .Y(_0120_),
    .B1(_0558_));
 sg13g2_xnor2_1 _1189_ (.Y(_0562_),
    .A(net171),
    .B(net227));
 sg13g2_o21ai_1 _1190_ (.B1(net173),
    .Y(_0563_),
    .A1(\u_lf.i_acc[9] ),
    .A2(\u_lf.i_acc[8] ));
 sg13g2_nand2_1 _1191_ (.Y(_0564_),
    .A(_0555_),
    .B(_0559_));
 sg13g2_a21oi_1 _1192_ (.A1(_0563_),
    .A2(_0564_),
    .Y(_0565_),
    .B1(_0562_));
 sg13g2_nand3_1 _1193_ (.B(_0563_),
    .C(_0564_),
    .A(_0562_),
    .Y(_0566_));
 sg13g2_nand2_1 _1194_ (.Y(_0567_),
    .A(net227),
    .B(net165));
 sg13g2_nand2_1 _1195_ (.Y(_0568_),
    .A(net158),
    .B(_0566_));
 sg13g2_o21ai_1 _1196_ (.B1(_0567_),
    .Y(_0121_),
    .A1(_0565_),
    .A2(_0568_));
 sg13g2_nor2_1 _1197_ (.A(net279),
    .B(net158),
    .Y(_0569_));
 sg13g2_a21oi_1 _1198_ (.A1(net172),
    .A2(net227),
    .Y(_0570_),
    .B1(_0565_));
 sg13g2_xnor2_1 _1199_ (.Y(_0571_),
    .A(_0434_),
    .B(_0570_));
 sg13g2_a21oi_1 _1200_ (.A1(net158),
    .A2(_0571_),
    .Y(_0122_),
    .B1(_0569_));
 sg13g2_nand2_1 _1201_ (.Y(_0572_),
    .A(net106),
    .B(net165));
 sg13g2_o21ai_1 _1202_ (.B1(net172),
    .Y(_0573_),
    .A1(\u_lf.i_acc[11] ),
    .A2(\u_lf.i_acc[10] ));
 sg13g2_nand2_1 _1203_ (.Y(_0574_),
    .A(_0563_),
    .B(_0573_));
 sg13g2_inv_1 _1204_ (.Y(_0575_),
    .A(_0574_));
 sg13g2_nor2_1 _1205_ (.A(_0434_),
    .B(_0562_),
    .Y(_0576_));
 sg13g2_nand4_1 _1206_ (.B(_0554_),
    .C(_0559_),
    .A(_0553_),
    .Y(_0577_),
    .D(_0576_));
 sg13g2_and2_1 _1207_ (.A(_0575_),
    .B(_0577_),
    .X(_0578_));
 sg13g2_a21oi_1 _1208_ (.A1(_0575_),
    .A2(_0577_),
    .Y(_0579_),
    .B1(_0424_));
 sg13g2_a21o_1 _1209_ (.A2(_0578_),
    .A1(_0424_),
    .B1(net165),
    .X(_0580_));
 sg13g2_o21ai_1 _1210_ (.B1(_0572_),
    .Y(_0123_),
    .A1(_0579_),
    .A2(_0580_));
 sg13g2_nor2_1 _1211_ (.A(net262),
    .B(net157),
    .Y(_0581_));
 sg13g2_o21ai_1 _1212_ (.B1(_0419_),
    .Y(_0582_),
    .A1(_0424_),
    .A2(_0578_));
 sg13g2_xnor2_1 _1213_ (.Y(_0583_),
    .A(_0428_),
    .B(_0582_));
 sg13g2_a21oi_1 _1214_ (.A1(net157),
    .A2(_0583_),
    .Y(_0124_),
    .B1(_0581_));
 sg13g2_nor2_1 _1215_ (.A(net259),
    .B(net157),
    .Y(_0584_));
 sg13g2_a21o_1 _1216_ (.A2(_0579_),
    .A1(_0428_),
    .B1(_0420_),
    .X(_0585_));
 sg13g2_xor2_1 _1217_ (.B(_0585_),
    .A(_0426_),
    .X(_0586_));
 sg13g2_a21oi_1 _1218_ (.A1(net157),
    .A2(_0586_),
    .Y(_0125_),
    .B1(_0584_));
 sg13g2_nor2_1 _1219_ (.A(net266),
    .B(net157),
    .Y(_0587_));
 sg13g2_a21oi_1 _1220_ (.A1(_0425_),
    .A2(_0585_),
    .Y(_0588_),
    .B1(_0421_));
 sg13g2_xor2_1 _1221_ (.B(_0588_),
    .A(_0429_),
    .X(_0589_));
 sg13g2_a21oi_1 _1222_ (.A1(net157),
    .A2(_0589_),
    .Y(_0126_),
    .B1(_0587_));
 sg13g2_nand2_1 _1223_ (.Y(_0590_),
    .A(net87),
    .B(net167));
 sg13g2_and4_1 _1224_ (.A(_0431_),
    .B(_0554_),
    .C(_0559_),
    .D(_0576_),
    .X(_0591_));
 sg13g2_or2_1 _1225_ (.X(_0592_),
    .B(_0574_),
    .A(_0423_));
 sg13g2_a21oi_1 _1226_ (.A1(_0553_),
    .A2(_0591_),
    .Y(_0593_),
    .B1(_0592_));
 sg13g2_a21o_2 _1227_ (.A2(_0591_),
    .A1(_0553_),
    .B1(_0592_),
    .X(_0594_));
 sg13g2_xnor2_1 _1228_ (.Y(_0595_),
    .A(_0469_),
    .B(_0594_));
 sg13g2_o21ai_1 _1229_ (.B1(_0590_),
    .Y(_0127_),
    .A1(net167),
    .A2(_0595_));
 sg13g2_nor2_1 _1230_ (.A(net230),
    .B(net163),
    .Y(_0596_));
 sg13g2_a21oi_1 _1231_ (.A1(_0469_),
    .A2(_0594_),
    .Y(_0597_),
    .B1(_0407_));
 sg13g2_xor2_1 _1232_ (.B(_0597_),
    .A(_0468_),
    .X(_0598_));
 sg13g2_a21oi_1 _1233_ (.A1(net163),
    .A2(_0598_),
    .Y(_0128_),
    .B1(_0596_));
 sg13g2_nand3_1 _1234_ (.B(_0469_),
    .C(_0594_),
    .A(_0468_),
    .Y(_0599_));
 sg13g2_a21oi_1 _1235_ (.A1(_0408_),
    .A2(_0599_),
    .Y(_0600_),
    .B1(_0470_));
 sg13g2_nand3_1 _1236_ (.B(_0470_),
    .C(_0599_),
    .A(_0408_),
    .Y(_0601_));
 sg13g2_nand2_1 _1237_ (.Y(_0602_),
    .A(net72),
    .B(net167));
 sg13g2_nand2_1 _1238_ (.Y(_0603_),
    .A(net163),
    .B(_0601_));
 sg13g2_o21ai_1 _1239_ (.B1(_0602_),
    .Y(_0129_),
    .A1(_0600_),
    .A2(_0603_));
 sg13g2_nor2_1 _1240_ (.A(net264),
    .B(net163),
    .Y(_0604_));
 sg13g2_a21oi_1 _1241_ (.A1(net178),
    .A2(net72),
    .Y(_0605_),
    .B1(_0600_));
 sg13g2_xnor2_1 _1242_ (.Y(_0606_),
    .A(_0467_),
    .B(_0605_));
 sg13g2_a21oi_1 _1243_ (.A1(net163),
    .A2(_0606_),
    .Y(_0130_),
    .B1(_0604_));
 sg13g2_nor2_1 _1244_ (.A(net273),
    .B(net161),
    .Y(_0607_));
 sg13g2_a21o_2 _1245_ (.A2(_0594_),
    .A1(_0473_),
    .B1(_0410_),
    .X(_0608_));
 sg13g2_nand2b_1 _1246_ (.Y(_0609_),
    .B(_0608_),
    .A_N(_0475_));
 sg13g2_xor2_1 _1247_ (.B(_0608_),
    .A(_0475_),
    .X(_0610_));
 sg13g2_a21oi_1 _1248_ (.A1(net161),
    .A2(_0610_),
    .Y(_0131_),
    .B1(_0607_));
 sg13g2_nor2_1 _1249_ (.A(net218),
    .B(net161),
    .Y(_0611_));
 sg13g2_nand2_1 _1250_ (.Y(_0612_),
    .A(_0412_),
    .B(_0609_));
 sg13g2_xor2_1 _1251_ (.B(_0612_),
    .A(_0474_),
    .X(_0613_));
 sg13g2_a21oi_1 _1252_ (.A1(net161),
    .A2(_0613_),
    .Y(_0132_),
    .B1(_0611_));
 sg13g2_a21oi_1 _1253_ (.A1(_0476_),
    .A2(_0608_),
    .Y(_0614_),
    .B1(_0414_));
 sg13g2_xnor2_1 _1254_ (.Y(_0615_),
    .A(_0479_),
    .B(_0614_));
 sg13g2_mux2_1 _1255_ (.A0(net283),
    .A1(_0615_),
    .S(net161),
    .X(_0133_));
 sg13g2_nor2_1 _1256_ (.A(net232),
    .B(net161),
    .Y(_0616_));
 sg13g2_o21ai_1 _1257_ (.B1(_0411_),
    .Y(_0617_),
    .A1(_0478_),
    .A2(_0614_));
 sg13g2_xnor2_1 _1258_ (.Y(_0618_),
    .A(_0477_),
    .B(_0617_));
 sg13g2_a21oi_1 _1259_ (.A1(net162),
    .A2(_0618_),
    .Y(_0134_),
    .B1(_0616_));
 sg13g2_o21ai_1 _1260_ (.B1(_0417_),
    .Y(_0619_),
    .A1(_0480_),
    .A2(_0593_));
 sg13g2_nand2b_1 _1261_ (.Y(_0620_),
    .B(_0619_),
    .A_N(_0483_));
 sg13g2_nor2_1 _1262_ (.A(net267),
    .B(net162),
    .Y(_0621_));
 sg13g2_xor2_1 _1263_ (.B(_0619_),
    .A(_0483_),
    .X(_0622_));
 sg13g2_a21oi_1 _1264_ (.A1(net162),
    .A2(_0622_),
    .Y(_0135_),
    .B1(_0621_));
 sg13g2_nor2_1 _1265_ (.A(net303),
    .B(net162),
    .Y(_0623_));
 sg13g2_nand2_1 _1266_ (.Y(_0624_),
    .A(_0404_),
    .B(_0620_));
 sg13g2_xnor2_1 _1267_ (.Y(_0625_),
    .A(_0484_),
    .B(_0624_));
 sg13g2_a21oi_1 _1268_ (.A1(net162),
    .A2(_0625_),
    .Y(_0136_),
    .B1(_0623_));
 sg13g2_nor2_1 _1269_ (.A(net252),
    .B(net160),
    .Y(_0626_));
 sg13g2_a21oi_1 _1270_ (.A1(_0485_),
    .A2(_0619_),
    .Y(_0627_),
    .B1(_0406_));
 sg13g2_xor2_1 _1271_ (.B(_0627_),
    .A(_0402_),
    .X(_0628_));
 sg13g2_a21oi_1 _1272_ (.A1(net160),
    .A2(_0628_),
    .Y(_0137_),
    .B1(_0626_));
 sg13g2_nor2_1 _1273_ (.A(net236),
    .B(net160),
    .Y(_0629_));
 sg13g2_o21ai_1 _1274_ (.B1(_0400_),
    .Y(_0630_),
    .A1(_0401_),
    .A2(_0627_));
 sg13g2_xnor2_1 _1275_ (.Y(_0631_),
    .A(_0399_),
    .B(_0630_));
 sg13g2_a21oi_1 _1276_ (.A1(net160),
    .A2(_0631_),
    .Y(_0138_),
    .B1(_0629_));
 sg13g2_nor2_1 _1277_ (.A(net257),
    .B(net160),
    .Y(_0632_));
 sg13g2_a21oi_1 _1278_ (.A1(_0501_),
    .A2(_0619_),
    .Y(_0633_),
    .B1(_0500_));
 sg13g2_xnor2_1 _1279_ (.Y(_0634_),
    .A(_0504_),
    .B(_0633_));
 sg13g2_a21oi_1 _1280_ (.A1(net161),
    .A2(_0634_),
    .Y(_0139_),
    .B1(_0632_));
 sg13g2_nor2_1 _1281_ (.A(net138),
    .B(net160),
    .Y(_0635_));
 sg13g2_o21ai_1 _1282_ (.B1(_0503_),
    .Y(_0636_),
    .A1(_0504_),
    .A2(_0633_));
 sg13g2_xnor2_1 _1283_ (.Y(_0637_),
    .A(_0508_),
    .B(_0636_));
 sg13g2_a21oi_1 _1284_ (.A1(net160),
    .A2(_0637_),
    .Y(_0140_),
    .B1(_0635_));
 sg13g2_dfrbpq_1 _1285_ (.RESET_B(net201),
    .D(net22),
    .Q(helper_msb_d),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1286_ (.RESET_B(net195),
    .D(net108),
    .Q(\u_core.ref_samp_d ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1287_ (.RESET_B(net193),
    .D(_0002_),
    .Q(\u_core.beat_cnt[0] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1288_ (.RESET_B(net191),
    .D(_0003_),
    .Q(\u_core.beat_cnt[1] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1289_ (.RESET_B(net190),
    .D(net28),
    .Q(\u_core.beat_cnt[2] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_2 _1290_ (.RESET_B(net190),
    .D(net55),
    .Q(\u_core.beat_cnt[3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1291_ (.RESET_B(net190),
    .D(_0006_),
    .Q(\u_core.beat_cnt[4] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1292_ (.RESET_B(net189),
    .D(net24),
    .Q(\u_core.beat_cnt[5] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1293_ (.RESET_B(net189),
    .D(net53),
    .Q(\u_core.beat_cnt[6] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1294_ (.RESET_B(net189),
    .D(_0009_),
    .Q(\u_core.beat_cnt[7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1295_ (.RESET_B(net189),
    .D(net26),
    .Q(\u_core.beat_cnt[8] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1296_ (.RESET_B(net185),
    .D(net36),
    .Q(\u_core.beat_cnt[9] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1297_ (.RESET_B(net184),
    .D(net47),
    .Q(\u_core.beat_cnt[10] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1298_ (.RESET_B(net184),
    .D(_0013_),
    .Q(\u_core.beat_cnt[11] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1299_ (.RESET_B(net183),
    .D(net60),
    .Q(\u_core.beat_cnt[12] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1300_ (.RESET_B(net183),
    .D(_0015_),
    .Q(\u_core.beat_cnt[13] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1301_ (.RESET_B(net183),
    .D(net62),
    .Q(\u_core.beat_cnt[14] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1302_ (.RESET_B(net186),
    .D(net44),
    .Q(\u_core.beat_cnt[15] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1303_ (.RESET_B(net194),
    .D(net38),
    .Q(\phase_err_beat[4] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1304_ (.RESET_B(net194),
    .D(net254),
    .Q(\phase_err_beat[5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1305_ (.RESET_B(net194),
    .D(_0020_),
    .Q(\phase_err_beat[6] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1306_ (.RESET_B(net194),
    .D(net244),
    .Q(\phase_err_beat[7] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1307_ (.RESET_B(net187),
    .D(net241),
    .Q(\phase_err_beat[8] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1308_ (.RESET_B(net187),
    .D(net261),
    .Q(\phase_err_beat[9] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1309_ (.RESET_B(net187),
    .D(net306),
    .Q(\phase_err_beat[10] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1310_ (.RESET_B(net187),
    .D(net226),
    .Q(\phase_err_beat[11] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_2 _1311_ (.RESET_B(net187),
    .D(net294),
    .Q(\phase_err_beat[12] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1312_ (.RESET_B(net187),
    .D(net133),
    .Q(\phase_err_beat[13] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1313_ (.RESET_B(net187),
    .D(_0028_),
    .Q(\phase_err_beat[14] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1314_ (.RESET_B(net188),
    .D(_0029_),
    .Q(\phase_err_beat[15] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1315_ (.RESET_B(net193),
    .D(_0030_),
    .Q(\u_core.t_ref[0] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1316_ (.RESET_B(net191),
    .D(net246),
    .Q(\u_core.t_ref[1] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1317_ (.RESET_B(net190),
    .D(_0032_),
    .Q(\u_core.t_ref[2] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1318_ (.RESET_B(net190),
    .D(_0033_),
    .Q(\u_core.t_ref[3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1319_ (.RESET_B(net191),
    .D(_0034_),
    .Q(\u_core.t_ref[4] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1320_ (.RESET_B(net192),
    .D(_0035_),
    .Q(\u_core.t_ref[5] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1321_ (.RESET_B(net189),
    .D(_0036_),
    .Q(\u_core.t_ref[6] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1322_ (.RESET_B(net189),
    .D(net278),
    .Q(\u_core.t_ref[7] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1323_ (.RESET_B(net184),
    .D(_0038_),
    .Q(\u_core.t_ref[8] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1324_ (.RESET_B(net185),
    .D(_0039_),
    .Q(\u_core.t_ref[9] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1325_ (.RESET_B(net184),
    .D(_0040_),
    .Q(\u_core.t_ref[10] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1326_ (.RESET_B(net184),
    .D(_0041_),
    .Q(\u_core.t_ref[11] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1327_ (.RESET_B(net183),
    .D(_0042_),
    .Q(\u_core.t_ref[12] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1328_ (.RESET_B(net183),
    .D(_0043_),
    .Q(\u_core.t_ref[13] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1329_ (.RESET_B(net183),
    .D(_0044_),
    .Q(\u_core.t_ref[14] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1330_ (.RESET_B(net188),
    .D(_0045_),
    .Q(\u_core.t_ref[15] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1331_ (.RESET_B(net206),
    .D(clk_fb),
    .Q(\u_core.fb_sync[0] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1332_ (.RESET_B(net202),
    .D(net20),
    .Q(\u_core.fb_sync[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1333_ (.RESET_B(net205),
    .D(net1),
    .Q(\u_core.ref_sync[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1334_ (.RESET_B(net205),
    .D(net21),
    .Q(\u_core.ref_sync[1] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1335_ (.RESET_B(net201),
    .D(net75),
    .Q(fb_samp),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1336_ (.RESET_B(net193),
    .D(_0047_),
    .Q(\u_core.t_fb[0] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1337_ (.RESET_B(net191),
    .D(net215),
    .Q(\u_core.t_fb[1] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1338_ (.RESET_B(net190),
    .D(_0049_),
    .Q(\u_core.t_fb[2] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1339_ (.RESET_B(net190),
    .D(_0050_),
    .Q(\u_core.t_fb[3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1340_ (.RESET_B(net190),
    .D(net281),
    .Q(\u_core.t_fb[4] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1341_ (.RESET_B(net192),
    .D(_0052_),
    .Q(\u_core.t_fb[5] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1342_ (.RESET_B(net189),
    .D(_0053_),
    .Q(\u_core.t_fb[6] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1343_ (.RESET_B(net189),
    .D(net286),
    .Q(\u_core.t_fb[7] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1344_ (.RESET_B(net184),
    .D(_0055_),
    .Q(\u_core.t_fb[8] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1345_ (.RESET_B(net185),
    .D(_0056_),
    .Q(\u_core.t_fb[9] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1346_ (.RESET_B(net184),
    .D(_0057_),
    .Q(\u_core.t_fb[10] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1347_ (.RESET_B(net184),
    .D(_0058_),
    .Q(\u_core.t_fb[11] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1348_ (.RESET_B(net183),
    .D(_0059_),
    .Q(\u_core.t_fb[12] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1349_ (.RESET_B(net186),
    .D(net86),
    .Q(\u_core.t_fb[13] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1350_ (.RESET_B(net183),
    .D(_0061_),
    .Q(\u_core.t_fb[14] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1351_ (.RESET_B(net188),
    .D(_0062_),
    .Q(\u_core.t_fb[15] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1352_ (.RESET_B(net201),
    .D(net126),
    .Q(ref_samp),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1353_ (.RESET_B(net195),
    .D(net58),
    .Q(\u_core.fb_samp_d ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1354_ (.RESET_B(net194),
    .D(net146),
    .Q(phase_valid),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1355_ (.RESET_B(net193),
    .D(_0065_),
    .Q(\u_core.have_ref ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1356_ (.RESET_B(net199),
    .D(net34),
    .Q(\nco_phase_acc[0] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1357_ (.RESET_B(net199),
    .D(_0067_),
    .Q(\nco_phase_acc[1] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1358_ (.RESET_B(net203),
    .D(net118),
    .Q(\nco_phase_acc[2] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1359_ (.RESET_B(net203),
    .D(_0069_),
    .Q(\nco_phase_acc[3] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1360_ (.RESET_B(net204),
    .D(net217),
    .Q(\nco_phase_acc[4] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1361_ (.RESET_B(net204),
    .D(net110),
    .Q(\nco_phase_acc[5] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1362_ (.RESET_B(net205),
    .D(net223),
    .Q(\nco_phase_acc[6] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1363_ (.RESET_B(net206),
    .D(net120),
    .Q(\nco_phase_acc[7] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1364_ (.RESET_B(net201),
    .D(_0074_),
    .Q(\nco_phase_acc[8] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1365_ (.RESET_B(net201),
    .D(net82),
    .Q(\nco_phase_acc[9] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1366_ (.RESET_B(net202),
    .D(_0076_),
    .Q(\nco_phase_acc[10] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _1367_ (.RESET_B(net202),
    .D(net124),
    .Q(\nco_phase_acc[11] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1368_ (.RESET_B(net202),
    .D(_0078_),
    .Q(\nco_phase_acc[12] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1369_ (.RESET_B(net203),
    .D(net100),
    .Q(\nco_phase_acc[13] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1370_ (.RESET_B(net203),
    .D(net113),
    .Q(\nco_phase_acc[14] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1371_ (.RESET_B(net203),
    .D(net248),
    .Q(\nco_phase_acc[15] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1372_ (.RESET_B(net206),
    .D(_0082_),
    .Q(\nco_phase_acc[16] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1373_ (.RESET_B(net206),
    .D(_0083_),
    .Q(\nco_phase_acc[17] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1374_ (.RESET_B(net206),
    .D(net32),
    .Q(\nco_phase_acc[18] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1375_ (.RESET_B(net205),
    .D(_0085_),
    .Q(\nco_phase_acc[19] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1376_ (.RESET_B(net205),
    .D(net40),
    .Q(\nco_phase_acc[20] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1377_ (.RESET_B(net205),
    .D(net78),
    .Q(\nco_phase_acc[21] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1378_ (.RESET_B(net207),
    .D(net30),
    .Q(\nco_phase_acc[22] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1379_ (.RESET_B(net206),
    .D(_0089_),
    .Q(clk_helper),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1380_ (.RESET_B(net201),
    .D(_0090_),
    .Q(\ctrl[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1381_ (.RESET_B(net193),
    .D(_0091_),
    .Q(\ctrl[1] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1382_ (.RESET_B(net193),
    .D(_0092_),
    .Q(\ctrl[2] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1383_ (.RESET_B(net193),
    .D(_0093_),
    .Q(\ctrl[3] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_1 _1384_ (.RESET_B(net199),
    .D(net68),
    .Q(\ctrl[8] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1385_ (.RESET_B(net199),
    .D(net129),
    .Q(\ctrl[9] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1386_ (.RESET_B(net199),
    .D(net103),
    .Q(\ctrl[10] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1387_ (.RESET_B(net204),
    .D(net49),
    .Q(\ctrl[11] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1388_ (.RESET_B(net204),
    .D(net105),
    .Q(\ctrl[12] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _1389_ (.RESET_B(net205),
    .D(net84),
    .Q(\ctrl[13] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1390_ (.RESET_B(net205),
    .D(net94),
    .Q(\ctrl[14] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1391_ (.RESET_B(net206),
    .D(net137),
    .Q(\ctrl[15] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_1 _1392_ (.RESET_B(net201),
    .D(net141),
    .Q(\ctrl[16] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1393_ (.RESET_B(net201),
    .D(net71),
    .Q(\ctrl[17] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1394_ (.RESET_B(net202),
    .D(_0104_),
    .Q(\ctrl[18] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1395_ (.RESET_B(net202),
    .D(_0105_),
    .Q(\ctrl[19] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1396_ (.RESET_B(net202),
    .D(net98),
    .Q(\ctrl[20] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1397_ (.RESET_B(net203),
    .D(net90),
    .Q(\ctrl[21] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1398_ (.RESET_B(net203),
    .D(net122),
    .Q(\ctrl[22] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1399_ (.RESET_B(net203),
    .D(net251),
    .Q(\ctrl[23] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1400_ (.RESET_B(net193),
    .D(_0110_),
    .Q(\u_core.have_fb ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_2 _1401_ (.RESET_B(net194),
    .D(net51),
    .Q(\u_lf.i_acc[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1402_ (.RESET_B(net194),
    .D(_0112_),
    .Q(\u_lf.i_acc[1] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1403_ (.RESET_B(net194),
    .D(net115),
    .Q(\u_lf.i_acc[2] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1404_ (.RESET_B(net196),
    .D(net271),
    .Q(\u_lf.i_acc[3] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1405_ (.RESET_B(net187),
    .D(net275),
    .Q(\u_lf.i_acc[4] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1406_ (.RESET_B(net188),
    .D(net291),
    .Q(\u_lf.i_acc[5] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1407_ (.RESET_B(net197),
    .D(_0117_),
    .Q(\u_lf.i_acc[6] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1408_ (.RESET_B(net200),
    .D(net299),
    .Q(\u_lf.i_acc[7] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1409_ (.RESET_B(net200),
    .D(_0119_),
    .Q(\u_lf.i_acc[8] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1410_ (.RESET_B(net197),
    .D(_0120_),
    .Q(\u_lf.i_acc[9] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1411_ (.RESET_B(net188),
    .D(net228),
    .Q(\u_lf.i_acc[10] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1412_ (.RESET_B(net188),
    .D(_0122_),
    .Q(\u_lf.i_acc[11] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1413_ (.RESET_B(net197),
    .D(_0123_),
    .Q(\u_lf.i_acc[12] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1414_ (.RESET_B(net197),
    .D(_0124_),
    .Q(\u_lf.i_acc[13] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1415_ (.RESET_B(net197),
    .D(_0125_),
    .Q(\u_lf.i_acc[14] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1416_ (.RESET_B(net188),
    .D(_0126_),
    .Q(\u_lf.i_acc[15] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1417_ (.RESET_B(net197),
    .D(net88),
    .Q(\u_lf.i_acc[16] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1418_ (.RESET_B(net199),
    .D(_0128_),
    .Q(\u_lf.i_acc[17] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1419_ (.RESET_B(net199),
    .D(net73),
    .Q(\u_lf.i_acc[18] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1420_ (.RESET_B(net199),
    .D(_0130_),
    .Q(\u_lf.i_acc[19] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1421_ (.RESET_B(net198),
    .D(_0131_),
    .Q(\u_lf.i_acc[20] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1422_ (.RESET_B(net198),
    .D(net219),
    .Q(\u_lf.i_acc[21] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1423_ (.RESET_B(net198),
    .D(_0133_),
    .Q(\u_lf.i_acc[22] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1424_ (.RESET_B(net198),
    .D(net233),
    .Q(\u_lf.i_acc[23] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1425_ (.RESET_B(net197),
    .D(net268),
    .Q(\u_lf.i_acc[24] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1426_ (.RESET_B(net197),
    .D(_0136_),
    .Q(\u_lf.i_acc[25] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1427_ (.RESET_B(net198),
    .D(_0137_),
    .Q(\u_lf.i_acc[26] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1428_ (.RESET_B(net198),
    .D(net237),
    .Q(\u_lf.i_acc[27] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1429_ (.RESET_B(net198),
    .D(net258),
    .Q(\u_lf.i_acc[28] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1430_ (.RESET_B(net198),
    .D(net139),
    .Q(\u_lf.i_acc[29] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_tielo tt_um_arthfink_ddmtd_5 (.L_LO(net5));
 sg13g2_tielo tt_um_arthfink_ddmtd_6 (.L_LO(net6));
 sg13g2_tielo tt_um_arthfink_ddmtd_7 (.L_LO(net7));
 sg13g2_tielo tt_um_arthfink_ddmtd_8 (.L_LO(net8));
 sg13g2_tielo tt_um_arthfink_ddmtd_9 (.L_LO(net9));
 sg13g2_tielo tt_um_arthfink_ddmtd_10 (.L_LO(net10));
 sg13g2_tielo tt_um_arthfink_ddmtd_11 (.L_LO(net11));
 sg13g2_tielo tt_um_arthfink_ddmtd_12 (.L_LO(net12));
 sg13g2_tielo tt_um_arthfink_ddmtd_13 (.L_LO(net13));
 sg13g2_tielo tt_um_arthfink_ddmtd_14 (.L_LO(net14));
 sg13g2_tielo tt_um_arthfink_ddmtd_15 (.L_LO(net15));
 sg13g2_tielo tt_um_arthfink_ddmtd_16 (.L_LO(net16));
 sg13g2_tielo tt_um_arthfink_ddmtd_17 (.L_LO(net17));
 sg13g2_tielo tt_um_arthfink_ddmtd_18 (.L_LO(net18));
 sg13g2_tielo tt_um_arthfink_ddmtd_19 (.L_LO(net19));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 fanout143 (.A(net145),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(net145),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0510_),
    .X(net145));
 sg13g2_buf_8 fanout146 (.A(_0000_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(net148),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(net150),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(_0282_),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(net152),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(net154),
    .X(net152));
 sg13g2_buf_8 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_8 fanout154 (.A(_0275_),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(_0183_),
    .X(net155));
 sg13g2_buf_1 fanout156 (.A(_0183_),
    .X(net156));
 sg13g2_buf_8 fanout157 (.A(net158),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_1 fanout159 (.A(uo_out[0]),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(net161),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(net162),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(net163),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(uo_out[0]),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(net164),
    .X(uo_out[0]));
 sg13g2_buf_8 fanout165 (.A(net166),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net170),
    .X(net166));
 sg13g2_buf_1 fanout167 (.A(net170),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net170),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(_0184_),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(net174),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_1 fanout175 (.A(net312),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(net180),
    .X(net176));
 sg13g2_buf_1 fanout177 (.A(net180),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net180),
    .X(net178));
 sg13g2_buf_1 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net181),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(\phase_err_beat[15] ),
    .X(net181));
 sg13g2_buf_8 fanout182 (.A(_0141_),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(net186),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(net185),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(net186),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(net196),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(net196),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(net192),
    .X(net189));
 sg13g2_buf_8 fanout190 (.A(net192),
    .X(net190));
 sg13g2_buf_1 fanout191 (.A(net192),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(net195),
    .X(net192));
 sg13g2_buf_8 fanout193 (.A(net195),
    .X(net193));
 sg13g2_buf_8 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_8 fanout195 (.A(net196),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(net208),
    .X(net196));
 sg13g2_buf_8 fanout197 (.A(net200),
    .X(net197));
 sg13g2_buf_8 fanout198 (.A(net200),
    .X(net198));
 sg13g2_buf_8 fanout199 (.A(net200),
    .X(net199));
 sg13g2_buf_8 fanout200 (.A(net208),
    .X(net200));
 sg13g2_buf_8 fanout201 (.A(net202),
    .X(net201));
 sg13g2_buf_8 fanout202 (.A(net208),
    .X(net202));
 sg13g2_buf_8 fanout203 (.A(net207),
    .X(net203));
 sg13g2_buf_1 fanout204 (.A(net207),
    .X(net204));
 sg13g2_buf_8 fanout205 (.A(net206),
    .X(net205));
 sg13g2_buf_8 fanout206 (.A(net207),
    .X(net206));
 sg13g2_buf_8 fanout207 (.A(net208),
    .X(net207));
 sg13g2_buf_8 fanout208 (.A(rst_n),
    .X(net208));
 sg13g2_buf_8 fanout209 (.A(net214),
    .X(net209));
 sg13g2_buf_8 fanout210 (.A(net214),
    .X(net210));
 sg13g2_buf_8 fanout211 (.A(net213),
    .X(net211));
 sg13g2_buf_1 fanout212 (.A(net213),
    .X(net212));
 sg13g2_buf_8 fanout213 (.A(net214),
    .X(net213));
 sg13g2_buf_8 fanout214 (.A(ena),
    .X(net214));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_tielo tt_um_arthfink_ddmtd_4 (.L_LO(net4));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_5_16__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload15 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_core.fb_sync[0] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_core.ref_sync[0] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold3 (.A(clk_helper),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold4 (.A(\u_core.beat_cnt[5] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0007_),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u_core.beat_cnt[8] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0010_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u_core.beat_cnt[2] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0004_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold10 (.A(\nco_phase_acc[22] ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0088_),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold12 (.A(\nco_phase_acc[18] ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0084_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold14 (.A(\nco_phase_acc[0] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0066_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u_core.beat_cnt[9] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0011_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold18 (.A(\phase_err_beat[4] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0018_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold20 (.A(\nco_phase_acc[20] ),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0086_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ctrl[0] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_core.beat_cnt[0] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold24 (.A(\u_core.beat_cnt[15] ),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0017_),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ctrl[1] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_core.beat_cnt[10] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0012_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ctrl[11] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0097_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_lf.i_acc[0] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0111_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_core.beat_cnt[6] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0008_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_core.beat_cnt[3] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0005_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold37 (.A(\ctrl[3] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u_core.fb_samp_d ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0064_),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u_core.beat_cnt[12] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0014_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold42 (.A(\u_core.beat_cnt[14] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0016_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold44 (.A(\ctrl[2] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold45 (.A(\nco_phase_acc[21] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0398_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u_core.t_ref[9] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold48 (.A(\ctrl[8] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0094_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u_core.beat_cnt[11] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold51 (.A(\ctrl[17] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0103_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u_lf.i_acc[18] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0129_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u_core.fb_sync[1] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0046_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold57 (.A(\nco_phase_acc[19] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0395_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0087_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold60 (.A(\nco_phase_acc[16] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0388_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold62 (.A(\nco_phase_acc[9] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0075_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ctrl[13] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0099_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_core.beat_cnt[13] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0060_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold68 (.A(\u_lf.i_acc[16] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0127_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold70 (.A(\ctrl[21] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold71 (.A(_0107_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold72 (.A(\u_core.t_ref[13] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold73 (.A(\nco_phase_acc[17] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold74 (.A(\ctrl[14] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold75 (.A(_0100_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold76 (.A(\ctrl[18] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold77 (.A(\u_core.t_fb[9] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold78 (.A(\ctrl[20] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0106_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold80 (.A(\nco_phase_acc[13] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0079_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold82 (.A(\u_core.t_fb[2] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ctrl[10] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0096_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ctrl[12] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0098_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold87 (.A(\u_lf.i_acc[12] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold88 (.A(\u_core.ref_samp_d ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0001_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold90 (.A(\nco_phase_acc[5] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0071_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold92 (.A(\u_core.t_ref[2] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold93 (.A(\nco_phase_acc[14] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0080_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold95 (.A(\u_lf.i_acc[2] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0113_),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_core.t_ref[0] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold98 (.A(\nco_phase_acc[2] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0068_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold100 (.A(\nco_phase_acc[7] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0073_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold102 (.A(\ctrl[22] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0108_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold104 (.A(\nco_phase_acc[11] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0077_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold106 (.A(\u_core.ref_sync[1] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0063_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold108 (.A(\nco_phase_acc[10] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ctrl[9] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0095_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold111 (.A(\nco_phase_acc[12] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold112 (.A(\phase_err_beat[13] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0262_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0027_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold115 (.A(\nco_phase_acc[1] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold116 (.A(\u_core.t_fb[0] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold117 (.A(\ctrl[15] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0101_),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold119 (.A(\u_lf.i_acc[29] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0140_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold121 (.A(\ctrl[16] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0102_),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_core.t_fb[1] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold124 (.A(_0048_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold125 (.A(\nco_phase_acc[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0070_),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_lf.i_acc[21] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0132_),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold129 (.A(\u_core.t_fb[11] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_core.t_ref[15] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold131 (.A(\nco_phase_acc[6] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold132 (.A(_0072_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold133 (.A(\phase_err_beat[11] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold134 (.A(_0252_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0025_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_lf.i_acc[10] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0121_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold138 (.A(\nco_phase_acc[3] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_lf.i_acc[17] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold140 (.A(\u_core.t_fb[8] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold141 (.A(\u_lf.i_acc[23] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0134_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold143 (.A(\u_core.t_fb[14] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold144 (.A(\u_core.t_ref[8] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_lf.i_acc[27] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0138_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_core.t_ref[11] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold148 (.A(\u_lf.i_acc[8] ),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold149 (.A(\phase_err_beat[8] ),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold150 (.A(_0022_),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold151 (.A(\phase_err_beat[6] ),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold152 (.A(\phase_err_beat[7] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold153 (.A(_0021_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_core.t_ref[1] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0031_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold156 (.A(\nco_phase_acc[15] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0081_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold158 (.A(\u_core.t_ref[14] ),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold159 (.A(\ctrl[23] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0109_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold161 (.A(\u_lf.i_acc[26] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold162 (.A(\phase_err_beat[5] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold163 (.A(_0019_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold164 (.A(\u_core.t_fb[5] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold165 (.A(\u_core.t_ref[5] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold166 (.A(\u_lf.i_acc[28] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0139_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold168 (.A(\u_lf.i_acc[14] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold169 (.A(\phase_err_beat[9] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0023_),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold171 (.A(\u_lf.i_acc[13] ),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_core.have_fb ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold173 (.A(\u_lf.i_acc[19] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_core.t_fb[15] ),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_lf.i_acc[15] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_lf.i_acc[24] ),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0135_),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold178 (.A(\u_core.t_ref[12] ),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_lf.i_acc[3] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0114_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_lf.i_acc[9] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold182 (.A(\u_lf.i_acc[20] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold183 (.A(\u_lf.i_acc[4] ),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0115_),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold185 (.A(\u_core.have_ref ),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_core.t_ref[7] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0037_),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold188 (.A(\u_lf.i_acc[11] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_core.beat_cnt[4] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold190 (.A(_0051_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold191 (.A(\ctrl[19] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold192 (.A(\u_lf.i_acc[22] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_core.t_ref[10] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold194 (.A(\u_core.t_fb[7] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0054_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold196 (.A(\u_core.t_fb[10] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_core.t_fb[6] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold198 (.A(\u_core.t_ref[6] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_lf.i_acc[5] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0116_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_core.t_ref[4] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold202 (.A(\phase_err_beat[12] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0026_),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold204 (.A(\u_core.t_fb[3] ),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_core.t_fb[12] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold206 (.A(\nco_phase_acc[8] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold207 (.A(\u_lf.i_acc[7] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold208 (.A(_0118_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold209 (.A(\u_lf.i_acc[6] ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold210 (.A(\u_lf.i_acc[1] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0518_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold212 (.A(\u_lf.i_acc[25] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold213 (.A(\u_core.t_ref[3] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold214 (.A(\phase_err_beat[10] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0024_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold216 (.A(\phase_err_beat[14] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold217 (.A(\u_core.beat_cnt[1] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold218 (.A(\nco_phase_acc[15] ),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold219 (.A(_0385_),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold220 (.A(\u_core.beat_cnt[7] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold221 (.A(\phase_err_beat[15] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold222 (.A(\u_lf.i_acc[13] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_core.t_ref[6] ),
    .X(net314));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_fill_2 FILLER_4_315 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_fill_1 FILLER_4_343 ();
 sg13g2_fill_2 FILLER_4_348 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_2 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_5_200 ();
 sg13g2_fill_1 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_215 ();
 sg13g2_decap_8 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_229 ();
 sg13g2_decap_8 FILLER_5_236 ();
 sg13g2_decap_8 FILLER_5_243 ();
 sg13g2_decap_8 FILLER_5_250 ();
 sg13g2_decap_8 FILLER_5_257 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_fill_2 FILLER_5_271 ();
 sg13g2_fill_1 FILLER_5_273 ();
 sg13g2_fill_2 FILLER_5_278 ();
 sg13g2_fill_1 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_4 FILLER_5_304 ();
 sg13g2_fill_2 FILLER_5_313 ();
 sg13g2_decap_4 FILLER_5_332 ();
 sg13g2_fill_2 FILLER_5_341 ();
 sg13g2_fill_1 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_377 ();
 sg13g2_decap_8 FILLER_6_384 ();
 sg13g2_decap_8 FILLER_6_391 ();
 sg13g2_decap_8 FILLER_6_398 ();
 sg13g2_decap_4 FILLER_6_405 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_4 FILLER_7_147 ();
 sg13g2_fill_1 FILLER_7_151 ();
 sg13g2_fill_2 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_181 ();
 sg13g2_decap_8 FILLER_7_242 ();
 sg13g2_decap_4 FILLER_7_249 ();
 sg13g2_fill_1 FILLER_7_305 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_fill_1 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_377 ();
 sg13g2_decap_8 FILLER_7_384 ();
 sg13g2_decap_8 FILLER_7_391 ();
 sg13g2_decap_8 FILLER_7_398 ();
 sg13g2_decap_4 FILLER_7_405 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_fill_2 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_47 ();
 sg13g2_fill_1 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_4 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_93 ();
 sg13g2_decap_8 FILLER_8_103 ();
 sg13g2_decap_8 FILLER_8_110 ();
 sg13g2_decap_8 FILLER_8_117 ();
 sg13g2_decap_8 FILLER_8_124 ();
 sg13g2_decap_8 FILLER_8_131 ();
 sg13g2_decap_8 FILLER_8_138 ();
 sg13g2_decap_8 FILLER_8_145 ();
 sg13g2_decap_8 FILLER_8_152 ();
 sg13g2_fill_2 FILLER_8_163 ();
 sg13g2_fill_1 FILLER_8_165 ();
 sg13g2_fill_2 FILLER_8_207 ();
 sg13g2_fill_1 FILLER_8_223 ();
 sg13g2_decap_8 FILLER_8_251 ();
 sg13g2_fill_2 FILLER_8_258 ();
 sg13g2_fill_1 FILLER_8_260 ();
 sg13g2_fill_2 FILLER_8_275 ();
 sg13g2_fill_1 FILLER_8_310 ();
 sg13g2_fill_1 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_329 ();
 sg13g2_fill_1 FILLER_8_331 ();
 sg13g2_fill_2 FILLER_8_353 ();
 sg13g2_fill_1 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_4 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_fill_2 FILLER_9_71 ();
 sg13g2_fill_1 FILLER_9_73 ();
 sg13g2_decap_8 FILLER_9_111 ();
 sg13g2_decap_8 FILLER_9_118 ();
 sg13g2_decap_8 FILLER_9_125 ();
 sg13g2_decap_8 FILLER_9_132 ();
 sg13g2_decap_8 FILLER_9_139 ();
 sg13g2_decap_4 FILLER_9_146 ();
 sg13g2_fill_1 FILLER_9_150 ();
 sg13g2_fill_1 FILLER_9_177 ();
 sg13g2_fill_2 FILLER_9_191 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_234 ();
 sg13g2_decap_8 FILLER_9_241 ();
 sg13g2_decap_8 FILLER_9_248 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_fill_1 FILLER_9_262 ();
 sg13g2_fill_2 FILLER_9_276 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_2 FILLER_9_306 ();
 sg13g2_fill_1 FILLER_9_313 ();
 sg13g2_fill_1 FILLER_9_319 ();
 sg13g2_fill_2 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_2 FILLER_10_11 ();
 sg13g2_fill_2 FILLER_10_41 ();
 sg13g2_fill_1 FILLER_10_83 ();
 sg13g2_decap_8 FILLER_10_111 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_decap_8 FILLER_10_125 ();
 sg13g2_decap_4 FILLER_10_132 ();
 sg13g2_fill_2 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_166 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_fill_2 FILLER_10_206 ();
 sg13g2_decap_4 FILLER_10_229 ();
 sg13g2_fill_2 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_fill_2 FILLER_10_255 ();
 sg13g2_fill_1 FILLER_10_257 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_fill_1 FILLER_10_329 ();
 sg13g2_decap_4 FILLER_10_338 ();
 sg13g2_fill_2 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_38 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_decap_4 FILLER_11_120 ();
 sg13g2_fill_2 FILLER_11_201 ();
 sg13g2_fill_1 FILLER_11_208 ();
 sg13g2_fill_1 FILLER_11_215 ();
 sg13g2_decap_4 FILLER_11_229 ();
 sg13g2_fill_2 FILLER_11_233 ();
 sg13g2_fill_1 FILLER_11_276 ();
 sg13g2_fill_1 FILLER_11_317 ();
 sg13g2_fill_2 FILLER_11_335 ();
 sg13g2_fill_2 FILLER_11_350 ();
 sg13g2_decap_4 FILLER_11_366 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_65 ();
 sg13g2_fill_2 FILLER_12_107 ();
 sg13g2_fill_1 FILLER_12_109 ();
 sg13g2_fill_2 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_decap_4 FILLER_12_133 ();
 sg13g2_fill_2 FILLER_12_137 ();
 sg13g2_fill_2 FILLER_12_179 ();
 sg13g2_fill_1 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_254 ();
 sg13g2_fill_2 FILLER_12_288 ();
 sg13g2_fill_1 FILLER_12_290 ();
 sg13g2_decap_8 FILLER_12_320 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_48 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_92 ();
 sg13g2_fill_2 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_fill_2 FILLER_13_138 ();
 sg13g2_fill_2 FILLER_13_149 ();
 sg13g2_fill_2 FILLER_13_160 ();
 sg13g2_fill_1 FILLER_13_162 ();
 sg13g2_fill_2 FILLER_13_176 ();
 sg13g2_fill_1 FILLER_13_178 ();
 sg13g2_fill_2 FILLER_13_199 ();
 sg13g2_fill_2 FILLER_13_223 ();
 sg13g2_decap_8 FILLER_13_239 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_decap_8 FILLER_13_253 ();
 sg13g2_decap_4 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_264 ();
 sg13g2_fill_1 FILLER_13_275 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_decap_4 FILLER_13_313 ();
 sg13g2_decap_8 FILLER_13_370 ();
 sg13g2_decap_8 FILLER_13_377 ();
 sg13g2_decap_8 FILLER_13_384 ();
 sg13g2_decap_8 FILLER_13_391 ();
 sg13g2_decap_8 FILLER_13_398 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_4 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_4 ();
 sg13g2_fill_2 FILLER_14_40 ();
 sg13g2_fill_1 FILLER_14_42 ();
 sg13g2_fill_1 FILLER_14_83 ();
 sg13g2_decap_4 FILLER_14_87 ();
 sg13g2_fill_1 FILLER_14_96 ();
 sg13g2_decap_4 FILLER_14_153 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_decap_4 FILLER_14_163 ();
 sg13g2_fill_1 FILLER_14_167 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_200 ();
 sg13g2_fill_1 FILLER_14_202 ();
 sg13g2_fill_1 FILLER_14_211 ();
 sg13g2_fill_1 FILLER_14_253 ();
 sg13g2_decap_4 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_288 ();
 sg13g2_decap_4 FILLER_14_314 ();
 sg13g2_fill_1 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_8 FILLER_14_384 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_fill_2 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_71 ();
 sg13g2_decap_4 FILLER_15_81 ();
 sg13g2_fill_2 FILLER_15_85 ();
 sg13g2_decap_4 FILLER_15_96 ();
 sg13g2_fill_2 FILLER_15_100 ();
 sg13g2_fill_2 FILLER_15_107 ();
 sg13g2_decap_8 FILLER_15_155 ();
 sg13g2_fill_1 FILLER_15_162 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_fill_2 FILLER_15_200 ();
 sg13g2_decap_4 FILLER_15_205 ();
 sg13g2_fill_1 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_222 ();
 sg13g2_decap_8 FILLER_15_229 ();
 sg13g2_decap_8 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_15_243 ();
 sg13g2_decap_4 FILLER_15_250 ();
 sg13g2_fill_2 FILLER_15_268 ();
 sg13g2_fill_1 FILLER_15_270 ();
 sg13g2_fill_2 FILLER_15_318 ();
 sg13g2_decap_4 FILLER_15_329 ();
 sg13g2_fill_1 FILLER_15_333 ();
 sg13g2_fill_2 FILLER_15_346 ();
 sg13g2_fill_1 FILLER_15_348 ();
 sg13g2_decap_4 FILLER_15_358 ();
 sg13g2_fill_1 FILLER_15_362 ();
 sg13g2_fill_2 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_55 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_4 FILLER_16_74 ();
 sg13g2_fill_1 FILLER_16_78 ();
 sg13g2_fill_1 FILLER_16_114 ();
 sg13g2_fill_1 FILLER_16_128 ();
 sg13g2_decap_8 FILLER_16_157 ();
 sg13g2_fill_2 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_1 FILLER_16_202 ();
 sg13g2_decap_4 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_296 ();
 sg13g2_fill_1 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_fill_2 FILLER_16_357 ();
 sg13g2_fill_1 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_4 ();
 sg13g2_fill_2 FILLER_17_19 ();
 sg13g2_fill_1 FILLER_17_21 ();
 sg13g2_decap_4 FILLER_17_41 ();
 sg13g2_decap_8 FILLER_17_54 ();
 sg13g2_fill_2 FILLER_17_61 ();
 sg13g2_fill_2 FILLER_17_68 ();
 sg13g2_decap_4 FILLER_17_148 ();
 sg13g2_fill_2 FILLER_17_152 ();
 sg13g2_fill_2 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_240 ();
 sg13g2_decap_4 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_4 FILLER_17_343 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_43 ();
 sg13g2_fill_1 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_107 ();
 sg13g2_decap_8 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_fill_2 FILLER_18_174 ();
 sg13g2_decap_8 FILLER_18_187 ();
 sg13g2_decap_8 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_201 ();
 sg13g2_fill_1 FILLER_18_219 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_fill_2 FILLER_18_255 ();
 sg13g2_fill_1 FILLER_18_257 ();
 sg13g2_decap_4 FILLER_18_285 ();
 sg13g2_fill_2 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_decap_4 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_331 ();
 sg13g2_fill_2 FILLER_18_372 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_7 ();
 sg13g2_fill_2 FILLER_19_11 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_fill_1 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_4 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_decap_4 FILLER_19_224 ();
 sg13g2_fill_1 FILLER_19_237 ();
 sg13g2_decap_4 FILLER_19_251 ();
 sg13g2_fill_2 FILLER_19_255 ();
 sg13g2_decap_4 FILLER_19_292 ();
 sg13g2_fill_1 FILLER_19_296 ();
 sg13g2_fill_2 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_313 ();
 sg13g2_decap_8 FILLER_19_320 ();
 sg13g2_fill_2 FILLER_19_327 ();
 sg13g2_fill_1 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_397 ();
 sg13g2_fill_1 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_13 ();
 sg13g2_decap_4 FILLER_20_57 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_184 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_fill_2 FILLER_20_228 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_fill_2 FILLER_20_346 ();
 sg13g2_fill_1 FILLER_20_348 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_1 FILLER_21_57 ();
 sg13g2_fill_1 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_98 ();
 sg13g2_fill_2 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_202 ();
 sg13g2_decap_4 FILLER_21_216 ();
 sg13g2_decap_4 FILLER_21_233 ();
 sg13g2_fill_1 FILLER_21_237 ();
 sg13g2_fill_2 FILLER_21_292 ();
 sg13g2_fill_2 FILLER_21_326 ();
 sg13g2_decap_4 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_362 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_152 ();
 sg13g2_fill_2 FILLER_22_178 ();
 sg13g2_decap_4 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_274 ();
 sg13g2_decap_4 FILLER_22_349 ();
 sg13g2_fill_2 FILLER_22_353 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_97 ();
 sg13g2_fill_1 FILLER_23_99 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_2 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_fill_2 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_fill_2 FILLER_23_288 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_364 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_fill_2 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_41 ();
 sg13g2_fill_1 FILLER_24_43 ();
 sg13g2_decap_8 FILLER_24_48 ();
 sg13g2_decap_4 FILLER_24_55 ();
 sg13g2_fill_2 FILLER_24_64 ();
 sg13g2_fill_2 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_98 ();
 sg13g2_fill_1 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_fill_2 FILLER_24_221 ();
 sg13g2_decap_4 FILLER_24_272 ();
 sg13g2_fill_2 FILLER_24_276 ();
 sg13g2_fill_1 FILLER_24_344 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_decap_4 FILLER_25_43 ();
 sg13g2_fill_2 FILLER_25_47 ();
 sg13g2_decap_4 FILLER_25_58 ();
 sg13g2_fill_2 FILLER_25_62 ();
 sg13g2_decap_4 FILLER_25_90 ();
 sg13g2_decap_4 FILLER_25_99 ();
 sg13g2_fill_1 FILLER_25_110 ();
 sg13g2_fill_2 FILLER_25_126 ();
 sg13g2_fill_2 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_190 ();
 sg13g2_fill_2 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_211 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_decap_4 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_287 ();
 sg13g2_fill_2 FILLER_25_350 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_decap_4 FILLER_26_60 ();
 sg13g2_fill_1 FILLER_26_64 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_fill_2 FILLER_26_111 ();
 sg13g2_fill_1 FILLER_26_113 ();
 sg13g2_decap_4 FILLER_26_149 ();
 sg13g2_fill_2 FILLER_26_173 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_decap_4 FILLER_26_215 ();
 sg13g2_fill_2 FILLER_26_219 ();
 sg13g2_fill_1 FILLER_26_252 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_fill_1 FILLER_26_340 ();
 sg13g2_fill_1 FILLER_26_358 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_fill_1 FILLER_26_401 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_fill_2 FILLER_27_62 ();
 sg13g2_fill_1 FILLER_27_64 ();
 sg13g2_fill_2 FILLER_27_92 ();
 sg13g2_decap_4 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_120 ();
 sg13g2_fill_2 FILLER_27_134 ();
 sg13g2_fill_2 FILLER_27_163 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_fill_2 FILLER_27_221 ();
 sg13g2_fill_1 FILLER_27_249 ();
 sg13g2_fill_1 FILLER_27_351 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_44 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_decap_4 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_166 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_fill_2 FILLER_28_231 ();
 sg13g2_fill_1 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_268 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_48 ();
 sg13g2_decap_8 FILLER_29_55 ();
 sg13g2_fill_1 FILLER_29_62 ();
 sg13g2_fill_1 FILLER_29_73 ();
 sg13g2_fill_2 FILLER_29_120 ();
 sg13g2_decap_4 FILLER_29_153 ();
 sg13g2_decap_8 FILLER_29_170 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_29_203 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_4 FILLER_29_223 ();
 sg13g2_fill_2 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_259 ();
 sg13g2_fill_2 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_306 ();
 sg13g2_fill_1 FILLER_29_354 ();
 sg13g2_fill_2 FILLER_29_392 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_48 ();
 sg13g2_decap_8 FILLER_30_55 ();
 sg13g2_fill_1 FILLER_30_62 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_44 ();
 sg13g2_fill_2 FILLER_31_51 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_17 ();
 sg13g2_fill_1 FILLER_32_19 ();
 sg13g2_decap_8 FILLER_32_48 ();
 sg13g2_fill_2 FILLER_32_55 ();
 sg13g2_fill_1 FILLER_32_57 ();
 sg13g2_fill_2 FILLER_32_99 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_fill_2 FILLER_32_134 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_167 ();
 sg13g2_decap_4 FILLER_32_174 ();
 sg13g2_fill_2 FILLER_32_205 ();
 sg13g2_fill_1 FILLER_32_221 ();
 sg13g2_fill_1 FILLER_32_301 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_2 ();
 sg13g2_decap_4 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_86 ();
 sg13g2_decap_8 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_decap_4 FILLER_33_165 ();
 sg13g2_fill_2 FILLER_33_185 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_213 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_299 ();
 sg13g2_fill_1 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_350 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_2 FILLER_34_11 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_87 ();
 sg13g2_decap_4 FILLER_34_111 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_2 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_decap_8 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_259 ();
 sg13g2_decap_8 FILLER_34_266 ();
 sg13g2_fill_1 FILLER_34_278 ();
 sg13g2_fill_1 FILLER_34_287 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_fill_1 FILLER_35_23 ();
 sg13g2_fill_2 FILLER_35_51 ();
 sg13g2_fill_2 FILLER_35_138 ();
 sg13g2_fill_1 FILLER_35_140 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_decap_4 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_298 ();
 sg13g2_fill_2 FILLER_35_320 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_28 ();
 sg13g2_fill_2 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_53 ();
 sg13g2_decap_4 FILLER_36_210 ();
 sg13g2_fill_2 FILLER_36_254 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_fill_2 FILLER_36_363 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_fill_2 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_40 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_fill_2 FILLER_37_153 ();
 sg13g2_fill_1 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_1 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_177 ();
 sg13g2_fill_1 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_267 ();
 sg13g2_fill_1 FILLER_37_296 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_fill_2 FILLER_38_71 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_134 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_212 ();
 sg13g2_fill_1 FILLER_38_214 ();
 sg13g2_decap_4 FILLER_38_238 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_fill_2 FILLER_38_277 ();
 sg13g2_fill_1 FILLER_38_279 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_fill_1 FILLER_38_347 ();
 assign uio_oe[0] = net4;
 assign uio_oe[1] = net5;
 assign uio_oe[2] = net6;
 assign uio_oe[3] = net7;
 assign uio_oe[4] = net8;
 assign uio_oe[5] = net9;
 assign uio_oe[6] = net10;
 assign uio_oe[7] = net11;
 assign uio_out[0] = net12;
 assign uio_out[1] = net13;
 assign uio_out[2] = net14;
 assign uio_out[3] = net15;
 assign uio_out[4] = net16;
 assign uio_out[5] = net17;
 assign uio_out[6] = net18;
 assign uio_out[7] = net19;
endmodule
