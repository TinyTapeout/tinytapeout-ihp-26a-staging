module tt_um_ygdes_hdsiso8 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire CLK_OUT;
 wire DL_out;
 wire \Decoded8[0] ;
 wire \Decoded8[1] ;
 wire \Decoded8[2] ;
 wire \Decoded8[3] ;
 wire \Decoded8[4] ;
 wire \Decoded8[5] ;
 wire \Decoded8[6] ;
 wire \Decoded8[7] ;
 wire INT_RESET;
 wire \J8.DecN[0] ;
 wire \J8.DecN[1] ;
 wire \J8.DecN[2] ;
 wire \J8.DecN[3] ;
 wire \J8.DecN[4] ;
 wire \J8.DecN[5] ;
 wire \J8.DecN[6] ;
 wire \J8.DecN[7] ;
 wire \J8.J4N[0] ;
 wire \J8.J4N[1] ;
 wire \J8.J4N[2] ;
 wire \J8.J4N[3] ;
 wire \J8.rst ;
 wire \J8.rst1 ;
 wire \J8.rst2 ;
 wire \J8.rst3 ;
 wire LFSR_BIT;
 wire LFSR_PERIOD;
 wire \LFSR_state8[1] ;
 wire \LFSR_state8[2] ;
 wire \LFSR_state8[3] ;
 wire \LFSR_state8[4] ;
 wire \LFSR_state8[5] ;
 wire \LFSR_state8[6] ;
 wire \LFSR_state8[7] ;
 wire MX_out;
 wire SISO_in;
 wire back;
 wire \chain4[0] ;
 wire \chain4[1] ;
 wire \chain4[2] ;
 wire \chain4[3] ;
 wire \lfsr.and8_1 ;
 wire \lfsr.and8_2 ;
 wire \lfsr.dum1 ;
 wire \lfsr.dum2 ;
 wire \lfsr.feedback ;
 wire \lfsr.x1 ;
 wire \lfsr.x2 ;
 wire \lfsr.x3 ;
 wire \siso256_1.Amp0.Y[0] ;
 wire \siso256_1.Amp0.Y[1] ;
 wire \siso256_1.Amp0.Y[2] ;
 wire \siso256_1.Amp0.Y[3] ;
 wire \siso256_1.Amp1.Y[0] ;
 wire \siso256_1.Amp1.Y[1] ;
 wire \siso256_1.Amp1.Y[2] ;
 wire \siso256_1.Amp1.Y[3] ;
 wire \siso256_1.Amp2.Y[0] ;
 wire \siso256_1.Amp2.Y[1] ;
 wire \siso256_1.Amp2.Y[2] ;
 wire \siso256_1.Amp2.Y[3] ;
 wire \siso256_1.Amp3.Y[0] ;
 wire \siso256_1.Amp3.Y[1] ;
 wire \siso256_1.Amp3.Y[2] ;
 wire \siso256_1.Amp3.Y[3] ;
 wire \siso256_1.Amp4.Y[0] ;
 wire \siso256_1.Amp4.Y[1] ;
 wire \siso256_1.Amp4.Y[2] ;
 wire \siso256_1.Amp4.Y[3] ;
 wire \siso256_1.siso_in[1] ;
 wire \siso256_1.siso_in[3] ;
 wire \siso256_1.t1[0] ;
 wire \siso256_1.t1[1] ;
 wire \siso256_1.t1[2] ;
 wire \siso256_1.t1[3] ;
 wire \siso256_1.t2[0] ;
 wire \siso256_1.t2[1] ;
 wire \siso256_1.t2[2] ;
 wire \siso256_1.t2[3] ;
 wire \siso256_1.t3[0] ;
 wire \siso256_1.t3[1] ;
 wire \siso256_1.t3[2] ;
 wire \siso256_1.t3[3] ;
 wire \siso256_1.tranche0.t1[0] ;
 wire \siso256_1.tranche0.t1[1] ;
 wire \siso256_1.tranche0.t1[2] ;
 wire \siso256_1.tranche0.t1[3] ;
 wire \siso256_1.tranche0.t2[0] ;
 wire \siso256_1.tranche0.t2[1] ;
 wire \siso256_1.tranche0.t2[2] ;
 wire \siso256_1.tranche0.t2[3] ;
 wire \siso256_1.tranche0.t3[0] ;
 wire \siso256_1.tranche0.t3[1] ;
 wire \siso256_1.tranche0.t3[2] ;
 wire \siso256_1.tranche0.t3[3] ;
 wire \siso256_1.tranche0.tranche0.slice0.latch ;
 wire \siso256_1.tranche0.tranche0.slice0.latch_n ;
 wire \siso256_1.tranche0.tranche0.slice0.siso_out[0] ;
 wire \siso256_1.tranche0.tranche0.slice0.siso_out[1] ;
 wire \siso256_1.tranche0.tranche0.slice0.siso_out[2] ;
 wire \siso256_1.tranche0.tranche0.slice0.siso_out[3] ;
 wire \siso256_1.tranche0.tranche0.slice1.latch ;
 wire \siso256_1.tranche0.tranche0.slice1.latch_n ;
 wire \siso256_1.tranche0.tranche0.slice1.siso_out[0] ;
 wire \siso256_1.tranche0.tranche0.slice1.siso_out[1] ;
 wire \siso256_1.tranche0.tranche0.slice1.siso_out[2] ;
 wire \siso256_1.tranche0.tranche0.slice1.siso_out[3] ;
 wire \siso256_1.tranche0.tranche0.slice2.latch ;
 wire \siso256_1.tranche0.tranche0.slice2.latch_n ;
 wire \siso256_1.tranche0.tranche0.slice2.siso_out[0] ;
 wire \siso256_1.tranche0.tranche0.slice2.siso_out[1] ;
 wire \siso256_1.tranche0.tranche0.slice2.siso_out[2] ;
 wire \siso256_1.tranche0.tranche0.slice2.siso_out[3] ;
 wire \siso256_1.tranche0.tranche0.slice3.latch ;
 wire \siso256_1.tranche0.tranche0.slice3.latch_n ;
 wire \siso256_1.tranche0.tranche1.slice0.latch_n ;
 wire \siso256_1.tranche0.tranche1.slice0.siso_out[0] ;
 wire \siso256_1.tranche0.tranche1.slice0.siso_out[1] ;
 wire \siso256_1.tranche0.tranche1.slice0.siso_out[2] ;
 wire \siso256_1.tranche0.tranche1.slice0.siso_out[3] ;
 wire \siso256_1.tranche0.tranche1.slice1.latch_n ;
 wire \siso256_1.tranche0.tranche1.slice1.siso_out[0] ;
 wire \siso256_1.tranche0.tranche1.slice1.siso_out[1] ;
 wire \siso256_1.tranche0.tranche1.slice1.siso_out[2] ;
 wire \siso256_1.tranche0.tranche1.slice1.siso_out[3] ;
 wire \siso256_1.tranche0.tranche1.slice2.latch_n ;
 wire \siso256_1.tranche0.tranche1.slice2.siso_out[0] ;
 wire \siso256_1.tranche0.tranche1.slice2.siso_out[1] ;
 wire \siso256_1.tranche0.tranche1.slice2.siso_out[2] ;
 wire \siso256_1.tranche0.tranche1.slice2.siso_out[3] ;
 wire \siso256_1.tranche0.tranche1.slice3.latch_n ;
 wire \siso256_1.tranche0.tranche2.slice0.latch_n ;
 wire \siso256_1.tranche0.tranche2.slice0.siso_out[0] ;
 wire \siso256_1.tranche0.tranche2.slice0.siso_out[1] ;
 wire \siso256_1.tranche0.tranche2.slice0.siso_out[2] ;
 wire \siso256_1.tranche0.tranche2.slice0.siso_out[3] ;
 wire \siso256_1.tranche0.tranche2.slice1.latch_n ;
 wire \siso256_1.tranche0.tranche2.slice1.siso_out[0] ;
 wire \siso256_1.tranche0.tranche2.slice1.siso_out[1] ;
 wire \siso256_1.tranche0.tranche2.slice1.siso_out[2] ;
 wire \siso256_1.tranche0.tranche2.slice1.siso_out[3] ;
 wire \siso256_1.tranche0.tranche2.slice2.latch_n ;
 wire \siso256_1.tranche0.tranche2.slice2.siso_out[0] ;
 wire \siso256_1.tranche0.tranche2.slice2.siso_out[1] ;
 wire \siso256_1.tranche0.tranche2.slice2.siso_out[2] ;
 wire \siso256_1.tranche0.tranche2.slice2.siso_out[3] ;
 wire \siso256_1.tranche0.tranche2.slice3.latch_n ;
 wire \siso256_1.tranche0.tranche3.slice0.latch_n ;
 wire \siso256_1.tranche0.tranche3.slice0.siso_out[0] ;
 wire \siso256_1.tranche0.tranche3.slice0.siso_out[1] ;
 wire \siso256_1.tranche0.tranche3.slice0.siso_out[2] ;
 wire \siso256_1.tranche0.tranche3.slice0.siso_out[3] ;
 wire \siso256_1.tranche0.tranche3.slice1.latch_n ;
 wire \siso256_1.tranche0.tranche3.slice1.siso_out[0] ;
 wire \siso256_1.tranche0.tranche3.slice1.siso_out[1] ;
 wire \siso256_1.tranche0.tranche3.slice1.siso_out[2] ;
 wire \siso256_1.tranche0.tranche3.slice1.siso_out[3] ;
 wire \siso256_1.tranche0.tranche3.slice2.latch_n ;
 wire \siso256_1.tranche0.tranche3.slice2.siso_out[0] ;
 wire \siso256_1.tranche0.tranche3.slice2.siso_out[1] ;
 wire \siso256_1.tranche0.tranche3.slice2.siso_out[2] ;
 wire \siso256_1.tranche0.tranche3.slice2.siso_out[3] ;
 wire \siso256_1.tranche0.tranche3.slice3.latch_n ;
 wire \siso256_1.tranche1.t1[0] ;
 wire \siso256_1.tranche1.t1[1] ;
 wire \siso256_1.tranche1.t1[2] ;
 wire \siso256_1.tranche1.t1[3] ;
 wire \siso256_1.tranche1.t2[0] ;
 wire \siso256_1.tranche1.t2[1] ;
 wire \siso256_1.tranche1.t2[2] ;
 wire \siso256_1.tranche1.t2[3] ;
 wire \siso256_1.tranche1.t3[0] ;
 wire \siso256_1.tranche1.t3[1] ;
 wire \siso256_1.tranche1.t3[2] ;
 wire \siso256_1.tranche1.t3[3] ;
 wire \siso256_1.tranche1.tranche0.slice0.latch ;
 wire \siso256_1.tranche1.tranche0.slice0.latch_n ;
 wire \siso256_1.tranche1.tranche0.slice0.siso_out[0] ;
 wire \siso256_1.tranche1.tranche0.slice0.siso_out[1] ;
 wire \siso256_1.tranche1.tranche0.slice0.siso_out[2] ;
 wire \siso256_1.tranche1.tranche0.slice0.siso_out[3] ;
 wire \siso256_1.tranche1.tranche0.slice1.latch ;
 wire \siso256_1.tranche1.tranche0.slice1.latch_n ;
 wire \siso256_1.tranche1.tranche0.slice1.siso_out[0] ;
 wire \siso256_1.tranche1.tranche0.slice1.siso_out[1] ;
 wire \siso256_1.tranche1.tranche0.slice1.siso_out[2] ;
 wire \siso256_1.tranche1.tranche0.slice1.siso_out[3] ;
 wire \siso256_1.tranche1.tranche0.slice2.latch ;
 wire \siso256_1.tranche1.tranche0.slice2.latch_n ;
 wire \siso256_1.tranche1.tranche0.slice2.siso_out[0] ;
 wire \siso256_1.tranche1.tranche0.slice2.siso_out[1] ;
 wire \siso256_1.tranche1.tranche0.slice2.siso_out[2] ;
 wire \siso256_1.tranche1.tranche0.slice2.siso_out[3] ;
 wire \siso256_1.tranche1.tranche0.slice3.latch ;
 wire \siso256_1.tranche1.tranche0.slice3.latch_n ;
 wire \siso256_1.tranche1.tranche1.slice0.latch_n ;
 wire \siso256_1.tranche1.tranche1.slice0.siso_out[0] ;
 wire \siso256_1.tranche1.tranche1.slice0.siso_out[1] ;
 wire \siso256_1.tranche1.tranche1.slice0.siso_out[2] ;
 wire \siso256_1.tranche1.tranche1.slice0.siso_out[3] ;
 wire \siso256_1.tranche1.tranche1.slice1.latch_n ;
 wire \siso256_1.tranche1.tranche1.slice1.siso_out[0] ;
 wire \siso256_1.tranche1.tranche1.slice1.siso_out[1] ;
 wire \siso256_1.tranche1.tranche1.slice1.siso_out[2] ;
 wire \siso256_1.tranche1.tranche1.slice1.siso_out[3] ;
 wire \siso256_1.tranche1.tranche1.slice2.latch_n ;
 wire \siso256_1.tranche1.tranche1.slice2.siso_out[0] ;
 wire \siso256_1.tranche1.tranche1.slice2.siso_out[1] ;
 wire \siso256_1.tranche1.tranche1.slice2.siso_out[2] ;
 wire \siso256_1.tranche1.tranche1.slice2.siso_out[3] ;
 wire \siso256_1.tranche1.tranche1.slice3.latch_n ;
 wire \siso256_1.tranche1.tranche2.slice0.latch_n ;
 wire \siso256_1.tranche1.tranche2.slice0.siso_out[0] ;
 wire \siso256_1.tranche1.tranche2.slice0.siso_out[1] ;
 wire \siso256_1.tranche1.tranche2.slice0.siso_out[2] ;
 wire \siso256_1.tranche1.tranche2.slice0.siso_out[3] ;
 wire \siso256_1.tranche1.tranche2.slice1.latch_n ;
 wire \siso256_1.tranche1.tranche2.slice1.siso_out[0] ;
 wire \siso256_1.tranche1.tranche2.slice1.siso_out[1] ;
 wire \siso256_1.tranche1.tranche2.slice1.siso_out[2] ;
 wire \siso256_1.tranche1.tranche2.slice1.siso_out[3] ;
 wire \siso256_1.tranche1.tranche2.slice2.latch_n ;
 wire \siso256_1.tranche1.tranche2.slice2.siso_out[0] ;
 wire \siso256_1.tranche1.tranche2.slice2.siso_out[1] ;
 wire \siso256_1.tranche1.tranche2.slice2.siso_out[2] ;
 wire \siso256_1.tranche1.tranche2.slice2.siso_out[3] ;
 wire \siso256_1.tranche1.tranche2.slice3.latch_n ;
 wire \siso256_1.tranche1.tranche3.slice0.latch_n ;
 wire \siso256_1.tranche1.tranche3.slice0.siso_out[0] ;
 wire \siso256_1.tranche1.tranche3.slice0.siso_out[1] ;
 wire \siso256_1.tranche1.tranche3.slice0.siso_out[2] ;
 wire \siso256_1.tranche1.tranche3.slice0.siso_out[3] ;
 wire \siso256_1.tranche1.tranche3.slice1.latch_n ;
 wire \siso256_1.tranche1.tranche3.slice1.siso_out[0] ;
 wire \siso256_1.tranche1.tranche3.slice1.siso_out[1] ;
 wire \siso256_1.tranche1.tranche3.slice1.siso_out[2] ;
 wire \siso256_1.tranche1.tranche3.slice1.siso_out[3] ;
 wire \siso256_1.tranche1.tranche3.slice2.latch_n ;
 wire \siso256_1.tranche1.tranche3.slice2.siso_out[0] ;
 wire \siso256_1.tranche1.tranche3.slice2.siso_out[1] ;
 wire \siso256_1.tranche1.tranche3.slice2.siso_out[2] ;
 wire \siso256_1.tranche1.tranche3.slice2.siso_out[3] ;
 wire \siso256_1.tranche1.tranche3.slice3.latch_n ;
 wire \siso256_1.tranche2.t1[0] ;
 wire \siso256_1.tranche2.t1[1] ;
 wire \siso256_1.tranche2.t1[2] ;
 wire \siso256_1.tranche2.t1[3] ;
 wire \siso256_1.tranche2.t2[0] ;
 wire \siso256_1.tranche2.t2[1] ;
 wire \siso256_1.tranche2.t2[2] ;
 wire \siso256_1.tranche2.t2[3] ;
 wire \siso256_1.tranche2.t3[0] ;
 wire \siso256_1.tranche2.t3[1] ;
 wire \siso256_1.tranche2.t3[2] ;
 wire \siso256_1.tranche2.t3[3] ;
 wire \siso256_1.tranche2.tranche0.slice0.latch ;
 wire \siso256_1.tranche2.tranche0.slice0.latch_n ;
 wire \siso256_1.tranche2.tranche0.slice0.siso_out[0] ;
 wire \siso256_1.tranche2.tranche0.slice0.siso_out[1] ;
 wire \siso256_1.tranche2.tranche0.slice0.siso_out[2] ;
 wire \siso256_1.tranche2.tranche0.slice0.siso_out[3] ;
 wire \siso256_1.tranche2.tranche0.slice1.latch ;
 wire \siso256_1.tranche2.tranche0.slice1.latch_n ;
 wire \siso256_1.tranche2.tranche0.slice1.siso_out[0] ;
 wire \siso256_1.tranche2.tranche0.slice1.siso_out[1] ;
 wire \siso256_1.tranche2.tranche0.slice1.siso_out[2] ;
 wire \siso256_1.tranche2.tranche0.slice1.siso_out[3] ;
 wire \siso256_1.tranche2.tranche0.slice2.latch ;
 wire \siso256_1.tranche2.tranche0.slice2.latch_n ;
 wire \siso256_1.tranche2.tranche0.slice2.siso_out[0] ;
 wire \siso256_1.tranche2.tranche0.slice2.siso_out[1] ;
 wire \siso256_1.tranche2.tranche0.slice2.siso_out[2] ;
 wire \siso256_1.tranche2.tranche0.slice2.siso_out[3] ;
 wire \siso256_1.tranche2.tranche0.slice3.latch ;
 wire \siso256_1.tranche2.tranche0.slice3.latch_n ;
 wire \siso256_1.tranche2.tranche1.slice0.latch_n ;
 wire \siso256_1.tranche2.tranche1.slice0.siso_out[0] ;
 wire \siso256_1.tranche2.tranche1.slice0.siso_out[1] ;
 wire \siso256_1.tranche2.tranche1.slice0.siso_out[2] ;
 wire \siso256_1.tranche2.tranche1.slice0.siso_out[3] ;
 wire \siso256_1.tranche2.tranche1.slice1.latch_n ;
 wire \siso256_1.tranche2.tranche1.slice1.siso_out[0] ;
 wire \siso256_1.tranche2.tranche1.slice1.siso_out[1] ;
 wire \siso256_1.tranche2.tranche1.slice1.siso_out[2] ;
 wire \siso256_1.tranche2.tranche1.slice1.siso_out[3] ;
 wire \siso256_1.tranche2.tranche1.slice2.latch_n ;
 wire \siso256_1.tranche2.tranche1.slice2.siso_out[0] ;
 wire \siso256_1.tranche2.tranche1.slice2.siso_out[1] ;
 wire \siso256_1.tranche2.tranche1.slice2.siso_out[2] ;
 wire \siso256_1.tranche2.tranche1.slice2.siso_out[3] ;
 wire \siso256_1.tranche2.tranche1.slice3.latch_n ;
 wire \siso256_1.tranche2.tranche2.slice0.latch_n ;
 wire \siso256_1.tranche2.tranche2.slice0.siso_out[0] ;
 wire \siso256_1.tranche2.tranche2.slice0.siso_out[1] ;
 wire \siso256_1.tranche2.tranche2.slice0.siso_out[2] ;
 wire \siso256_1.tranche2.tranche2.slice0.siso_out[3] ;
 wire \siso256_1.tranche2.tranche2.slice1.latch_n ;
 wire \siso256_1.tranche2.tranche2.slice1.siso_out[0] ;
 wire \siso256_1.tranche2.tranche2.slice1.siso_out[1] ;
 wire \siso256_1.tranche2.tranche2.slice1.siso_out[2] ;
 wire \siso256_1.tranche2.tranche2.slice1.siso_out[3] ;
 wire \siso256_1.tranche2.tranche2.slice2.latch_n ;
 wire \siso256_1.tranche2.tranche2.slice2.siso_out[0] ;
 wire \siso256_1.tranche2.tranche2.slice2.siso_out[1] ;
 wire \siso256_1.tranche2.tranche2.slice2.siso_out[2] ;
 wire \siso256_1.tranche2.tranche2.slice2.siso_out[3] ;
 wire \siso256_1.tranche2.tranche2.slice3.latch_n ;
 wire \siso256_1.tranche2.tranche3.slice0.latch_n ;
 wire \siso256_1.tranche2.tranche3.slice0.siso_out[0] ;
 wire \siso256_1.tranche2.tranche3.slice0.siso_out[1] ;
 wire \siso256_1.tranche2.tranche3.slice0.siso_out[2] ;
 wire \siso256_1.tranche2.tranche3.slice0.siso_out[3] ;
 wire \siso256_1.tranche2.tranche3.slice1.latch_n ;
 wire \siso256_1.tranche2.tranche3.slice1.siso_out[0] ;
 wire \siso256_1.tranche2.tranche3.slice1.siso_out[1] ;
 wire \siso256_1.tranche2.tranche3.slice1.siso_out[2] ;
 wire \siso256_1.tranche2.tranche3.slice1.siso_out[3] ;
 wire \siso256_1.tranche2.tranche3.slice2.latch_n ;
 wire \siso256_1.tranche2.tranche3.slice2.siso_out[0] ;
 wire \siso256_1.tranche2.tranche3.slice2.siso_out[1] ;
 wire \siso256_1.tranche2.tranche3.slice2.siso_out[2] ;
 wire \siso256_1.tranche2.tranche3.slice2.siso_out[3] ;
 wire \siso256_1.tranche2.tranche3.slice3.latch_n ;
 wire \siso256_1.tranche3.t1[0] ;
 wire \siso256_1.tranche3.t1[1] ;
 wire \siso256_1.tranche3.t1[2] ;
 wire \siso256_1.tranche3.t1[3] ;
 wire \siso256_1.tranche3.t2[0] ;
 wire \siso256_1.tranche3.t2[1] ;
 wire \siso256_1.tranche3.t2[2] ;
 wire \siso256_1.tranche3.t2[3] ;
 wire \siso256_1.tranche3.t3[0] ;
 wire \siso256_1.tranche3.t3[1] ;
 wire \siso256_1.tranche3.t3[2] ;
 wire \siso256_1.tranche3.t3[3] ;
 wire \siso256_1.tranche3.tranche0.slice0.latch ;
 wire \siso256_1.tranche3.tranche0.slice0.latch_n ;
 wire \siso256_1.tranche3.tranche0.slice0.siso_out[0] ;
 wire \siso256_1.tranche3.tranche0.slice0.siso_out[1] ;
 wire \siso256_1.tranche3.tranche0.slice0.siso_out[2] ;
 wire \siso256_1.tranche3.tranche0.slice0.siso_out[3] ;
 wire \siso256_1.tranche3.tranche0.slice1.latch ;
 wire \siso256_1.tranche3.tranche0.slice1.latch_n ;
 wire \siso256_1.tranche3.tranche0.slice1.siso_out[0] ;
 wire \siso256_1.tranche3.tranche0.slice1.siso_out[1] ;
 wire \siso256_1.tranche3.tranche0.slice1.siso_out[2] ;
 wire \siso256_1.tranche3.tranche0.slice1.siso_out[3] ;
 wire \siso256_1.tranche3.tranche0.slice2.latch ;
 wire \siso256_1.tranche3.tranche0.slice2.latch_n ;
 wire \siso256_1.tranche3.tranche0.slice2.siso_out[0] ;
 wire \siso256_1.tranche3.tranche0.slice2.siso_out[1] ;
 wire \siso256_1.tranche3.tranche0.slice2.siso_out[2] ;
 wire \siso256_1.tranche3.tranche0.slice2.siso_out[3] ;
 wire \siso256_1.tranche3.tranche0.slice3.latch ;
 wire \siso256_1.tranche3.tranche0.slice3.latch_n ;
 wire \siso256_1.tranche3.tranche1.slice0.latch_n ;
 wire \siso256_1.tranche3.tranche1.slice0.siso_out[0] ;
 wire \siso256_1.tranche3.tranche1.slice0.siso_out[1] ;
 wire \siso256_1.tranche3.tranche1.slice0.siso_out[2] ;
 wire \siso256_1.tranche3.tranche1.slice0.siso_out[3] ;
 wire \siso256_1.tranche3.tranche1.slice1.latch_n ;
 wire \siso256_1.tranche3.tranche1.slice1.siso_out[0] ;
 wire \siso256_1.tranche3.tranche1.slice1.siso_out[1] ;
 wire \siso256_1.tranche3.tranche1.slice1.siso_out[2] ;
 wire \siso256_1.tranche3.tranche1.slice1.siso_out[3] ;
 wire \siso256_1.tranche3.tranche1.slice2.latch_n ;
 wire \siso256_1.tranche3.tranche1.slice2.siso_out[0] ;
 wire \siso256_1.tranche3.tranche1.slice2.siso_out[1] ;
 wire \siso256_1.tranche3.tranche1.slice2.siso_out[2] ;
 wire \siso256_1.tranche3.tranche1.slice2.siso_out[3] ;
 wire \siso256_1.tranche3.tranche1.slice3.latch_n ;
 wire \siso256_1.tranche3.tranche2.slice0.latch_n ;
 wire \siso256_1.tranche3.tranche2.slice0.siso_out[0] ;
 wire \siso256_1.tranche3.tranche2.slice0.siso_out[1] ;
 wire \siso256_1.tranche3.tranche2.slice0.siso_out[2] ;
 wire \siso256_1.tranche3.tranche2.slice0.siso_out[3] ;
 wire \siso256_1.tranche3.tranche2.slice1.latch_n ;
 wire \siso256_1.tranche3.tranche2.slice1.siso_out[0] ;
 wire \siso256_1.tranche3.tranche2.slice1.siso_out[1] ;
 wire \siso256_1.tranche3.tranche2.slice1.siso_out[2] ;
 wire \siso256_1.tranche3.tranche2.slice1.siso_out[3] ;
 wire \siso256_1.tranche3.tranche2.slice2.latch_n ;
 wire \siso256_1.tranche3.tranche2.slice2.siso_out[0] ;
 wire \siso256_1.tranche3.tranche2.slice2.siso_out[1] ;
 wire \siso256_1.tranche3.tranche2.slice2.siso_out[2] ;
 wire \siso256_1.tranche3.tranche2.slice2.siso_out[3] ;
 wire \siso256_1.tranche3.tranche2.slice3.latch_n ;
 wire \siso256_1.tranche3.tranche3.slice0.latch_n ;
 wire \siso256_1.tranche3.tranche3.slice0.siso_out[0] ;
 wire \siso256_1.tranche3.tranche3.slice0.siso_out[1] ;
 wire \siso256_1.tranche3.tranche3.slice0.siso_out[2] ;
 wire \siso256_1.tranche3.tranche3.slice0.siso_out[3] ;
 wire \siso256_1.tranche3.tranche3.slice1.latch_n ;
 wire \siso256_1.tranche3.tranche3.slice1.siso_out[0] ;
 wire \siso256_1.tranche3.tranche3.slice1.siso_out[1] ;
 wire \siso256_1.tranche3.tranche3.slice1.siso_out[2] ;
 wire \siso256_1.tranche3.tranche3.slice1.siso_out[3] ;
 wire \siso256_1.tranche3.tranche3.slice2.latch_n ;
 wire \siso256_1.tranche3.tranche3.slice2.siso_out[0] ;
 wire \siso256_1.tranche3.tranche3.slice2.siso_out[1] ;
 wire \siso256_1.tranche3.tranche3.slice2.siso_out[2] ;
 wire \siso256_1.tranche3.tranche3.slice2.siso_out[3] ;
 wire \siso256_1.tranche3.tranche3.slice3.latch_n ;
 wire \siso256_2.Amp0.Y[0] ;
 wire \siso256_2.Amp0.Y[1] ;
 wire \siso256_2.Amp0.Y[2] ;
 wire \siso256_2.Amp0.Y[3] ;
 wire \siso256_2.Amp1.Y[0] ;
 wire \siso256_2.Amp1.Y[1] ;
 wire \siso256_2.Amp1.Y[2] ;
 wire \siso256_2.Amp1.Y[3] ;
 wire \siso256_2.Amp2.Y[0] ;
 wire \siso256_2.Amp2.Y[1] ;
 wire \siso256_2.Amp2.Y[2] ;
 wire \siso256_2.Amp2.Y[3] ;
 wire \siso256_2.Amp3.Y[0] ;
 wire \siso256_2.Amp3.Y[1] ;
 wire \siso256_2.Amp3.Y[2] ;
 wire \siso256_2.Amp3.Y[3] ;
 wire \siso256_2.Amp4.Y[0] ;
 wire \siso256_2.Amp4.Y[1] ;
 wire \siso256_2.Amp4.Y[2] ;
 wire \siso256_2.Amp4.Y[3] ;
 wire \siso256_2.t1[0] ;
 wire \siso256_2.t1[1] ;
 wire \siso256_2.t1[2] ;
 wire \siso256_2.t1[3] ;
 wire \siso256_2.t2[0] ;
 wire \siso256_2.t2[1] ;
 wire \siso256_2.t2[2] ;
 wire \siso256_2.t2[3] ;
 wire \siso256_2.t3[0] ;
 wire \siso256_2.t3[1] ;
 wire \siso256_2.t3[2] ;
 wire \siso256_2.t3[3] ;
 wire \siso256_2.tranche0.t1[0] ;
 wire \siso256_2.tranche0.t1[1] ;
 wire \siso256_2.tranche0.t1[2] ;
 wire \siso256_2.tranche0.t1[3] ;
 wire \siso256_2.tranche0.t2[0] ;
 wire \siso256_2.tranche0.t2[1] ;
 wire \siso256_2.tranche0.t2[2] ;
 wire \siso256_2.tranche0.t2[3] ;
 wire \siso256_2.tranche0.t3[0] ;
 wire \siso256_2.tranche0.t3[1] ;
 wire \siso256_2.tranche0.t3[2] ;
 wire \siso256_2.tranche0.t3[3] ;
 wire \siso256_2.tranche0.tranche0.slice0.latch ;
 wire \siso256_2.tranche0.tranche0.slice0.latch_n ;
 wire \siso256_2.tranche0.tranche0.slice0.siso_out[0] ;
 wire \siso256_2.tranche0.tranche0.slice0.siso_out[1] ;
 wire \siso256_2.tranche0.tranche0.slice0.siso_out[2] ;
 wire \siso256_2.tranche0.tranche0.slice0.siso_out[3] ;
 wire \siso256_2.tranche0.tranche0.slice1.latch ;
 wire \siso256_2.tranche0.tranche0.slice1.latch_n ;
 wire \siso256_2.tranche0.tranche0.slice1.siso_out[0] ;
 wire \siso256_2.tranche0.tranche0.slice1.siso_out[1] ;
 wire \siso256_2.tranche0.tranche0.slice1.siso_out[2] ;
 wire \siso256_2.tranche0.tranche0.slice1.siso_out[3] ;
 wire \siso256_2.tranche0.tranche0.slice2.latch ;
 wire \siso256_2.tranche0.tranche0.slice2.latch_n ;
 wire \siso256_2.tranche0.tranche0.slice2.siso_out[0] ;
 wire \siso256_2.tranche0.tranche0.slice2.siso_out[1] ;
 wire \siso256_2.tranche0.tranche0.slice2.siso_out[2] ;
 wire \siso256_2.tranche0.tranche0.slice2.siso_out[3] ;
 wire \siso256_2.tranche0.tranche0.slice3.latch ;
 wire \siso256_2.tranche0.tranche0.slice3.latch_n ;
 wire \siso256_2.tranche0.tranche1.slice0.latch_n ;
 wire \siso256_2.tranche0.tranche1.slice0.siso_out[0] ;
 wire \siso256_2.tranche0.tranche1.slice0.siso_out[1] ;
 wire \siso256_2.tranche0.tranche1.slice0.siso_out[2] ;
 wire \siso256_2.tranche0.tranche1.slice0.siso_out[3] ;
 wire \siso256_2.tranche0.tranche1.slice1.latch_n ;
 wire \siso256_2.tranche0.tranche1.slice1.siso_out[0] ;
 wire \siso256_2.tranche0.tranche1.slice1.siso_out[1] ;
 wire \siso256_2.tranche0.tranche1.slice1.siso_out[2] ;
 wire \siso256_2.tranche0.tranche1.slice1.siso_out[3] ;
 wire \siso256_2.tranche0.tranche1.slice2.latch_n ;
 wire \siso256_2.tranche0.tranche1.slice2.siso_out[0] ;
 wire \siso256_2.tranche0.tranche1.slice2.siso_out[1] ;
 wire \siso256_2.tranche0.tranche1.slice2.siso_out[2] ;
 wire \siso256_2.tranche0.tranche1.slice2.siso_out[3] ;
 wire \siso256_2.tranche0.tranche1.slice3.latch_n ;
 wire \siso256_2.tranche0.tranche2.slice0.latch_n ;
 wire \siso256_2.tranche0.tranche2.slice0.siso_out[0] ;
 wire \siso256_2.tranche0.tranche2.slice0.siso_out[1] ;
 wire \siso256_2.tranche0.tranche2.slice0.siso_out[2] ;
 wire \siso256_2.tranche0.tranche2.slice0.siso_out[3] ;
 wire \siso256_2.tranche0.tranche2.slice1.latch_n ;
 wire \siso256_2.tranche0.tranche2.slice1.siso_out[0] ;
 wire \siso256_2.tranche0.tranche2.slice1.siso_out[1] ;
 wire \siso256_2.tranche0.tranche2.slice1.siso_out[2] ;
 wire \siso256_2.tranche0.tranche2.slice1.siso_out[3] ;
 wire \siso256_2.tranche0.tranche2.slice2.latch_n ;
 wire \siso256_2.tranche0.tranche2.slice2.siso_out[0] ;
 wire \siso256_2.tranche0.tranche2.slice2.siso_out[1] ;
 wire \siso256_2.tranche0.tranche2.slice2.siso_out[2] ;
 wire \siso256_2.tranche0.tranche2.slice2.siso_out[3] ;
 wire \siso256_2.tranche0.tranche2.slice3.latch_n ;
 wire \siso256_2.tranche0.tranche3.slice0.latch_n ;
 wire \siso256_2.tranche0.tranche3.slice0.siso_out[0] ;
 wire \siso256_2.tranche0.tranche3.slice0.siso_out[1] ;
 wire \siso256_2.tranche0.tranche3.slice0.siso_out[2] ;
 wire \siso256_2.tranche0.tranche3.slice0.siso_out[3] ;
 wire \siso256_2.tranche0.tranche3.slice1.latch_n ;
 wire \siso256_2.tranche0.tranche3.slice1.siso_out[0] ;
 wire \siso256_2.tranche0.tranche3.slice1.siso_out[1] ;
 wire \siso256_2.tranche0.tranche3.slice1.siso_out[2] ;
 wire \siso256_2.tranche0.tranche3.slice1.siso_out[3] ;
 wire \siso256_2.tranche0.tranche3.slice2.latch_n ;
 wire \siso256_2.tranche0.tranche3.slice2.siso_out[0] ;
 wire \siso256_2.tranche0.tranche3.slice2.siso_out[1] ;
 wire \siso256_2.tranche0.tranche3.slice2.siso_out[2] ;
 wire \siso256_2.tranche0.tranche3.slice2.siso_out[3] ;
 wire \siso256_2.tranche0.tranche3.slice3.latch_n ;
 wire \siso256_2.tranche1.t1[0] ;
 wire \siso256_2.tranche1.t1[1] ;
 wire \siso256_2.tranche1.t1[2] ;
 wire \siso256_2.tranche1.t1[3] ;
 wire \siso256_2.tranche1.t2[0] ;
 wire \siso256_2.tranche1.t2[1] ;
 wire \siso256_2.tranche1.t2[2] ;
 wire \siso256_2.tranche1.t2[3] ;
 wire \siso256_2.tranche1.t3[0] ;
 wire \siso256_2.tranche1.t3[1] ;
 wire \siso256_2.tranche1.t3[2] ;
 wire \siso256_2.tranche1.t3[3] ;
 wire \siso256_2.tranche1.tranche0.slice0.latch ;
 wire \siso256_2.tranche1.tranche0.slice0.latch_n ;
 wire \siso256_2.tranche1.tranche0.slice0.siso_out[0] ;
 wire \siso256_2.tranche1.tranche0.slice0.siso_out[1] ;
 wire \siso256_2.tranche1.tranche0.slice0.siso_out[2] ;
 wire \siso256_2.tranche1.tranche0.slice0.siso_out[3] ;
 wire \siso256_2.tranche1.tranche0.slice1.latch ;
 wire \siso256_2.tranche1.tranche0.slice1.latch_n ;
 wire \siso256_2.tranche1.tranche0.slice1.siso_out[0] ;
 wire \siso256_2.tranche1.tranche0.slice1.siso_out[1] ;
 wire \siso256_2.tranche1.tranche0.slice1.siso_out[2] ;
 wire \siso256_2.tranche1.tranche0.slice1.siso_out[3] ;
 wire \siso256_2.tranche1.tranche0.slice2.latch ;
 wire \siso256_2.tranche1.tranche0.slice2.latch_n ;
 wire \siso256_2.tranche1.tranche0.slice2.siso_out[0] ;
 wire \siso256_2.tranche1.tranche0.slice2.siso_out[1] ;
 wire \siso256_2.tranche1.tranche0.slice2.siso_out[2] ;
 wire \siso256_2.tranche1.tranche0.slice2.siso_out[3] ;
 wire \siso256_2.tranche1.tranche0.slice3.latch ;
 wire \siso256_2.tranche1.tranche0.slice3.latch_n ;
 wire \siso256_2.tranche1.tranche1.slice0.latch_n ;
 wire \siso256_2.tranche1.tranche1.slice0.siso_out[0] ;
 wire \siso256_2.tranche1.tranche1.slice0.siso_out[1] ;
 wire \siso256_2.tranche1.tranche1.slice0.siso_out[2] ;
 wire \siso256_2.tranche1.tranche1.slice0.siso_out[3] ;
 wire \siso256_2.tranche1.tranche1.slice1.latch_n ;
 wire \siso256_2.tranche1.tranche1.slice1.siso_out[0] ;
 wire \siso256_2.tranche1.tranche1.slice1.siso_out[1] ;
 wire \siso256_2.tranche1.tranche1.slice1.siso_out[2] ;
 wire \siso256_2.tranche1.tranche1.slice1.siso_out[3] ;
 wire \siso256_2.tranche1.tranche1.slice2.latch_n ;
 wire \siso256_2.tranche1.tranche1.slice2.siso_out[0] ;
 wire \siso256_2.tranche1.tranche1.slice2.siso_out[1] ;
 wire \siso256_2.tranche1.tranche1.slice2.siso_out[2] ;
 wire \siso256_2.tranche1.tranche1.slice2.siso_out[3] ;
 wire \siso256_2.tranche1.tranche1.slice3.latch_n ;
 wire \siso256_2.tranche1.tranche2.slice0.latch_n ;
 wire \siso256_2.tranche1.tranche2.slice0.siso_out[0] ;
 wire \siso256_2.tranche1.tranche2.slice0.siso_out[1] ;
 wire \siso256_2.tranche1.tranche2.slice0.siso_out[2] ;
 wire \siso256_2.tranche1.tranche2.slice0.siso_out[3] ;
 wire \siso256_2.tranche1.tranche2.slice1.latch_n ;
 wire \siso256_2.tranche1.tranche2.slice1.siso_out[0] ;
 wire \siso256_2.tranche1.tranche2.slice1.siso_out[1] ;
 wire \siso256_2.tranche1.tranche2.slice1.siso_out[2] ;
 wire \siso256_2.tranche1.tranche2.slice1.siso_out[3] ;
 wire \siso256_2.tranche1.tranche2.slice2.latch_n ;
 wire \siso256_2.tranche1.tranche2.slice2.siso_out[0] ;
 wire \siso256_2.tranche1.tranche2.slice2.siso_out[1] ;
 wire \siso256_2.tranche1.tranche2.slice2.siso_out[2] ;
 wire \siso256_2.tranche1.tranche2.slice2.siso_out[3] ;
 wire \siso256_2.tranche1.tranche2.slice3.latch_n ;
 wire \siso256_2.tranche1.tranche3.slice0.latch_n ;
 wire \siso256_2.tranche1.tranche3.slice0.siso_out[0] ;
 wire \siso256_2.tranche1.tranche3.slice0.siso_out[1] ;
 wire \siso256_2.tranche1.tranche3.slice0.siso_out[2] ;
 wire \siso256_2.tranche1.tranche3.slice0.siso_out[3] ;
 wire \siso256_2.tranche1.tranche3.slice1.latch_n ;
 wire \siso256_2.tranche1.tranche3.slice1.siso_out[0] ;
 wire \siso256_2.tranche1.tranche3.slice1.siso_out[1] ;
 wire \siso256_2.tranche1.tranche3.slice1.siso_out[2] ;
 wire \siso256_2.tranche1.tranche3.slice1.siso_out[3] ;
 wire \siso256_2.tranche1.tranche3.slice2.latch_n ;
 wire \siso256_2.tranche1.tranche3.slice2.siso_out[0] ;
 wire \siso256_2.tranche1.tranche3.slice2.siso_out[1] ;
 wire \siso256_2.tranche1.tranche3.slice2.siso_out[2] ;
 wire \siso256_2.tranche1.tranche3.slice2.siso_out[3] ;
 wire \siso256_2.tranche1.tranche3.slice3.latch_n ;
 wire \siso256_2.tranche2.t1[0] ;
 wire \siso256_2.tranche2.t1[1] ;
 wire \siso256_2.tranche2.t1[2] ;
 wire \siso256_2.tranche2.t1[3] ;
 wire \siso256_2.tranche2.t2[0] ;
 wire \siso256_2.tranche2.t2[1] ;
 wire \siso256_2.tranche2.t2[2] ;
 wire \siso256_2.tranche2.t2[3] ;
 wire \siso256_2.tranche2.t3[0] ;
 wire \siso256_2.tranche2.t3[1] ;
 wire \siso256_2.tranche2.t3[2] ;
 wire \siso256_2.tranche2.t3[3] ;
 wire \siso256_2.tranche2.tranche0.slice0.latch ;
 wire \siso256_2.tranche2.tranche0.slice0.latch_n ;
 wire \siso256_2.tranche2.tranche0.slice0.siso_out[0] ;
 wire \siso256_2.tranche2.tranche0.slice0.siso_out[1] ;
 wire \siso256_2.tranche2.tranche0.slice0.siso_out[2] ;
 wire \siso256_2.tranche2.tranche0.slice0.siso_out[3] ;
 wire \siso256_2.tranche2.tranche0.slice1.latch ;
 wire \siso256_2.tranche2.tranche0.slice1.latch_n ;
 wire \siso256_2.tranche2.tranche0.slice1.siso_out[0] ;
 wire \siso256_2.tranche2.tranche0.slice1.siso_out[1] ;
 wire \siso256_2.tranche2.tranche0.slice1.siso_out[2] ;
 wire \siso256_2.tranche2.tranche0.slice1.siso_out[3] ;
 wire \siso256_2.tranche2.tranche0.slice2.latch ;
 wire \siso256_2.tranche2.tranche0.slice2.latch_n ;
 wire \siso256_2.tranche2.tranche0.slice2.siso_out[0] ;
 wire \siso256_2.tranche2.tranche0.slice2.siso_out[1] ;
 wire \siso256_2.tranche2.tranche0.slice2.siso_out[2] ;
 wire \siso256_2.tranche2.tranche0.slice2.siso_out[3] ;
 wire \siso256_2.tranche2.tranche0.slice3.latch ;
 wire \siso256_2.tranche2.tranche0.slice3.latch_n ;
 wire \siso256_2.tranche2.tranche1.slice0.latch_n ;
 wire \siso256_2.tranche2.tranche1.slice0.siso_out[0] ;
 wire \siso256_2.tranche2.tranche1.slice0.siso_out[1] ;
 wire \siso256_2.tranche2.tranche1.slice0.siso_out[2] ;
 wire \siso256_2.tranche2.tranche1.slice0.siso_out[3] ;
 wire \siso256_2.tranche2.tranche1.slice1.latch_n ;
 wire \siso256_2.tranche2.tranche1.slice1.siso_out[0] ;
 wire \siso256_2.tranche2.tranche1.slice1.siso_out[1] ;
 wire \siso256_2.tranche2.tranche1.slice1.siso_out[2] ;
 wire \siso256_2.tranche2.tranche1.slice1.siso_out[3] ;
 wire \siso256_2.tranche2.tranche1.slice2.latch_n ;
 wire \siso256_2.tranche2.tranche1.slice2.siso_out[0] ;
 wire \siso256_2.tranche2.tranche1.slice2.siso_out[1] ;
 wire \siso256_2.tranche2.tranche1.slice2.siso_out[2] ;
 wire \siso256_2.tranche2.tranche1.slice2.siso_out[3] ;
 wire \siso256_2.tranche2.tranche1.slice3.latch_n ;
 wire \siso256_2.tranche2.tranche2.slice0.latch_n ;
 wire \siso256_2.tranche2.tranche2.slice0.siso_out[0] ;
 wire \siso256_2.tranche2.tranche2.slice0.siso_out[1] ;
 wire \siso256_2.tranche2.tranche2.slice0.siso_out[2] ;
 wire \siso256_2.tranche2.tranche2.slice0.siso_out[3] ;
 wire \siso256_2.tranche2.tranche2.slice1.latch_n ;
 wire \siso256_2.tranche2.tranche2.slice1.siso_out[0] ;
 wire \siso256_2.tranche2.tranche2.slice1.siso_out[1] ;
 wire \siso256_2.tranche2.tranche2.slice1.siso_out[2] ;
 wire \siso256_2.tranche2.tranche2.slice1.siso_out[3] ;
 wire \siso256_2.tranche2.tranche2.slice2.latch_n ;
 wire \siso256_2.tranche2.tranche2.slice2.siso_out[0] ;
 wire \siso256_2.tranche2.tranche2.slice2.siso_out[1] ;
 wire \siso256_2.tranche2.tranche2.slice2.siso_out[2] ;
 wire \siso256_2.tranche2.tranche2.slice2.siso_out[3] ;
 wire \siso256_2.tranche2.tranche2.slice3.latch_n ;
 wire \siso256_2.tranche2.tranche3.slice0.latch_n ;
 wire \siso256_2.tranche2.tranche3.slice0.siso_out[0] ;
 wire \siso256_2.tranche2.tranche3.slice0.siso_out[1] ;
 wire \siso256_2.tranche2.tranche3.slice0.siso_out[2] ;
 wire \siso256_2.tranche2.tranche3.slice0.siso_out[3] ;
 wire \siso256_2.tranche2.tranche3.slice1.latch_n ;
 wire \siso256_2.tranche2.tranche3.slice1.siso_out[0] ;
 wire \siso256_2.tranche2.tranche3.slice1.siso_out[1] ;
 wire \siso256_2.tranche2.tranche3.slice1.siso_out[2] ;
 wire \siso256_2.tranche2.tranche3.slice1.siso_out[3] ;
 wire \siso256_2.tranche2.tranche3.slice2.latch_n ;
 wire \siso256_2.tranche2.tranche3.slice2.siso_out[0] ;
 wire \siso256_2.tranche2.tranche3.slice2.siso_out[1] ;
 wire \siso256_2.tranche2.tranche3.slice2.siso_out[2] ;
 wire \siso256_2.tranche2.tranche3.slice2.siso_out[3] ;
 wire \siso256_2.tranche2.tranche3.slice3.latch_n ;
 wire \siso256_2.tranche3.t1[0] ;
 wire \siso256_2.tranche3.t1[1] ;
 wire \siso256_2.tranche3.t1[2] ;
 wire \siso256_2.tranche3.t1[3] ;
 wire \siso256_2.tranche3.t2[0] ;
 wire \siso256_2.tranche3.t2[1] ;
 wire \siso256_2.tranche3.t2[2] ;
 wire \siso256_2.tranche3.t2[3] ;
 wire \siso256_2.tranche3.t3[0] ;
 wire \siso256_2.tranche3.t3[1] ;
 wire \siso256_2.tranche3.t3[2] ;
 wire \siso256_2.tranche3.t3[3] ;
 wire \siso256_2.tranche3.tranche0.slice0.latch ;
 wire \siso256_2.tranche3.tranche0.slice0.latch_n ;
 wire \siso256_2.tranche3.tranche0.slice0.siso_out[0] ;
 wire \siso256_2.tranche3.tranche0.slice0.siso_out[1] ;
 wire \siso256_2.tranche3.tranche0.slice0.siso_out[2] ;
 wire \siso256_2.tranche3.tranche0.slice0.siso_out[3] ;
 wire \siso256_2.tranche3.tranche0.slice1.latch ;
 wire \siso256_2.tranche3.tranche0.slice1.latch_n ;
 wire \siso256_2.tranche3.tranche0.slice1.siso_out[0] ;
 wire \siso256_2.tranche3.tranche0.slice1.siso_out[1] ;
 wire \siso256_2.tranche3.tranche0.slice1.siso_out[2] ;
 wire \siso256_2.tranche3.tranche0.slice1.siso_out[3] ;
 wire \siso256_2.tranche3.tranche0.slice2.latch ;
 wire \siso256_2.tranche3.tranche0.slice2.latch_n ;
 wire \siso256_2.tranche3.tranche0.slice2.siso_out[0] ;
 wire \siso256_2.tranche3.tranche0.slice2.siso_out[1] ;
 wire \siso256_2.tranche3.tranche0.slice2.siso_out[2] ;
 wire \siso256_2.tranche3.tranche0.slice2.siso_out[3] ;
 wire \siso256_2.tranche3.tranche0.slice3.latch ;
 wire \siso256_2.tranche3.tranche0.slice3.latch_n ;
 wire \siso256_2.tranche3.tranche1.slice0.latch_n ;
 wire \siso256_2.tranche3.tranche1.slice0.siso_out[0] ;
 wire \siso256_2.tranche3.tranche1.slice0.siso_out[1] ;
 wire \siso256_2.tranche3.tranche1.slice0.siso_out[2] ;
 wire \siso256_2.tranche3.tranche1.slice0.siso_out[3] ;
 wire \siso256_2.tranche3.tranche1.slice1.latch_n ;
 wire \siso256_2.tranche3.tranche1.slice1.siso_out[0] ;
 wire \siso256_2.tranche3.tranche1.slice1.siso_out[1] ;
 wire \siso256_2.tranche3.tranche1.slice1.siso_out[2] ;
 wire \siso256_2.tranche3.tranche1.slice1.siso_out[3] ;
 wire \siso256_2.tranche3.tranche1.slice2.latch_n ;
 wire \siso256_2.tranche3.tranche1.slice2.siso_out[0] ;
 wire \siso256_2.tranche3.tranche1.slice2.siso_out[1] ;
 wire \siso256_2.tranche3.tranche1.slice2.siso_out[2] ;
 wire \siso256_2.tranche3.tranche1.slice2.siso_out[3] ;
 wire \siso256_2.tranche3.tranche1.slice3.latch_n ;
 wire \siso256_2.tranche3.tranche2.slice0.latch_n ;
 wire \siso256_2.tranche3.tranche2.slice0.siso_out[0] ;
 wire \siso256_2.tranche3.tranche2.slice0.siso_out[1] ;
 wire \siso256_2.tranche3.tranche2.slice0.siso_out[2] ;
 wire \siso256_2.tranche3.tranche2.slice0.siso_out[3] ;
 wire \siso256_2.tranche3.tranche2.slice1.latch_n ;
 wire \siso256_2.tranche3.tranche2.slice1.siso_out[0] ;
 wire \siso256_2.tranche3.tranche2.slice1.siso_out[1] ;
 wire \siso256_2.tranche3.tranche2.slice1.siso_out[2] ;
 wire \siso256_2.tranche3.tranche2.slice1.siso_out[3] ;
 wire \siso256_2.tranche3.tranche2.slice2.latch_n ;
 wire \siso256_2.tranche3.tranche2.slice2.siso_out[0] ;
 wire \siso256_2.tranche3.tranche2.slice2.siso_out[1] ;
 wire \siso256_2.tranche3.tranche2.slice2.siso_out[2] ;
 wire \siso256_2.tranche3.tranche2.slice2.siso_out[3] ;
 wire \siso256_2.tranche3.tranche2.slice3.latch_n ;
 wire \siso256_2.tranche3.tranche3.slice0.latch_n ;
 wire \siso256_2.tranche3.tranche3.slice0.siso_out[0] ;
 wire \siso256_2.tranche3.tranche3.slice0.siso_out[1] ;
 wire \siso256_2.tranche3.tranche3.slice0.siso_out[2] ;
 wire \siso256_2.tranche3.tranche3.slice0.siso_out[3] ;
 wire \siso256_2.tranche3.tranche3.slice1.latch_n ;
 wire \siso256_2.tranche3.tranche3.slice1.siso_out[0] ;
 wire \siso256_2.tranche3.tranche3.slice1.siso_out[1] ;
 wire \siso256_2.tranche3.tranche3.slice1.siso_out[2] ;
 wire \siso256_2.tranche3.tranche3.slice1.siso_out[3] ;
 wire \siso256_2.tranche3.tranche3.slice2.latch_n ;
 wire \siso256_2.tranche3.tranche3.slice2.siso_out[0] ;
 wire \siso256_2.tranche3.tranche3.slice2.siso_out[1] ;
 wire \siso256_2.tranche3.tranche3.slice2.siso_out[2] ;
 wire \siso256_2.tranche3.tranche3.slice2.siso_out[3] ;
 wire \siso256_2.tranche3.tranche3.slice3.latch_n ;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire CLK_OUT_regs;
 wire net3;
 wire net4;
 wire net1;
 wire net2;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_0_CLK_OUT;
 wire clknet_1_0__leaf_CLK_OUT;
 wire clknet_0_CLK_OUT_regs;
 wire clknet_2_0__leaf_CLK_OUT_regs;
 wire clknet_2_1__leaf_CLK_OUT_regs;
 wire clknet_2_2__leaf_CLK_OUT_regs;
 wire clknet_2_3__leaf_CLK_OUT_regs;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;

 sg13g2_dfrbpq_1 DFF_reset (.RESET_B(net1),
    .D(net6),
    .Q(INT_RESET),
    .CLK(clknet_2_1__leaf_CLK_OUT_regs));
 sg13g2_dfrbp_1 \J8.DFF_J1  (.RESET_B(\J8.rst1 ),
    .D(net24),
    .Q(uo_out[2]),
    .Q_N(\J8.J4N[0] ),
    .CLK(clknet_2_0__leaf_CLK_OUT_regs));
 sg13g2_dfrbp_1 \J8.DFF_J2  (.RESET_B(\J8.rst1 ),
    .D(net25),
    .Q(uo_out[3]),
    .Q_N(\J8.J4N[1] ),
    .CLK(clknet_2_0__leaf_CLK_OUT_regs));
 sg13g2_dfrbp_1 \J8.DFF_J3  (.RESET_B(\J8.rst1 ),
    .D(net27),
    .Q(uo_out[4]),
    .Q_N(\J8.J4N[2] ),
    .CLK(clknet_2_0__leaf_CLK_OUT_regs));
 sg13g2_dfrbp_1 \J8.DFF_J4  (.RESET_B(\J8.rst1 ),
    .D(net26),
    .Q(uo_out[5]),
    .Q_N(\J8.J4N[3] ),
    .CLK(clknet_2_0__leaf_CLK_OUT_regs));
 sg13g2_inv_2 \J8.boost0  (.Y(\J8.rst ),
    .A(net4));
 sg13g2_inv_2 \J8.boost1  (.Y(\J8.rst1 ),
    .A(\J8.rst ));
 sg13g2_inv_2 \J8.boost2  (.Y(\J8.rst2 ),
    .A(\J8.rst ));
 sg13g2_inv_2 \J8.boost3  (.Y(\J8.rst3 ),
    .A(\J8.rst ));
 sg13g2_inv_2 \J8.boosta  (.Y(\Decoded8[0] ),
    .A(\J8.DecN[0] ));
 sg13g2_inv_1 \J8.boostb  (.Y(\Decoded8[1] ),
    .A(\J8.DecN[1] ));
 sg13g2_inv_2 \J8.boostc  (.Y(\Decoded8[2] ),
    .A(\J8.DecN[2] ));
 sg13g2_inv_1 \J8.boostd  (.Y(\Decoded8[3] ),
    .A(\J8.DecN[3] ));
 sg13g2_inv_2 \J8.booste  (.Y(\Decoded8[4] ),
    .A(\J8.DecN[4] ));
 sg13g2_inv_1 \J8.boostf  (.Y(\Decoded8[5] ),
    .A(\J8.DecN[5] ));
 sg13g2_inv_2 \J8.boostg  (.Y(\Decoded8[6] ),
    .A(\J8.DecN[6] ));
 sg13g2_inv_1 \J8.boosth  (.Y(\Decoded8[7] ),
    .A(\J8.DecN[7] ));
 sg13g2_nand3_1 \J8.dec0  (.B(\J8.J4N[0] ),
    .C(\J8.rst2 ),
    .A(\J8.J4N[3] ),
    .Y(\J8.DecN[0] ));
 sg13g2_nand3_1 \J8.dec1  (.B(\J8.J4N[1] ),
    .C(\J8.rst2 ),
    .A(uo_out[2]),
    .Y(\J8.DecN[1] ));
 sg13g2_nand3_1 \J8.dec2  (.B(\J8.J4N[2] ),
    .C(\J8.rst2 ),
    .A(uo_out[3]),
    .Y(\J8.DecN[2] ));
 sg13g2_nand3_1 \J8.dec3  (.B(\J8.J4N[3] ),
    .C(\J8.rst2 ),
    .A(uo_out[4]),
    .Y(\J8.DecN[3] ));
 sg13g2_nand3_1 \J8.dec4  (.B(uo_out[2]),
    .C(\J8.rst3 ),
    .A(uo_out[5]),
    .Y(\J8.DecN[4] ));
 sg13g2_nand3_1 \J8.dec5  (.B(net27),
    .C(\J8.rst3 ),
    .A(net38),
    .Y(\J8.DecN[5] ));
 sg13g2_nand3_1 \J8.dec6  (.B(uo_out[4]),
    .C(\J8.rst3 ),
    .A(\J8.J4N[1] ),
    .Y(\J8.DecN[6] ));
 sg13g2_nand3_1 \J8.dec7  (.B(uo_out[5]),
    .C(\J8.rst3 ),
    .A(\J8.J4N[2] ),
    .Y(\J8.DecN[7] ));
 sg13g2_mux2_1 _00_ (.A0(\Decoded8[0] ),
    .A1(LFSR_BIT),
    .S(net9),
    .X(uio_out[0]));
 sg13g2_mux2_1 _01_ (.A0(\Decoded8[1] ),
    .A1(\LFSR_state8[1] ),
    .S(net9),
    .X(uio_out[1]));
 sg13g2_mux2_1 _02_ (.A0(\Decoded8[2] ),
    .A1(\LFSR_state8[2] ),
    .S(net9),
    .X(uio_out[2]));
 sg13g2_mux2_1 _03_ (.A0(\Decoded8[3] ),
    .A1(\LFSR_state8[3] ),
    .S(net9),
    .X(uio_out[3]));
 sg13g2_mux2_1 _04_ (.A0(\Decoded8[4] ),
    .A1(\LFSR_state8[4] ),
    .S(net9),
    .X(uio_out[4]));
 sg13g2_mux2_1 _05_ (.A0(\Decoded8[5] ),
    .A1(\LFSR_state8[5] ),
    .S(net9),
    .X(uio_out[5]));
 sg13g2_mux2_1 _06_ (.A0(\Decoded8[6] ),
    .A1(\LFSR_state8[6] ),
    .S(net9),
    .X(uio_out[6]));
 sg13g2_mux2_1 _07_ (.A0(\Decoded8[7] ),
    .A1(\LFSR_state8[7] ),
    .S(net9),
    .X(uio_out[7]));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_11 (.L_HI(net13));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_12 (.L_HI(net14));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_13 (.L_HI(net15));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_14 (.L_HI(net16));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_15 (.L_HI(net17));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_16 (.L_HI(net18));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_17 (.L_HI(net19));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(CLK_OUT),
    .X(CLK_OUT_regs));
 sg13g2_buf_1 _16_ (.A(clknet_1_0__leaf_CLK_OUT),
    .X(uo_out[1]));
 sg13g2_buf_1 _17_ (.A(LFSR_PERIOD),
    .X(uo_out[6]));
 sg13g2_buf_1 _18_ (.A(LFSR_BIT),
    .X(uo_out[7]));
 sg13g2_dfrbpq_2 \lfsr.lfsr0  (.RESET_B(net3),
    .D(net33),
    .Q(LFSR_BIT),
    .CLK(clknet_2_3__leaf_CLK_OUT_regs));
 sg13g2_dfrbp_1 \lfsr.lfsr1  (.RESET_B(net3),
    .D(net23),
    .Q(\lfsr.dum2 ),
    .Q_N(\LFSR_state8[1] ),
    .CLK(clknet_2_2__leaf_CLK_OUT_regs));
 sg13g2_dfrbp_1 \lfsr.lfsr2  (.RESET_B(net3),
    .D(net29),
    .Q(\lfsr.dum1 ),
    .Q_N(\LFSR_state8[2] ),
    .CLK(clknet_2_3__leaf_CLK_OUT_regs));
 sg13g2_dfrbpq_1 \lfsr.lfsr3  (.RESET_B(net3),
    .D(net20),
    .Q(\LFSR_state8[3] ),
    .CLK(clknet_2_2__leaf_CLK_OUT_regs));
 sg13g2_dfrbpq_1 \lfsr.lfsr4  (.RESET_B(net3),
    .D(net31),
    .Q(\LFSR_state8[4] ),
    .CLK(clknet_2_1__leaf_CLK_OUT_regs));
 sg13g2_dfrbpq_1 \lfsr.lfsr5  (.RESET_B(net3),
    .D(net21),
    .Q(\LFSR_state8[5] ),
    .CLK(clknet_2_2__leaf_CLK_OUT_regs));
 sg13g2_dfrbpq_1 \lfsr.lfsr6  (.RESET_B(net3),
    .D(net22),
    .Q(\LFSR_state8[6] ),
    .CLK(clknet_2_1__leaf_CLK_OUT_regs));
 sg13g2_dfrbpq_1 \lfsr.lfsr7  (.RESET_B(net3),
    .D(\lfsr.feedback ),
    .Q(\LFSR_state8[7] ),
    .CLK(clknet_2_1__leaf_CLK_OUT_regs));
 sg13g2_and4_1 \lfsr.period4_1  (.A(LFSR_BIT),
    .B(\LFSR_state8[1] ),
    .C(\LFSR_state8[2] ),
    .D(\LFSR_state8[3] ),
    .X(\lfsr.and8_1 ));
 sg13g2_and4_1 \lfsr.period4_2  (.A(\LFSR_state8[4] ),
    .B(\LFSR_state8[5] ),
    .C(\LFSR_state8[6] ),
    .D(\LFSR_state8[7] ),
    .X(\lfsr.and8_2 ));
 sg13g2_and2_1 \lfsr.period8  (.A(\lfsr.and8_1 ),
    .B(\lfsr.and8_2 ),
    .X(LFSR_PERIOD));
 sg13g2_and2_1 \lfsr.stall  (.A(net35),
    .B(net10),
    .X(\lfsr.feedback ));
 sg13g2_xor2_1 \lfsr.x_a  (.B(net30),
    .A(\lfsr.feedback ),
    .X(\lfsr.x1 ));
 sg13g2_xor2_1 \lfsr.x_b  (.B(net28),
    .A(\lfsr.feedback ),
    .X(\lfsr.x2 ));
 sg13g2_xor2_1 \lfsr.x_c  (.B(net32),
    .A(\lfsr.feedback ),
    .X(\lfsr.x3 ));
 sg13g2_mux2_1 mux2_Din (.A0(DL_out),
    .A1(MX_out),
    .S(net8),
    .X(uo_out[0]));
 sg13g2_mux2_2 mux_clk (.A0(clk),
    .A1(net5),
    .S(net2),
    .X(CLK_OUT));
 sg13g2_inv_2 \siso256_1.Amp0.Amp0  (.Y(\siso256_1.Amp0.Y[0] ),
    .A(\Decoded8[6] ));
 sg13g2_inv_2 \siso256_1.Amp0.Amp1  (.Y(\siso256_1.Amp0.Y[1] ),
    .A(\Decoded8[4] ));
 sg13g2_inv_2 \siso256_1.Amp0.Amp2  (.Y(\siso256_1.Amp0.Y[2] ),
    .A(\Decoded8[2] ));
 sg13g2_inv_2 \siso256_1.Amp0.Amp3  (.Y(\siso256_1.Amp0.Y[3] ),
    .A(\Decoded8[0] ));
 sg13g2_inv_1 \siso256_1.Amp1.Amp0  (.Y(\siso256_1.Amp1.Y[0] ),
    .A(\siso256_1.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_1.Amp1.Amp1  (.Y(\siso256_1.Amp1.Y[1] ),
    .A(\siso256_1.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_1.Amp1.Amp2  (.Y(\siso256_1.Amp1.Y[2] ),
    .A(\siso256_1.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_1.Amp1.Amp3  (.Y(\siso256_1.Amp1.Y[3] ),
    .A(\siso256_1.Amp0.Y[3] ));
 sg13g2_inv_1 \siso256_1.Amp2.Amp0  (.Y(\siso256_1.Amp2.Y[0] ),
    .A(\siso256_1.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_1.Amp2.Amp1  (.Y(\siso256_1.Amp2.Y[1] ),
    .A(\siso256_1.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_1.Amp2.Amp2  (.Y(\siso256_1.Amp2.Y[2] ),
    .A(\siso256_1.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_1.Amp2.Amp3  (.Y(\siso256_1.Amp2.Y[3] ),
    .A(\siso256_1.Amp0.Y[3] ));
 sg13g2_inv_1 \siso256_1.Amp3.Amp0  (.Y(\siso256_1.Amp3.Y[0] ),
    .A(\siso256_1.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_1.Amp3.Amp1  (.Y(\siso256_1.Amp3.Y[1] ),
    .A(\siso256_1.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_1.Amp3.Amp2  (.Y(\siso256_1.Amp3.Y[2] ),
    .A(\siso256_1.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_1.Amp3.Amp3  (.Y(\siso256_1.Amp3.Y[3] ),
    .A(\siso256_1.Amp0.Y[3] ));
 sg13g2_inv_1 \siso256_1.Amp4.Amp0  (.Y(\siso256_1.Amp4.Y[0] ),
    .A(\siso256_1.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_1.Amp4.Amp1  (.Y(\siso256_1.Amp4.Y[1] ),
    .A(\siso256_1.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_1.Amp4.Amp2  (.Y(\siso256_1.Amp4.Y[2] ),
    .A(\siso256_1.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_1.Amp4.Amp3  (.Y(\siso256_1.Amp4.Y[3] ),
    .A(\siso256_1.Amp0.Y[3] ));
 sg13g2_inv_2 \siso256_1.tranche0.Amp.Amp0  (.Y(\siso256_1.tranche0.tranche0.slice3.latch ),
    .A(\siso256_1.Amp1.Y[0] ));
 sg13g2_inv_2 \siso256_1.tranche0.Amp.Amp1  (.Y(\siso256_1.tranche0.tranche0.slice2.latch ),
    .A(\siso256_1.Amp1.Y[1] ));
 sg13g2_inv_2 \siso256_1.tranche0.Amp.Amp2  (.Y(\siso256_1.tranche0.tranche0.slice1.latch ),
    .A(\siso256_1.Amp1.Y[2] ));
 sg13g2_inv_2 \siso256_1.tranche0.Amp.Amp3  (.Y(\siso256_1.tranche0.tranche0.slice0.latch ),
    .A(\siso256_1.Amp1.Y[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche0.slice0.Amp  (.Y(\siso256_1.tranche0.tranche0.slice0.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice0.l0  (.D(back),
    .GATE(\siso256_1.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice0.l1  (.D(\siso256_1.siso_in[1] ),
    .GATE(\siso256_1.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice0.l2  (.D(MX_out),
    .GATE(\siso256_1.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice0.l3  (.D(\siso256_1.siso_in[3] ),
    .GATE(\siso256_1.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche0.slice1.Amp  (.Y(\siso256_1.tranche0.tranche0.slice1.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice1.l0  (.D(\siso256_1.tranche0.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice1.l1  (.D(\siso256_1.tranche0.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice1.l2  (.D(\siso256_1.tranche0.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice1.l3  (.D(\siso256_1.tranche0.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche0.slice2.Amp  (.Y(\siso256_1.tranche0.tranche0.slice2.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice2.l0  (.D(\siso256_1.tranche0.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice2.l1  (.D(\siso256_1.tranche0.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice2.l2  (.D(\siso256_1.tranche0.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice2.l3  (.D(\siso256_1.tranche0.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche0.slice3.Amp  (.Y(\siso256_1.tranche0.tranche0.slice3.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice3.l0  (.D(\siso256_1.tranche0.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t1[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice3.l1  (.D(\siso256_1.tranche0.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t1[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice3.l2  (.D(\siso256_1.tranche0.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t1[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche0.slice3.l3  (.D(\siso256_1.tranche0.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t1[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche1.slice0.Amp  (.Y(\siso256_1.tranche0.tranche1.slice0.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice0.l0  (.D(\siso256_1.tranche0.t1[0] ),
    .GATE(\siso256_1.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice0.l1  (.D(\siso256_1.tranche0.t1[1] ),
    .GATE(\siso256_1.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice0.l2  (.D(\siso256_1.tranche0.t1[2] ),
    .GATE(\siso256_1.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice0.l3  (.D(\siso256_1.tranche0.t1[3] ),
    .GATE(\siso256_1.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche1.slice1.Amp  (.Y(\siso256_1.tranche0.tranche1.slice1.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice1.l0  (.D(\siso256_1.tranche0.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice1.l1  (.D(\siso256_1.tranche0.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice1.l2  (.D(\siso256_1.tranche0.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice1.l3  (.D(\siso256_1.tranche0.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_2 \siso256_1.tranche0.tranche1.slice2.Amp  (.Y(\siso256_1.tranche0.tranche1.slice2.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice2.l0  (.D(\siso256_1.tranche0.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice2.l1  (.D(\siso256_1.tranche0.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice2.l2  (.D(\siso256_1.tranche0.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice2.l3  (.D(\siso256_1.tranche0.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche1.slice3.Amp  (.Y(\siso256_1.tranche0.tranche1.slice3.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice3.l0  (.D(\siso256_1.tranche0.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t2[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice3.l1  (.D(\siso256_1.tranche0.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t2[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice3.l2  (.D(\siso256_1.tranche0.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t2[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche1.slice3.l3  (.D(\siso256_1.tranche0.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t2[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche2.slice0.Amp  (.Y(\siso256_1.tranche0.tranche2.slice0.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice0.l0  (.D(\siso256_1.tranche0.t2[0] ),
    .GATE(\siso256_1.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice0.l1  (.D(\siso256_1.tranche0.t2[1] ),
    .GATE(\siso256_1.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice0.l2  (.D(\siso256_1.tranche0.t2[2] ),
    .GATE(\siso256_1.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice0.l3  (.D(\siso256_1.tranche0.t2[3] ),
    .GATE(\siso256_1.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche2.slice1.Amp  (.Y(\siso256_1.tranche0.tranche2.slice1.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice1.l0  (.D(\siso256_1.tranche0.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice1.l1  (.D(\siso256_1.tranche0.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice1.l2  (.D(\siso256_1.tranche0.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice1.l3  (.D(\siso256_1.tranche0.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche2.slice2.Amp  (.Y(\siso256_1.tranche0.tranche2.slice2.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice2.l0  (.D(\siso256_1.tranche0.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice2.l1  (.D(\siso256_1.tranche0.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice2.l2  (.D(\siso256_1.tranche0.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice2.l3  (.D(\siso256_1.tranche0.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche2.slice3.Amp  (.Y(\siso256_1.tranche0.tranche2.slice3.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice3.l0  (.D(\siso256_1.tranche0.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t3[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice3.l1  (.D(\siso256_1.tranche0.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t3[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice3.l2  (.D(\siso256_1.tranche0.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t3[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche2.slice3.l3  (.D(\siso256_1.tranche0.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche0.t3[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche3.slice0.Amp  (.Y(\siso256_1.tranche0.tranche3.slice0.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice0.l0  (.D(\siso256_1.tranche0.t3[0] ),
    .GATE(\siso256_1.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice0.l1  (.D(\siso256_1.tranche0.t3[1] ),
    .GATE(\siso256_1.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice0.l2  (.D(\siso256_1.tranche0.t3[2] ),
    .GATE(\siso256_1.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice0.l3  (.D(\siso256_1.tranche0.t3[3] ),
    .GATE(\siso256_1.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche3.slice1.Amp  (.Y(\siso256_1.tranche0.tranche3.slice1.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice1.l0  (.D(\siso256_1.tranche0.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice1.l1  (.D(\siso256_1.tranche0.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice1.l2  (.D(\siso256_1.tranche0.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice1.l3  (.D(\siso256_1.tranche0.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche3.slice2.Amp  (.Y(\siso256_1.tranche0.tranche3.slice2.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice2.l0  (.D(\siso256_1.tranche0.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice2.l1  (.D(\siso256_1.tranche0.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice2.l2  (.D(\siso256_1.tranche0.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice2.l3  (.D(\siso256_1.tranche0.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche0.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche0.tranche3.slice3.Amp  (.Y(\siso256_1.tranche0.tranche3.slice3.latch_n ),
    .A(\siso256_1.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice3.l0  (.D(\siso256_1.tranche0.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t1[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice3.l1  (.D(\siso256_1.tranche0.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t1[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice3.l2  (.D(\siso256_1.tranche0.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t1[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche0.tranche3.slice3.l3  (.D(\siso256_1.tranche0.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t1[3] ));
 sg13g2_inv_2 \siso256_1.tranche1.Amp.Amp0  (.Y(\siso256_1.tranche1.tranche0.slice3.latch ),
    .A(\siso256_1.Amp2.Y[0] ));
 sg13g2_inv_2 \siso256_1.tranche1.Amp.Amp1  (.Y(\siso256_1.tranche1.tranche0.slice2.latch ),
    .A(\siso256_1.Amp2.Y[1] ));
 sg13g2_inv_2 \siso256_1.tranche1.Amp.Amp2  (.Y(\siso256_1.tranche1.tranche0.slice1.latch ),
    .A(\siso256_1.Amp2.Y[2] ));
 sg13g2_inv_2 \siso256_1.tranche1.Amp.Amp3  (.Y(\siso256_1.tranche1.tranche0.slice0.latch ),
    .A(\siso256_1.Amp2.Y[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche0.slice0.Amp  (.Y(\siso256_1.tranche1.tranche0.slice0.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice0.l0  (.D(\siso256_1.t1[0] ),
    .GATE(\siso256_1.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice0.l1  (.D(\siso256_1.t1[1] ),
    .GATE(\siso256_1.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice0.l2  (.D(\siso256_1.t1[2] ),
    .GATE(\siso256_1.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice0.l3  (.D(\siso256_1.t1[3] ),
    .GATE(\siso256_1.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche0.slice1.Amp  (.Y(\siso256_1.tranche1.tranche0.slice1.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice1.l0  (.D(\siso256_1.tranche1.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice1.l1  (.D(\siso256_1.tranche1.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice1.l2  (.D(\siso256_1.tranche1.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice1.l3  (.D(\siso256_1.tranche1.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche0.slice2.Amp  (.Y(\siso256_1.tranche1.tranche0.slice2.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice2.l0  (.D(\siso256_1.tranche1.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice2.l1  (.D(\siso256_1.tranche1.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice2.l2  (.D(\siso256_1.tranche1.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice2.l3  (.D(\siso256_1.tranche1.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche0.slice3.Amp  (.Y(\siso256_1.tranche1.tranche0.slice3.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice3.l0  (.D(\siso256_1.tranche1.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t1[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice3.l1  (.D(\siso256_1.tranche1.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t1[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice3.l2  (.D(\siso256_1.tranche1.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t1[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche0.slice3.l3  (.D(\siso256_1.tranche1.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t1[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche1.slice0.Amp  (.Y(\siso256_1.tranche1.tranche1.slice0.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice0.l0  (.D(\siso256_1.tranche1.t1[0] ),
    .GATE(\siso256_1.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice0.l1  (.D(\siso256_1.tranche1.t1[1] ),
    .GATE(\siso256_1.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice0.l2  (.D(\siso256_1.tranche1.t1[2] ),
    .GATE(\siso256_1.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice0.l3  (.D(\siso256_1.tranche1.t1[3] ),
    .GATE(\siso256_1.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche1.slice1.Amp  (.Y(\siso256_1.tranche1.tranche1.slice1.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice1.l0  (.D(\siso256_1.tranche1.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice1.l1  (.D(\siso256_1.tranche1.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice1.l2  (.D(\siso256_1.tranche1.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice1.l3  (.D(\siso256_1.tranche1.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche1.slice2.Amp  (.Y(\siso256_1.tranche1.tranche1.slice2.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice2.l0  (.D(\siso256_1.tranche1.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice2.l1  (.D(\siso256_1.tranche1.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice2.l2  (.D(\siso256_1.tranche1.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice2.l3  (.D(\siso256_1.tranche1.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche1.slice3.Amp  (.Y(\siso256_1.tranche1.tranche1.slice3.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice3.l0  (.D(\siso256_1.tranche1.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t2[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice3.l1  (.D(\siso256_1.tranche1.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t2[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice3.l2  (.D(\siso256_1.tranche1.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t2[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche1.slice3.l3  (.D(\siso256_1.tranche1.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t2[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche2.slice0.Amp  (.Y(\siso256_1.tranche1.tranche2.slice0.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice0.l0  (.D(\siso256_1.tranche1.t2[0] ),
    .GATE(\siso256_1.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice0.l1  (.D(\siso256_1.tranche1.t2[1] ),
    .GATE(\siso256_1.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice0.l2  (.D(\siso256_1.tranche1.t2[2] ),
    .GATE(\siso256_1.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice0.l3  (.D(\siso256_1.tranche1.t2[3] ),
    .GATE(\siso256_1.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche2.slice1.Amp  (.Y(\siso256_1.tranche1.tranche2.slice1.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice1.l0  (.D(\siso256_1.tranche1.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice1.l1  (.D(\siso256_1.tranche1.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice1.l2  (.D(\siso256_1.tranche1.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice1.l3  (.D(\siso256_1.tranche1.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche2.slice2.Amp  (.Y(\siso256_1.tranche1.tranche2.slice2.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice2.l0  (.D(\siso256_1.tranche1.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice2.l1  (.D(\siso256_1.tranche1.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice2.l2  (.D(\siso256_1.tranche1.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice2.l3  (.D(\siso256_1.tranche1.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche2.slice3.Amp  (.Y(\siso256_1.tranche1.tranche2.slice3.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice3.l0  (.D(\siso256_1.tranche1.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t3[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice3.l1  (.D(\siso256_1.tranche1.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t3[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice3.l2  (.D(\siso256_1.tranche1.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t3[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche2.slice3.l3  (.D(\siso256_1.tranche1.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche1.t3[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche3.slice0.Amp  (.Y(\siso256_1.tranche1.tranche3.slice0.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice0.l0  (.D(\siso256_1.tranche1.t3[0] ),
    .GATE(\siso256_1.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice0.l1  (.D(\siso256_1.tranche1.t3[1] ),
    .GATE(\siso256_1.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice0.l2  (.D(\siso256_1.tranche1.t3[2] ),
    .GATE(\siso256_1.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice0.l3  (.D(\siso256_1.tranche1.t3[3] ),
    .GATE(\siso256_1.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche3.slice1.Amp  (.Y(\siso256_1.tranche1.tranche3.slice1.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice1.l0  (.D(\siso256_1.tranche1.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice1.l1  (.D(\siso256_1.tranche1.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice1.l2  (.D(\siso256_1.tranche1.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice1.l3  (.D(\siso256_1.tranche1.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche3.slice2.Amp  (.Y(\siso256_1.tranche1.tranche3.slice2.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice2.l0  (.D(\siso256_1.tranche1.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice2.l1  (.D(\siso256_1.tranche1.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice2.l2  (.D(\siso256_1.tranche1.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice2.l3  (.D(\siso256_1.tranche1.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche1.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche1.tranche3.slice3.Amp  (.Y(\siso256_1.tranche1.tranche3.slice3.latch_n ),
    .A(\siso256_1.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice3.l0  (.D(\siso256_1.tranche1.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t2[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice3.l1  (.D(\siso256_1.tranche1.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t2[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice3.l2  (.D(\siso256_1.tranche1.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t2[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche1.tranche3.slice3.l3  (.D(\siso256_1.tranche1.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t2[3] ));
 sg13g2_inv_2 \siso256_1.tranche2.Amp.Amp0  (.Y(\siso256_1.tranche2.tranche0.slice3.latch ),
    .A(\siso256_1.Amp3.Y[0] ));
 sg13g2_inv_2 \siso256_1.tranche2.Amp.Amp1  (.Y(\siso256_1.tranche2.tranche0.slice2.latch ),
    .A(\siso256_1.Amp3.Y[1] ));
 sg13g2_inv_2 \siso256_1.tranche2.Amp.Amp2  (.Y(\siso256_1.tranche2.tranche0.slice1.latch ),
    .A(\siso256_1.Amp3.Y[2] ));
 sg13g2_inv_2 \siso256_1.tranche2.Amp.Amp3  (.Y(\siso256_1.tranche2.tranche0.slice0.latch ),
    .A(\siso256_1.Amp3.Y[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche0.slice0.Amp  (.Y(\siso256_1.tranche2.tranche0.slice0.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice0.l0  (.D(\siso256_1.t2[0] ),
    .GATE(\siso256_1.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice0.l1  (.D(\siso256_1.t2[1] ),
    .GATE(\siso256_1.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice0.l2  (.D(\siso256_1.t2[2] ),
    .GATE(\siso256_1.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice0.l3  (.D(\siso256_1.t2[3] ),
    .GATE(\siso256_1.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche0.slice1.Amp  (.Y(\siso256_1.tranche2.tranche0.slice1.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice1.l0  (.D(\siso256_1.tranche2.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice1.l1  (.D(\siso256_1.tranche2.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice1.l2  (.D(\siso256_1.tranche2.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice1.l3  (.D(\siso256_1.tranche2.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche0.slice2.Amp  (.Y(\siso256_1.tranche2.tranche0.slice2.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice2.l0  (.D(\siso256_1.tranche2.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice2.l1  (.D(\siso256_1.tranche2.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice2.l2  (.D(\siso256_1.tranche2.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice2.l3  (.D(\siso256_1.tranche2.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche0.slice3.Amp  (.Y(\siso256_1.tranche2.tranche0.slice3.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice3.l0  (.D(\siso256_1.tranche2.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t1[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice3.l1  (.D(\siso256_1.tranche2.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t1[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice3.l2  (.D(\siso256_1.tranche2.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t1[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche0.slice3.l3  (.D(\siso256_1.tranche2.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t1[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche1.slice0.Amp  (.Y(\siso256_1.tranche2.tranche1.slice0.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice0.l0  (.D(\siso256_1.tranche2.t1[0] ),
    .GATE(\siso256_1.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice0.l1  (.D(\siso256_1.tranche2.t1[1] ),
    .GATE(\siso256_1.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice0.l2  (.D(\siso256_1.tranche2.t1[2] ),
    .GATE(\siso256_1.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice0.l3  (.D(\siso256_1.tranche2.t1[3] ),
    .GATE(\siso256_1.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche1.slice1.Amp  (.Y(\siso256_1.tranche2.tranche1.slice1.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice1.l0  (.D(\siso256_1.tranche2.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice1.l1  (.D(\siso256_1.tranche2.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice1.l2  (.D(\siso256_1.tranche2.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice1.l3  (.D(\siso256_1.tranche2.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche1.slice2.Amp  (.Y(\siso256_1.tranche2.tranche1.slice2.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice2.l0  (.D(\siso256_1.tranche2.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice2.l1  (.D(\siso256_1.tranche2.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice2.l2  (.D(\siso256_1.tranche2.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice2.l3  (.D(\siso256_1.tranche2.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche1.slice3.Amp  (.Y(\siso256_1.tranche2.tranche1.slice3.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice3.l0  (.D(\siso256_1.tranche2.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t2[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice3.l1  (.D(\siso256_1.tranche2.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t2[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice3.l2  (.D(\siso256_1.tranche2.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t2[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche1.slice3.l3  (.D(\siso256_1.tranche2.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t2[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche2.slice0.Amp  (.Y(\siso256_1.tranche2.tranche2.slice0.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice0.l0  (.D(\siso256_1.tranche2.t2[0] ),
    .GATE(\siso256_1.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice0.l1  (.D(\siso256_1.tranche2.t2[1] ),
    .GATE(\siso256_1.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice0.l2  (.D(\siso256_1.tranche2.t2[2] ),
    .GATE(\siso256_1.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice0.l3  (.D(\siso256_1.tranche2.t2[3] ),
    .GATE(\siso256_1.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche2.slice1.Amp  (.Y(\siso256_1.tranche2.tranche2.slice1.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice1.l0  (.D(\siso256_1.tranche2.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice1.l1  (.D(\siso256_1.tranche2.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice1.l2  (.D(\siso256_1.tranche2.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice1.l3  (.D(\siso256_1.tranche2.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche2.slice2.Amp  (.Y(\siso256_1.tranche2.tranche2.slice2.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice2.l0  (.D(\siso256_1.tranche2.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice2.l1  (.D(\siso256_1.tranche2.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice2.l2  (.D(\siso256_1.tranche2.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice2.l3  (.D(\siso256_1.tranche2.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche2.slice3.Amp  (.Y(\siso256_1.tranche2.tranche2.slice3.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice3.l0  (.D(\siso256_1.tranche2.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t3[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice3.l1  (.D(\siso256_1.tranche2.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t3[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice3.l2  (.D(\siso256_1.tranche2.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t3[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche2.slice3.l3  (.D(\siso256_1.tranche2.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche2.t3[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche3.slice0.Amp  (.Y(\siso256_1.tranche2.tranche3.slice0.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice0.l0  (.D(\siso256_1.tranche2.t3[0] ),
    .GATE(\siso256_1.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice0.l1  (.D(\siso256_1.tranche2.t3[1] ),
    .GATE(\siso256_1.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice0.l2  (.D(\siso256_1.tranche2.t3[2] ),
    .GATE(\siso256_1.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice0.l3  (.D(\siso256_1.tranche2.t3[3] ),
    .GATE(\siso256_1.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche3.slice1.Amp  (.Y(\siso256_1.tranche2.tranche3.slice1.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice1.l0  (.D(\siso256_1.tranche2.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice1.l1  (.D(\siso256_1.tranche2.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice1.l2  (.D(\siso256_1.tranche2.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice1.l3  (.D(\siso256_1.tranche2.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche3.slice2.Amp  (.Y(\siso256_1.tranche2.tranche3.slice2.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice2.l0  (.D(\siso256_1.tranche2.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice2.l1  (.D(\siso256_1.tranche2.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice2.l2  (.D(\siso256_1.tranche2.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice2.l3  (.D(\siso256_1.tranche2.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche2.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche2.tranche3.slice3.Amp  (.Y(\siso256_1.tranche2.tranche3.slice3.latch_n ),
    .A(\siso256_1.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice3.l0  (.D(\siso256_1.tranche2.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t3[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice3.l1  (.D(\siso256_1.tranche2.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t3[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice3.l2  (.D(\siso256_1.tranche2.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t3[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche2.tranche3.slice3.l3  (.D(\siso256_1.tranche2.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_1.t3[3] ));
 sg13g2_inv_2 \siso256_1.tranche3.Amp.Amp0  (.Y(\siso256_1.tranche3.tranche0.slice3.latch ),
    .A(\siso256_1.Amp4.Y[0] ));
 sg13g2_inv_2 \siso256_1.tranche3.Amp.Amp1  (.Y(\siso256_1.tranche3.tranche0.slice2.latch ),
    .A(\siso256_1.Amp4.Y[1] ));
 sg13g2_inv_2 \siso256_1.tranche3.Amp.Amp2  (.Y(\siso256_1.tranche3.tranche0.slice1.latch ),
    .A(\siso256_1.Amp4.Y[2] ));
 sg13g2_inv_2 \siso256_1.tranche3.Amp.Amp3  (.Y(\siso256_1.tranche3.tranche0.slice0.latch ),
    .A(\siso256_1.Amp4.Y[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche0.slice0.Amp  (.Y(\siso256_1.tranche3.tranche0.slice0.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice0.l0  (.D(\siso256_1.t3[0] ),
    .GATE(\siso256_1.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice0.l1  (.D(\siso256_1.t3[1] ),
    .GATE(\siso256_1.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice0.l2  (.D(\siso256_1.t3[2] ),
    .GATE(\siso256_1.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice0.l3  (.D(\siso256_1.t3[3] ),
    .GATE(\siso256_1.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche0.slice1.Amp  (.Y(\siso256_1.tranche3.tranche0.slice1.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice1.l0  (.D(\siso256_1.tranche3.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice1.l1  (.D(\siso256_1.tranche3.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice1.l2  (.D(\siso256_1.tranche3.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice1.l3  (.D(\siso256_1.tranche3.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche0.slice2.Amp  (.Y(\siso256_1.tranche3.tranche0.slice2.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice2.l0  (.D(\siso256_1.tranche3.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice2.l1  (.D(\siso256_1.tranche3.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice2.l2  (.D(\siso256_1.tranche3.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice2.l3  (.D(\siso256_1.tranche3.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche0.slice3.Amp  (.Y(\siso256_1.tranche3.tranche0.slice3.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice3.l0  (.D(\siso256_1.tranche3.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t1[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice3.l1  (.D(\siso256_1.tranche3.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t1[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice3.l2  (.D(\siso256_1.tranche3.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t1[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche0.slice3.l3  (.D(\siso256_1.tranche3.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t1[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche1.slice0.Amp  (.Y(\siso256_1.tranche3.tranche1.slice0.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice0.l0  (.D(\siso256_1.tranche3.t1[0] ),
    .GATE(\siso256_1.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice0.l1  (.D(\siso256_1.tranche3.t1[1] ),
    .GATE(\siso256_1.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice0.l2  (.D(\siso256_1.tranche3.t1[2] ),
    .GATE(\siso256_1.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice0.l3  (.D(\siso256_1.tranche3.t1[3] ),
    .GATE(\siso256_1.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche1.slice1.Amp  (.Y(\siso256_1.tranche3.tranche1.slice1.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice1.l0  (.D(\siso256_1.tranche3.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice1.l1  (.D(\siso256_1.tranche3.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice1.l2  (.D(\siso256_1.tranche3.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice1.l3  (.D(\siso256_1.tranche3.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche1.slice2.Amp  (.Y(\siso256_1.tranche3.tranche1.slice2.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice2.l0  (.D(\siso256_1.tranche3.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice2.l1  (.D(\siso256_1.tranche3.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice2.l2  (.D(\siso256_1.tranche3.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice2.l3  (.D(\siso256_1.tranche3.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche1.slice3.Amp  (.Y(\siso256_1.tranche3.tranche1.slice3.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice3.l0  (.D(\siso256_1.tranche3.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t2[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice3.l1  (.D(\siso256_1.tranche3.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t2[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice3.l2  (.D(\siso256_1.tranche3.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t2[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche1.slice3.l3  (.D(\siso256_1.tranche3.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t2[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche2.slice0.Amp  (.Y(\siso256_1.tranche3.tranche2.slice0.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice0.l0  (.D(\siso256_1.tranche3.t2[0] ),
    .GATE(\siso256_1.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice0.l1  (.D(\siso256_1.tranche3.t2[1] ),
    .GATE(\siso256_1.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice0.l2  (.D(\siso256_1.tranche3.t2[2] ),
    .GATE(\siso256_1.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice0.l3  (.D(\siso256_1.tranche3.t2[3] ),
    .GATE(\siso256_1.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche2.slice1.Amp  (.Y(\siso256_1.tranche3.tranche2.slice1.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice1.l0  (.D(\siso256_1.tranche3.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice1.l1  (.D(\siso256_1.tranche3.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice1.l2  (.D(\siso256_1.tranche3.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice1.l3  (.D(\siso256_1.tranche3.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche2.slice2.Amp  (.Y(\siso256_1.tranche3.tranche2.slice2.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice2.l0  (.D(\siso256_1.tranche3.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice2.l1  (.D(\siso256_1.tranche3.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice2.l2  (.D(\siso256_1.tranche3.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice2.l3  (.D(\siso256_1.tranche3.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche2.slice3.Amp  (.Y(\siso256_1.tranche3.tranche2.slice3.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice3.l0  (.D(\siso256_1.tranche3.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t3[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice3.l1  (.D(\siso256_1.tranche3.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t3[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice3.l2  (.D(\siso256_1.tranche3.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t3[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche2.slice3.l3  (.D(\siso256_1.tranche3.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_1.tranche3.t3[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche3.slice0.Amp  (.Y(\siso256_1.tranche3.tranche3.slice0.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice0.l0  (.D(\siso256_1.tranche3.t3[0] ),
    .GATE(\siso256_1.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice0.l1  (.D(\siso256_1.tranche3.t3[1] ),
    .GATE(\siso256_1.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice0.l2  (.D(\siso256_1.tranche3.t3[2] ),
    .GATE(\siso256_1.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice0.l3  (.D(\siso256_1.tranche3.t3[3] ),
    .GATE(\siso256_1.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche3.slice1.Amp  (.Y(\siso256_1.tranche3.tranche3.slice1.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice1.l0  (.D(\siso256_1.tranche3.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice1.l1  (.D(\siso256_1.tranche3.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice1.l2  (.D(\siso256_1.tranche3.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice1.l3  (.D(\siso256_1.tranche3.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche3.slice2.Amp  (.Y(\siso256_1.tranche3.tranche3.slice2.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice2.l0  (.D(\siso256_1.tranche3.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice2.l1  (.D(\siso256_1.tranche3.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice2.l2  (.D(\siso256_1.tranche3.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice2.l3  (.D(\siso256_1.tranche3.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_1.tranche3.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_1.tranche3.tranche3.slice3.Amp  (.Y(\siso256_1.tranche3.tranche3.slice3.latch_n ),
    .A(\siso256_1.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice3.l0  (.D(\siso256_1.tranche3.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_1.tranche3.tranche3.slice3.latch_n ),
    .Q(\chain4[0] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice3.l1  (.D(\siso256_1.tranche3.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_1.tranche3.tranche3.slice3.latch_n ),
    .Q(\chain4[1] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice3.l2  (.D(\siso256_1.tranche3.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_1.tranche3.tranche3.slice3.latch_n ),
    .Q(\chain4[2] ));
 sg13g2_dlhq_1 \siso256_1.tranche3.tranche3.slice3.l3  (.D(\siso256_1.tranche3.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_1.tranche3.tranche3.slice3.latch_n ),
    .Q(\chain4[3] ));
 sg13g2_inv_4 \siso256_2.Amp0.Amp0  (.A(\Decoded8[6] ),
    .Y(\siso256_2.Amp0.Y[0] ));
 sg13g2_inv_4 \siso256_2.Amp0.Amp1  (.A(\Decoded8[4] ),
    .Y(\siso256_2.Amp0.Y[1] ));
 sg13g2_inv_4 \siso256_2.Amp0.Amp2  (.A(\Decoded8[2] ),
    .Y(\siso256_2.Amp0.Y[2] ));
 sg13g2_inv_4 \siso256_2.Amp0.Amp3  (.A(\Decoded8[0] ),
    .Y(\siso256_2.Amp0.Y[3] ));
 sg13g2_inv_1 \siso256_2.Amp1.Amp0  (.Y(\siso256_2.Amp1.Y[0] ),
    .A(\siso256_2.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_2.Amp1.Amp1  (.Y(\siso256_2.Amp1.Y[1] ),
    .A(\siso256_2.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_2.Amp1.Amp2  (.Y(\siso256_2.Amp1.Y[2] ),
    .A(\siso256_2.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_2.Amp1.Amp3  (.Y(\siso256_2.Amp1.Y[3] ),
    .A(\siso256_2.Amp0.Y[3] ));
 sg13g2_inv_1 \siso256_2.Amp2.Amp0  (.Y(\siso256_2.Amp2.Y[0] ),
    .A(\siso256_2.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_2.Amp2.Amp1  (.Y(\siso256_2.Amp2.Y[1] ),
    .A(\siso256_2.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_2.Amp2.Amp2  (.Y(\siso256_2.Amp2.Y[2] ),
    .A(\siso256_2.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_2.Amp2.Amp3  (.Y(\siso256_2.Amp2.Y[3] ),
    .A(\siso256_2.Amp0.Y[3] ));
 sg13g2_inv_1 \siso256_2.Amp3.Amp0  (.Y(\siso256_2.Amp3.Y[0] ),
    .A(\siso256_2.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_2.Amp3.Amp1  (.Y(\siso256_2.Amp3.Y[1] ),
    .A(\siso256_2.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_2.Amp3.Amp2  (.Y(\siso256_2.Amp3.Y[2] ),
    .A(\siso256_2.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_2.Amp3.Amp3  (.Y(\siso256_2.Amp3.Y[3] ),
    .A(\siso256_2.Amp0.Y[3] ));
 sg13g2_inv_1 \siso256_2.Amp4.Amp0  (.Y(\siso256_2.Amp4.Y[0] ),
    .A(\siso256_2.Amp0.Y[0] ));
 sg13g2_inv_1 \siso256_2.Amp4.Amp1  (.Y(\siso256_2.Amp4.Y[1] ),
    .A(\siso256_2.Amp0.Y[1] ));
 sg13g2_inv_1 \siso256_2.Amp4.Amp2  (.Y(\siso256_2.Amp4.Y[2] ),
    .A(\siso256_2.Amp0.Y[2] ));
 sg13g2_inv_1 \siso256_2.Amp4.Amp3  (.Y(\siso256_2.Amp4.Y[3] ),
    .A(\siso256_2.Amp0.Y[3] ));
 sg13g2_inv_2 \siso256_2.tranche0.Amp.Amp0  (.Y(\siso256_2.tranche0.tranche0.slice3.latch ),
    .A(\siso256_2.Amp1.Y[0] ));
 sg13g2_inv_2 \siso256_2.tranche0.Amp.Amp1  (.Y(\siso256_2.tranche0.tranche0.slice2.latch ),
    .A(\siso256_2.Amp1.Y[1] ));
 sg13g2_inv_2 \siso256_2.tranche0.Amp.Amp2  (.Y(\siso256_2.tranche0.tranche0.slice1.latch ),
    .A(\siso256_2.Amp1.Y[2] ));
 sg13g2_inv_2 \siso256_2.tranche0.Amp.Amp3  (.Y(\siso256_2.tranche0.tranche0.slice0.latch ),
    .A(\siso256_2.Amp1.Y[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche0.slice0.Amp  (.Y(\siso256_2.tranche0.tranche0.slice0.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice0.l0  (.D(\chain4[0] ),
    .GATE(\siso256_2.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice0.l1  (.D(\chain4[1] ),
    .GATE(\siso256_2.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice0.l2  (.D(\chain4[2] ),
    .GATE(\siso256_2.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice0.l3  (.D(\chain4[3] ),
    .GATE(\siso256_2.tranche0.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche0.slice1.Amp  (.Y(\siso256_2.tranche0.tranche0.slice1.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice1.l0  (.D(\siso256_2.tranche0.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice1.l1  (.D(\siso256_2.tranche0.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice1.l2  (.D(\siso256_2.tranche0.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice1.l3  (.D(\siso256_2.tranche0.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche0.slice2.Amp  (.Y(\siso256_2.tranche0.tranche0.slice2.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice2.l0  (.D(\siso256_2.tranche0.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice2.l1  (.D(\siso256_2.tranche0.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice2.l2  (.D(\siso256_2.tranche0.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice2.l3  (.D(\siso256_2.tranche0.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche0.slice3.Amp  (.Y(\siso256_2.tranche0.tranche0.slice3.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice3.l0  (.D(\siso256_2.tranche0.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t1[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice3.l1  (.D(\siso256_2.tranche0.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t1[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice3.l2  (.D(\siso256_2.tranche0.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t1[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche0.slice3.l3  (.D(\siso256_2.tranche0.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t1[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche1.slice0.Amp  (.Y(\siso256_2.tranche0.tranche1.slice0.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice0.l0  (.D(\siso256_2.tranche0.t1[0] ),
    .GATE(\siso256_2.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice0.l1  (.D(\siso256_2.tranche0.t1[1] ),
    .GATE(\siso256_2.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice0.l2  (.D(\siso256_2.tranche0.t1[2] ),
    .GATE(\siso256_2.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice0.l3  (.D(\siso256_2.tranche0.t1[3] ),
    .GATE(\siso256_2.tranche0.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche1.slice1.Amp  (.Y(\siso256_2.tranche0.tranche1.slice1.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice1.l0  (.D(\siso256_2.tranche0.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice1.l1  (.D(\siso256_2.tranche0.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice1.l2  (.D(\siso256_2.tranche0.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice1.l3  (.D(\siso256_2.tranche0.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche1.slice2.Amp  (.Y(\siso256_2.tranche0.tranche1.slice2.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice2.l0  (.D(\siso256_2.tranche0.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice2.l1  (.D(\siso256_2.tranche0.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice2.l2  (.D(\siso256_2.tranche0.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice2.l3  (.D(\siso256_2.tranche0.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche1.slice3.Amp  (.Y(\siso256_2.tranche0.tranche1.slice3.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice3.l0  (.D(\siso256_2.tranche0.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t2[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice3.l1  (.D(\siso256_2.tranche0.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t2[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice3.l2  (.D(\siso256_2.tranche0.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t2[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche1.slice3.l3  (.D(\siso256_2.tranche0.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t2[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche2.slice0.Amp  (.Y(\siso256_2.tranche0.tranche2.slice0.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice0.l0  (.D(\siso256_2.tranche0.t2[0] ),
    .GATE(\siso256_2.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice0.l1  (.D(\siso256_2.tranche0.t2[1] ),
    .GATE(\siso256_2.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice0.l2  (.D(\siso256_2.tranche0.t2[2] ),
    .GATE(\siso256_2.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice0.l3  (.D(\siso256_2.tranche0.t2[3] ),
    .GATE(\siso256_2.tranche0.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche2.slice1.Amp  (.Y(\siso256_2.tranche0.tranche2.slice1.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice1.l0  (.D(\siso256_2.tranche0.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice1.l1  (.D(\siso256_2.tranche0.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice1.l2  (.D(\siso256_2.tranche0.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice1.l3  (.D(\siso256_2.tranche0.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche2.slice2.Amp  (.Y(\siso256_2.tranche0.tranche2.slice2.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice2.l0  (.D(\siso256_2.tranche0.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice2.l1  (.D(\siso256_2.tranche0.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice2.l2  (.D(\siso256_2.tranche0.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice2.l3  (.D(\siso256_2.tranche0.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche2.slice3.Amp  (.Y(\siso256_2.tranche0.tranche2.slice3.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice3.l0  (.D(\siso256_2.tranche0.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t3[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice3.l1  (.D(\siso256_2.tranche0.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t3[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice3.l2  (.D(\siso256_2.tranche0.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t3[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche2.slice3.l3  (.D(\siso256_2.tranche0.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche0.t3[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche3.slice0.Amp  (.Y(\siso256_2.tranche0.tranche3.slice0.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice0.l0  (.D(\siso256_2.tranche0.t3[0] ),
    .GATE(\siso256_2.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice0.l1  (.D(\siso256_2.tranche0.t3[1] ),
    .GATE(\siso256_2.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice0.l2  (.D(\siso256_2.tranche0.t3[2] ),
    .GATE(\siso256_2.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice0.l3  (.D(\siso256_2.tranche0.t3[3] ),
    .GATE(\siso256_2.tranche0.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche3.slice1.Amp  (.Y(\siso256_2.tranche0.tranche3.slice1.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice1.l0  (.D(\siso256_2.tranche0.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice1.l1  (.D(\siso256_2.tranche0.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice1.l2  (.D(\siso256_2.tranche0.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice1.l3  (.D(\siso256_2.tranche0.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche3.slice2.Amp  (.Y(\siso256_2.tranche0.tranche3.slice2.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice2.l0  (.D(\siso256_2.tranche0.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice2.l1  (.D(\siso256_2.tranche0.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice2.l2  (.D(\siso256_2.tranche0.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice2.l3  (.D(\siso256_2.tranche0.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche0.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche0.tranche3.slice3.Amp  (.Y(\siso256_2.tranche0.tranche3.slice3.latch_n ),
    .A(\siso256_2.tranche0.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice3.l0  (.D(\siso256_2.tranche0.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t1[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice3.l1  (.D(\siso256_2.tranche0.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t1[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice3.l2  (.D(\siso256_2.tranche0.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t1[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche0.tranche3.slice3.l3  (.D(\siso256_2.tranche0.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche0.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t1[3] ));
 sg13g2_inv_2 \siso256_2.tranche1.Amp.Amp0  (.Y(\siso256_2.tranche1.tranche0.slice3.latch ),
    .A(\siso256_2.Amp2.Y[0] ));
 sg13g2_inv_2 \siso256_2.tranche1.Amp.Amp1  (.Y(\siso256_2.tranche1.tranche0.slice2.latch ),
    .A(\siso256_2.Amp2.Y[1] ));
 sg13g2_inv_2 \siso256_2.tranche1.Amp.Amp2  (.Y(\siso256_2.tranche1.tranche0.slice1.latch ),
    .A(\siso256_2.Amp2.Y[2] ));
 sg13g2_inv_2 \siso256_2.tranche1.Amp.Amp3  (.Y(\siso256_2.tranche1.tranche0.slice0.latch ),
    .A(\siso256_2.Amp2.Y[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche0.slice0.Amp  (.Y(\siso256_2.tranche1.tranche0.slice0.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice0.l0  (.D(\siso256_2.t1[0] ),
    .GATE(\siso256_2.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice0.l1  (.D(\siso256_2.t1[1] ),
    .GATE(\siso256_2.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice0.l2  (.D(\siso256_2.t1[2] ),
    .GATE(\siso256_2.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice0.l3  (.D(\siso256_2.t1[3] ),
    .GATE(\siso256_2.tranche1.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche0.slice1.Amp  (.Y(\siso256_2.tranche1.tranche0.slice1.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice1.l0  (.D(\siso256_2.tranche1.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice1.l1  (.D(\siso256_2.tranche1.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice1.l2  (.D(\siso256_2.tranche1.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice1.l3  (.D(\siso256_2.tranche1.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche0.slice2.Amp  (.Y(\siso256_2.tranche1.tranche0.slice2.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice2.l0  (.D(\siso256_2.tranche1.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice2.l1  (.D(\siso256_2.tranche1.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice2.l2  (.D(\siso256_2.tranche1.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice2.l3  (.D(\siso256_2.tranche1.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche0.slice3.Amp  (.Y(\siso256_2.tranche1.tranche0.slice3.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice3.l0  (.D(\siso256_2.tranche1.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t1[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice3.l1  (.D(\siso256_2.tranche1.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t1[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice3.l2  (.D(\siso256_2.tranche1.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t1[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche0.slice3.l3  (.D(\siso256_2.tranche1.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t1[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche1.slice0.Amp  (.Y(\siso256_2.tranche1.tranche1.slice0.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice0.l0  (.D(\siso256_2.tranche1.t1[0] ),
    .GATE(\siso256_2.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice0.l1  (.D(\siso256_2.tranche1.t1[1] ),
    .GATE(\siso256_2.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice0.l2  (.D(\siso256_2.tranche1.t1[2] ),
    .GATE(\siso256_2.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice0.l3  (.D(\siso256_2.tranche1.t1[3] ),
    .GATE(\siso256_2.tranche1.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche1.slice1.Amp  (.Y(\siso256_2.tranche1.tranche1.slice1.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice1.l0  (.D(\siso256_2.tranche1.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice1.l1  (.D(\siso256_2.tranche1.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice1.l2  (.D(\siso256_2.tranche1.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice1.l3  (.D(\siso256_2.tranche1.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche1.slice2.Amp  (.Y(\siso256_2.tranche1.tranche1.slice2.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice2.l0  (.D(\siso256_2.tranche1.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice2.l1  (.D(\siso256_2.tranche1.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice2.l2  (.D(\siso256_2.tranche1.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice2.l3  (.D(\siso256_2.tranche1.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche1.slice3.Amp  (.Y(\siso256_2.tranche1.tranche1.slice3.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice3.l0  (.D(\siso256_2.tranche1.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t2[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice3.l1  (.D(\siso256_2.tranche1.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t2[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice3.l2  (.D(\siso256_2.tranche1.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t2[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche1.slice3.l3  (.D(\siso256_2.tranche1.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t2[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche2.slice0.Amp  (.Y(\siso256_2.tranche1.tranche2.slice0.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice0.l0  (.D(\siso256_2.tranche1.t2[0] ),
    .GATE(\siso256_2.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice0.l1  (.D(\siso256_2.tranche1.t2[1] ),
    .GATE(\siso256_2.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice0.l2  (.D(\siso256_2.tranche1.t2[2] ),
    .GATE(\siso256_2.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice0.l3  (.D(\siso256_2.tranche1.t2[3] ),
    .GATE(\siso256_2.tranche1.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche2.slice1.Amp  (.Y(\siso256_2.tranche1.tranche2.slice1.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice1.l0  (.D(\siso256_2.tranche1.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice1.l1  (.D(\siso256_2.tranche1.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice1.l2  (.D(\siso256_2.tranche1.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice1.l3  (.D(\siso256_2.tranche1.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche2.slice2.Amp  (.Y(\siso256_2.tranche1.tranche2.slice2.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice2.l0  (.D(\siso256_2.tranche1.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice2.l1  (.D(\siso256_2.tranche1.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice2.l2  (.D(\siso256_2.tranche1.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice2.l3  (.D(\siso256_2.tranche1.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche2.slice3.Amp  (.Y(\siso256_2.tranche1.tranche2.slice3.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice3.l0  (.D(\siso256_2.tranche1.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t3[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice3.l1  (.D(\siso256_2.tranche1.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t3[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice3.l2  (.D(\siso256_2.tranche1.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t3[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche2.slice3.l3  (.D(\siso256_2.tranche1.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche1.t3[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche3.slice0.Amp  (.Y(\siso256_2.tranche1.tranche3.slice0.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice0.l0  (.D(\siso256_2.tranche1.t3[0] ),
    .GATE(\siso256_2.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice0.l1  (.D(\siso256_2.tranche1.t3[1] ),
    .GATE(\siso256_2.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice0.l2  (.D(\siso256_2.tranche1.t3[2] ),
    .GATE(\siso256_2.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice0.l3  (.D(\siso256_2.tranche1.t3[3] ),
    .GATE(\siso256_2.tranche1.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche3.slice1.Amp  (.Y(\siso256_2.tranche1.tranche3.slice1.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice1.l0  (.D(\siso256_2.tranche1.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice1.l1  (.D(\siso256_2.tranche1.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice1.l2  (.D(\siso256_2.tranche1.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice1.l3  (.D(\siso256_2.tranche1.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche3.slice2.Amp  (.Y(\siso256_2.tranche1.tranche3.slice2.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice2.l0  (.D(\siso256_2.tranche1.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice2.l1  (.D(\siso256_2.tranche1.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice2.l2  (.D(\siso256_2.tranche1.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice2.l3  (.D(\siso256_2.tranche1.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche1.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche1.tranche3.slice3.Amp  (.Y(\siso256_2.tranche1.tranche3.slice3.latch_n ),
    .A(\siso256_2.tranche1.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice3.l0  (.D(\siso256_2.tranche1.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t2[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice3.l1  (.D(\siso256_2.tranche1.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t2[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice3.l2  (.D(\siso256_2.tranche1.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t2[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche1.tranche3.slice3.l3  (.D(\siso256_2.tranche1.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche1.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t2[3] ));
 sg13g2_inv_2 \siso256_2.tranche2.Amp.Amp0  (.Y(\siso256_2.tranche2.tranche0.slice3.latch ),
    .A(\siso256_2.Amp3.Y[0] ));
 sg13g2_inv_2 \siso256_2.tranche2.Amp.Amp1  (.Y(\siso256_2.tranche2.tranche0.slice2.latch ),
    .A(\siso256_2.Amp3.Y[1] ));
 sg13g2_inv_2 \siso256_2.tranche2.Amp.Amp2  (.Y(\siso256_2.tranche2.tranche0.slice1.latch ),
    .A(\siso256_2.Amp3.Y[2] ));
 sg13g2_inv_2 \siso256_2.tranche2.Amp.Amp3  (.Y(\siso256_2.tranche2.tranche0.slice0.latch ),
    .A(\siso256_2.Amp3.Y[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche0.slice0.Amp  (.Y(\siso256_2.tranche2.tranche0.slice0.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice0.l0  (.D(\siso256_2.t2[0] ),
    .GATE(\siso256_2.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice0.l1  (.D(\siso256_2.t2[1] ),
    .GATE(\siso256_2.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice0.l2  (.D(\siso256_2.t2[2] ),
    .GATE(\siso256_2.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice0.l3  (.D(\siso256_2.t2[3] ),
    .GATE(\siso256_2.tranche2.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche0.slice1.Amp  (.Y(\siso256_2.tranche2.tranche0.slice1.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice1.l0  (.D(\siso256_2.tranche2.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice1.l1  (.D(\siso256_2.tranche2.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice1.l2  (.D(\siso256_2.tranche2.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice1.l3  (.D(\siso256_2.tranche2.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche0.slice2.Amp  (.Y(\siso256_2.tranche2.tranche0.slice2.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice2.l0  (.D(\siso256_2.tranche2.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice2.l1  (.D(\siso256_2.tranche2.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice2.l2  (.D(\siso256_2.tranche2.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice2.l3  (.D(\siso256_2.tranche2.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche0.slice3.Amp  (.Y(\siso256_2.tranche2.tranche0.slice3.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice3.l0  (.D(\siso256_2.tranche2.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t1[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice3.l1  (.D(\siso256_2.tranche2.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t1[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice3.l2  (.D(\siso256_2.tranche2.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t1[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche0.slice3.l3  (.D(\siso256_2.tranche2.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t1[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche1.slice0.Amp  (.Y(\siso256_2.tranche2.tranche1.slice0.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice0.l0  (.D(\siso256_2.tranche2.t1[0] ),
    .GATE(\siso256_2.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice0.l1  (.D(\siso256_2.tranche2.t1[1] ),
    .GATE(\siso256_2.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice0.l2  (.D(\siso256_2.tranche2.t1[2] ),
    .GATE(\siso256_2.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice0.l3  (.D(\siso256_2.tranche2.t1[3] ),
    .GATE(\siso256_2.tranche2.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche1.slice1.Amp  (.Y(\siso256_2.tranche2.tranche1.slice1.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice1.l0  (.D(\siso256_2.tranche2.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice1.l1  (.D(\siso256_2.tranche2.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice1.l2  (.D(\siso256_2.tranche2.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice1.l3  (.D(\siso256_2.tranche2.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche1.slice2.Amp  (.Y(\siso256_2.tranche2.tranche1.slice2.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice2.l0  (.D(\siso256_2.tranche2.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice2.l1  (.D(\siso256_2.tranche2.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice2.l2  (.D(\siso256_2.tranche2.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice2.l3  (.D(\siso256_2.tranche2.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche1.slice3.Amp  (.Y(\siso256_2.tranche2.tranche1.slice3.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice3.l0  (.D(\siso256_2.tranche2.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t2[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice3.l1  (.D(\siso256_2.tranche2.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t2[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice3.l2  (.D(\siso256_2.tranche2.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t2[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche1.slice3.l3  (.D(\siso256_2.tranche2.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t2[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche2.slice0.Amp  (.Y(\siso256_2.tranche2.tranche2.slice0.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice0.l0  (.D(\siso256_2.tranche2.t2[0] ),
    .GATE(\siso256_2.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice0.l1  (.D(\siso256_2.tranche2.t2[1] ),
    .GATE(\siso256_2.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice0.l2  (.D(\siso256_2.tranche2.t2[2] ),
    .GATE(\siso256_2.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice0.l3  (.D(\siso256_2.tranche2.t2[3] ),
    .GATE(\siso256_2.tranche2.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche2.slice1.Amp  (.Y(\siso256_2.tranche2.tranche2.slice1.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice1.l0  (.D(\siso256_2.tranche2.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice1.l1  (.D(\siso256_2.tranche2.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice1.l2  (.D(\siso256_2.tranche2.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice1.l3  (.D(\siso256_2.tranche2.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche2.slice2.Amp  (.Y(\siso256_2.tranche2.tranche2.slice2.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice2.l0  (.D(\siso256_2.tranche2.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice2.l1  (.D(\siso256_2.tranche2.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice2.l2  (.D(\siso256_2.tranche2.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice2.l3  (.D(\siso256_2.tranche2.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche2.slice3.Amp  (.Y(\siso256_2.tranche2.tranche2.slice3.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice3.l0  (.D(\siso256_2.tranche2.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t3[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice3.l1  (.D(\siso256_2.tranche2.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t3[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice3.l2  (.D(\siso256_2.tranche2.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t3[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche2.slice3.l3  (.D(\siso256_2.tranche2.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche2.t3[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche3.slice0.Amp  (.Y(\siso256_2.tranche2.tranche3.slice0.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice0.l0  (.D(\siso256_2.tranche2.t3[0] ),
    .GATE(\siso256_2.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice0.l1  (.D(\siso256_2.tranche2.t3[1] ),
    .GATE(\siso256_2.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice0.l2  (.D(\siso256_2.tranche2.t3[2] ),
    .GATE(\siso256_2.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice0.l3  (.D(\siso256_2.tranche2.t3[3] ),
    .GATE(\siso256_2.tranche2.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche3.slice1.Amp  (.Y(\siso256_2.tranche2.tranche3.slice1.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice1.l0  (.D(\siso256_2.tranche2.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice1.l1  (.D(\siso256_2.tranche2.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice1.l2  (.D(\siso256_2.tranche2.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice1.l3  (.D(\siso256_2.tranche2.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche3.slice2.Amp  (.Y(\siso256_2.tranche2.tranche3.slice2.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice2.l0  (.D(\siso256_2.tranche2.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice2.l1  (.D(\siso256_2.tranche2.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice2.l2  (.D(\siso256_2.tranche2.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice2.l3  (.D(\siso256_2.tranche2.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche2.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche2.tranche3.slice3.Amp  (.Y(\siso256_2.tranche2.tranche3.slice3.latch_n ),
    .A(\siso256_2.tranche2.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice3.l0  (.D(\siso256_2.tranche2.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t3[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice3.l1  (.D(\siso256_2.tranche2.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t3[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice3.l2  (.D(\siso256_2.tranche2.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t3[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche2.tranche3.slice3.l3  (.D(\siso256_2.tranche2.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche2.tranche3.slice3.latch_n ),
    .Q(\siso256_2.t3[3] ));
 sg13g2_inv_2 \siso256_2.tranche3.Amp.Amp0  (.Y(\siso256_2.tranche3.tranche0.slice3.latch ),
    .A(\siso256_2.Amp4.Y[0] ));
 sg13g2_inv_2 \siso256_2.tranche3.Amp.Amp1  (.Y(\siso256_2.tranche3.tranche0.slice2.latch ),
    .A(\siso256_2.Amp4.Y[1] ));
 sg13g2_inv_2 \siso256_2.tranche3.Amp.Amp2  (.Y(\siso256_2.tranche3.tranche0.slice1.latch ),
    .A(\siso256_2.Amp4.Y[2] ));
 sg13g2_inv_2 \siso256_2.tranche3.Amp.Amp3  (.Y(\siso256_2.tranche3.tranche0.slice0.latch ),
    .A(\siso256_2.Amp4.Y[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche0.slice0.Amp  (.Y(\siso256_2.tranche3.tranche0.slice0.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice0.l0  (.D(\siso256_2.t3[0] ),
    .GATE(\siso256_2.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice0.l1  (.D(\siso256_2.t3[1] ),
    .GATE(\siso256_2.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice0.l2  (.D(\siso256_2.t3[2] ),
    .GATE(\siso256_2.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice0.l3  (.D(\siso256_2.t3[3] ),
    .GATE(\siso256_2.tranche3.tranche0.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche0.slice1.Amp  (.Y(\siso256_2.tranche3.tranche0.slice1.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice1.l0  (.D(\siso256_2.tranche3.tranche0.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice1.l1  (.D(\siso256_2.tranche3.tranche0.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice1.l2  (.D(\siso256_2.tranche3.tranche0.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice1.l3  (.D(\siso256_2.tranche3.tranche0.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche0.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche0.slice2.Amp  (.Y(\siso256_2.tranche3.tranche0.slice2.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice2.l0  (.D(\siso256_2.tranche3.tranche0.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice2.l1  (.D(\siso256_2.tranche3.tranche0.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice2.l2  (.D(\siso256_2.tranche3.tranche0.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice2.l3  (.D(\siso256_2.tranche3.tranche0.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche0.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche0.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche0.slice3.Amp  (.Y(\siso256_2.tranche3.tranche0.slice3.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice3.l0  (.D(\siso256_2.tranche3.tranche0.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t1[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice3.l1  (.D(\siso256_2.tranche3.tranche0.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t1[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice3.l2  (.D(\siso256_2.tranche3.tranche0.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t1[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche0.slice3.l3  (.D(\siso256_2.tranche3.tranche0.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche0.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t1[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche1.slice0.Amp  (.Y(\siso256_2.tranche3.tranche1.slice0.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice0.l0  (.D(\siso256_2.tranche3.t1[0] ),
    .GATE(\siso256_2.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice0.l1  (.D(\siso256_2.tranche3.t1[1] ),
    .GATE(\siso256_2.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice0.l2  (.D(\siso256_2.tranche3.t1[2] ),
    .GATE(\siso256_2.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice0.l3  (.D(\siso256_2.tranche3.t1[3] ),
    .GATE(\siso256_2.tranche3.tranche1.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche1.slice1.Amp  (.Y(\siso256_2.tranche3.tranche1.slice1.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice1.l0  (.D(\siso256_2.tranche3.tranche1.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice1.l1  (.D(\siso256_2.tranche3.tranche1.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice1.l2  (.D(\siso256_2.tranche3.tranche1.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice1.l3  (.D(\siso256_2.tranche3.tranche1.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche1.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche1.slice2.Amp  (.Y(\siso256_2.tranche3.tranche1.slice2.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice2.l0  (.D(\siso256_2.tranche3.tranche1.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice2.l1  (.D(\siso256_2.tranche3.tranche1.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice2.l2  (.D(\siso256_2.tranche3.tranche1.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice2.l3  (.D(\siso256_2.tranche3.tranche1.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche1.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche1.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche1.slice3.Amp  (.Y(\siso256_2.tranche3.tranche1.slice3.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice3.l0  (.D(\siso256_2.tranche3.tranche1.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t2[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice3.l1  (.D(\siso256_2.tranche3.tranche1.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t2[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice3.l2  (.D(\siso256_2.tranche3.tranche1.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t2[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche1.slice3.l3  (.D(\siso256_2.tranche3.tranche1.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche1.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t2[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche2.slice0.Amp  (.Y(\siso256_2.tranche3.tranche2.slice0.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice0.l0  (.D(\siso256_2.tranche3.t2[0] ),
    .GATE(\siso256_2.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice0.l1  (.D(\siso256_2.tranche3.t2[1] ),
    .GATE(\siso256_2.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice0.l2  (.D(\siso256_2.tranche3.t2[2] ),
    .GATE(\siso256_2.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice0.l3  (.D(\siso256_2.tranche3.t2[3] ),
    .GATE(\siso256_2.tranche3.tranche2.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche2.slice1.Amp  (.Y(\siso256_2.tranche3.tranche2.slice1.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice1.l0  (.D(\siso256_2.tranche3.tranche2.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice1.l1  (.D(\siso256_2.tranche3.tranche2.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice1.l2  (.D(\siso256_2.tranche3.tranche2.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice1.l3  (.D(\siso256_2.tranche3.tranche2.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche2.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice1.siso_out[3] ));
 sg13g2_inv_2 \siso256_2.tranche3.tranche2.slice2.Amp  (.Y(\siso256_2.tranche3.tranche2.slice2.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice2.l0  (.D(\siso256_2.tranche3.tranche2.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice2.l1  (.D(\siso256_2.tranche3.tranche2.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice2.l2  (.D(\siso256_2.tranche3.tranche2.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice2.l3  (.D(\siso256_2.tranche3.tranche2.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche2.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche2.slice2.siso_out[3] ));
 sg13g2_inv_2 \siso256_2.tranche3.tranche2.slice3.Amp  (.Y(\siso256_2.tranche3.tranche2.slice3.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice3.l0  (.D(\siso256_2.tranche3.tranche2.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t3[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice3.l1  (.D(\siso256_2.tranche3.tranche2.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t3[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice3.l2  (.D(\siso256_2.tranche3.tranche2.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t3[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche2.slice3.l3  (.D(\siso256_2.tranche3.tranche2.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche2.slice3.latch_n ),
    .Q(\siso256_2.tranche3.t3[3] ));
 sg13g2_inv_2 \siso256_2.tranche3.tranche3.slice0.Amp  (.Y(\siso256_2.tranche3.tranche3.slice0.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice0.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice0.l0  (.D(\siso256_2.tranche3.t3[0] ),
    .GATE(\siso256_2.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice0.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice0.l1  (.D(\siso256_2.tranche3.t3[1] ),
    .GATE(\siso256_2.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice0.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice0.l2  (.D(\siso256_2.tranche3.t3[2] ),
    .GATE(\siso256_2.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice0.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice0.l3  (.D(\siso256_2.tranche3.t3[3] ),
    .GATE(\siso256_2.tranche3.tranche3.slice0.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice0.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche3.slice1.Amp  (.Y(\siso256_2.tranche3.tranche3.slice1.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice1.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice1.l0  (.D(\siso256_2.tranche3.tranche3.slice0.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice1.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice1.l1  (.D(\siso256_2.tranche3.tranche3.slice0.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice1.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice1.l2  (.D(\siso256_2.tranche3.tranche3.slice0.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice1.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice1.l3  (.D(\siso256_2.tranche3.tranche3.slice0.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche3.slice1.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice1.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche3.slice2.Amp  (.Y(\siso256_2.tranche3.tranche3.slice2.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice2.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice2.l0  (.D(\siso256_2.tranche3.tranche3.slice1.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice2.siso_out[0] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice2.l1  (.D(\siso256_2.tranche3.tranche3.slice1.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice2.siso_out[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice2.l2  (.D(\siso256_2.tranche3.tranche3.slice1.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice2.siso_out[2] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice2.l3  (.D(\siso256_2.tranche3.tranche3.slice1.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche3.slice2.latch_n ),
    .Q(\siso256_2.tranche3.tranche3.slice2.siso_out[3] ));
 sg13g2_inv_1 \siso256_2.tranche3.tranche3.slice3.Amp  (.Y(\siso256_2.tranche3.tranche3.slice3.latch_n ),
    .A(\siso256_2.tranche3.tranche0.slice3.latch ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice3.l0  (.D(\siso256_2.tranche3.tranche3.slice2.siso_out[0] ),
    .GATE(\siso256_2.tranche3.tranche3.slice3.latch_n ),
    .Q(\siso256_1.siso_in[1] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice3.l1  (.D(\siso256_2.tranche3.tranche3.slice2.siso_out[1] ),
    .GATE(\siso256_2.tranche3.tranche3.slice3.latch_n ),
    .Q(MX_out));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice3.l2  (.D(\siso256_2.tranche3.tranche3.slice2.siso_out[2] ),
    .GATE(\siso256_2.tranche3.tranche3.slice3.latch_n ),
    .Q(\siso256_1.siso_in[3] ));
 sg13g2_dlhq_1 \siso256_2.tranche3.tranche3.slice3.l3  (.D(\siso256_2.tranche3.tranche3.slice2.siso_out[3] ),
    .GATE(\siso256_2.tranche3.tranche3.slice3.latch_n ),
    .Q(DL_out));
 sg13g2_sdfrbpq_1 sync8 (.Q(back),
    .CLK(clknet_2_3__leaf_CLK_OUT_regs),
    .RESET_B(net4),
    .SCD(net34),
    .D(net36),
    .SCE(\Decoded8[5] ));
 sg13g2_sdfrbpq_1 sync_Din (.Q(SISO_in),
    .CLK(clknet_2_2__leaf_CLK_OUT_regs),
    .RESET_B(net4),
    .SCD(net35),
    .D(net7),
    .SCE(net11));
 sg13g2_buf_8 fanout3 (.A(net4),
    .X(net3));
 sg13g2_buf_8 fanout4 (.A(net37),
    .X(net4));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net5));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net6));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net7));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net8));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net9));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net10));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net11));
 sg13g2_tiehi tt_um_ygdes_hdsiso8_10 (.L_HI(net12));
 sg13g2_buf_8 clkbuf_0_CLK_OUT (.A(CLK_OUT),
    .X(clknet_0_CLK_OUT));
 sg13g2_buf_8 clkbuf_1_0__f_CLK_OUT (.A(clknet_0_CLK_OUT),
    .X(clknet_1_0__leaf_CLK_OUT));
 sg13g2_buf_8 clkbuf_0_CLK_OUT_regs (.A(CLK_OUT_regs),
    .X(clknet_0_CLK_OUT_regs));
 sg13g2_buf_8 clkbuf_2_0__f_CLK_OUT_regs (.A(clknet_0_CLK_OUT_regs),
    .X(clknet_2_0__leaf_CLK_OUT_regs));
 sg13g2_buf_8 clkbuf_2_1__f_CLK_OUT_regs (.A(clknet_0_CLK_OUT_regs),
    .X(clknet_2_1__leaf_CLK_OUT_regs));
 sg13g2_buf_8 clkbuf_2_2__f_CLK_OUT_regs (.A(clknet_0_CLK_OUT_regs),
    .X(clknet_2_2__leaf_CLK_OUT_regs));
 sg13g2_buf_8 clkbuf_2_3__f_CLK_OUT_regs (.A(clknet_0_CLK_OUT_regs),
    .X(clknet_2_3__leaf_CLK_OUT_regs));
 sg13g2_buf_1 clkload0 (.A(clknet_2_0__leaf_CLK_OUT_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_2_1__leaf_CLK_OUT_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_CLK_OUT_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\LFSR_state8[4] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold2 (.A(\LFSR_state8[6] ),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold3 (.A(\LFSR_state8[7] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold4 (.A(\LFSR_state8[2] ),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold5 (.A(\J8.J4N[3] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold6 (.A(uo_out[2]),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold7 (.A(uo_out[4]),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold8 (.A(uo_out[3]),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold9 (.A(\LFSR_state8[3] ),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold10 (.A(\lfsr.x2 ),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold11 (.A(\LFSR_state8[5] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold12 (.A(\lfsr.x1 ),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold13 (.A(\LFSR_state8[1] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold14 (.A(\lfsr.x3 ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold15 (.A(SISO_in),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold16 (.A(LFSR_BIT),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold17 (.A(back),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold18 (.A(INT_RESET),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold19 (.A(\J8.J4N[0] ),
    .X(net38));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_4 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_181 ();
 sg13g2_decap_8 FILLER_0_188 ();
 sg13g2_decap_8 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_219 ();
 sg13g2_decap_8 FILLER_0_226 ();
 sg13g2_decap_8 FILLER_0_233 ();
 sg13g2_decap_8 FILLER_0_240 ();
 sg13g2_decap_8 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_254 ();
 sg13g2_decap_8 FILLER_0_261 ();
 sg13g2_decap_8 FILLER_0_268 ();
 sg13g2_decap_8 FILLER_0_275 ();
 sg13g2_decap_8 FILLER_0_282 ();
 sg13g2_decap_8 FILLER_0_289 ();
 sg13g2_decap_8 FILLER_0_296 ();
 sg13g2_decap_8 FILLER_0_303 ();
 sg13g2_decap_8 FILLER_0_310 ();
 sg13g2_decap_8 FILLER_0_317 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_decap_8 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_338 ();
 sg13g2_decap_8 FILLER_0_345 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_4 FILLER_1_133 ();
 sg13g2_fill_1 FILLER_1_137 ();
 sg13g2_decap_8 FILLER_1_155 ();
 sg13g2_fill_2 FILLER_1_162 ();
 sg13g2_fill_1 FILLER_1_164 ();
 sg13g2_decap_8 FILLER_1_233 ();
 sg13g2_decap_8 FILLER_1_240 ();
 sg13g2_decap_8 FILLER_1_247 ();
 sg13g2_decap_8 FILLER_1_254 ();
 sg13g2_decap_8 FILLER_1_261 ();
 sg13g2_decap_8 FILLER_1_268 ();
 sg13g2_decap_8 FILLER_1_275 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_289 ();
 sg13g2_decap_8 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_fill_2 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_155 ();
 sg13g2_fill_2 FILLER_2_162 ();
 sg13g2_fill_1 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_8 FILLER_2_247 ();
 sg13g2_decap_8 FILLER_2_254 ();
 sg13g2_decap_8 FILLER_2_261 ();
 sg13g2_decap_8 FILLER_2_268 ();
 sg13g2_decap_8 FILLER_2_275 ();
 sg13g2_decap_8 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_289 ();
 sg13g2_decap_8 FILLER_2_296 ();
 sg13g2_decap_8 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_310 ();
 sg13g2_decap_8 FILLER_2_317 ();
 sg13g2_decap_8 FILLER_2_324 ();
 sg13g2_decap_8 FILLER_2_331 ();
 sg13g2_decap_8 FILLER_2_338 ();
 sg13g2_decap_8 FILLER_2_345 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_4 FILLER_3_133 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_decap_4 FILLER_3_155 ();
 sg13g2_fill_2 FILLER_3_159 ();
 sg13g2_fill_1 FILLER_3_164 ();
 sg13g2_decap_8 FILLER_3_233 ();
 sg13g2_decap_8 FILLER_3_240 ();
 sg13g2_decap_8 FILLER_3_247 ();
 sg13g2_decap_8 FILLER_3_254 ();
 sg13g2_decap_8 FILLER_3_261 ();
 sg13g2_decap_8 FILLER_3_268 ();
 sg13g2_decap_8 FILLER_3_275 ();
 sg13g2_decap_8 FILLER_3_282 ();
 sg13g2_decap_8 FILLER_3_289 ();
 sg13g2_decap_8 FILLER_3_296 ();
 sg13g2_decap_8 FILLER_3_303 ();
 sg13g2_decap_8 FILLER_3_310 ();
 sg13g2_decap_8 FILLER_3_317 ();
 sg13g2_decap_8 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_331 ();
 sg13g2_decap_8 FILLER_3_338 ();
 sg13g2_decap_8 FILLER_3_345 ();
 sg13g2_decap_8 FILLER_3_352 ();
 sg13g2_decap_8 FILLER_3_359 ();
 sg13g2_decap_8 FILLER_3_366 ();
 sg13g2_decap_8 FILLER_3_373 ();
 sg13g2_fill_1 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_398 ();
 sg13g2_decap_4 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_126 ();
 sg13g2_fill_1 FILLER_4_128 ();
 sg13g2_fill_2 FILLER_4_163 ();
 sg13g2_fill_2 FILLER_4_182 ();
 sg13g2_fill_1 FILLER_4_184 ();
 sg13g2_fill_2 FILLER_4_219 ();
 sg13g2_fill_1 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_239 ();
 sg13g2_decap_8 FILLER_4_246 ();
 sg13g2_decap_8 FILLER_4_253 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_267 ();
 sg13g2_decap_8 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_281 ();
 sg13g2_decap_8 FILLER_4_288 ();
 sg13g2_decap_8 FILLER_4_295 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_316 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_decap_8 FILLER_4_330 ();
 sg13g2_decap_8 FILLER_4_337 ();
 sg13g2_decap_8 FILLER_4_344 ();
 sg13g2_decap_8 FILLER_4_351 ();
 sg13g2_decap_8 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_365 ();
 sg13g2_decap_8 FILLER_4_372 ();
 sg13g2_fill_2 FILLER_4_379 ();
 sg13g2_decap_8 FILLER_4_398 ();
 sg13g2_decap_4 FILLER_4_405 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_fill_2 FILLER_5_126 ();
 sg13g2_fill_1 FILLER_5_128 ();
 sg13g2_fill_2 FILLER_5_163 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_fill_2 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_177 ();
 sg13g2_fill_2 FILLER_5_204 ();
 sg13g2_fill_1 FILLER_5_206 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_239 ();
 sg13g2_decap_8 FILLER_5_246 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_274 ();
 sg13g2_decap_8 FILLER_5_281 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_decap_8 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_302 ();
 sg13g2_decap_8 FILLER_5_309 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_decap_8 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_330 ();
 sg13g2_decap_8 FILLER_5_337 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_351 ();
 sg13g2_decap_8 FILLER_5_358 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_126 ();
 sg13g2_fill_1 FILLER_6_128 ();
 sg13g2_decap_8 FILLER_6_163 ();
 sg13g2_decap_4 FILLER_6_170 ();
 sg13g2_fill_1 FILLER_6_174 ();
 sg13g2_fill_2 FILLER_6_178 ();
 sg13g2_fill_1 FILLER_6_180 ();
 sg13g2_decap_8 FILLER_6_198 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_4 FILLER_6_280 ();
 sg13g2_decap_4 FILLER_6_301 ();
 sg13g2_fill_1 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_323 ();
 sg13g2_decap_8 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_fill_1 FILLER_7_128 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_fill_1 FILLER_7_165 ();
 sg13g2_decap_8 FILLER_7_206 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_fill_2 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_239 ();
 sg13g2_decap_4 FILLER_7_246 ();
 sg13g2_decap_4 FILLER_7_301 ();
 sg13g2_fill_1 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_4 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_213 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_decap_8 FILLER_8_239 ();
 sg13g2_decap_4 FILLER_8_246 ();
 sg13g2_decap_4 FILLER_8_301 ();
 sg13g2_fill_1 FILLER_8_305 ();
 sg13g2_fill_1 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_341 ();
 sg13g2_fill_1 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_4 FILLER_9_119 ();
 sg13g2_fill_2 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_142 ();
 sg13g2_decap_8 FILLER_9_169 ();
 sg13g2_fill_2 FILLER_9_176 ();
 sg13g2_fill_1 FILLER_9_178 ();
 sg13g2_decap_8 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_239 ();
 sg13g2_decap_4 FILLER_9_246 ();
 sg13g2_fill_2 FILLER_9_301 ();
 sg13g2_fill_1 FILLER_9_323 ();
 sg13g2_fill_2 FILLER_9_341 ();
 sg13g2_fill_1 FILLER_9_343 ();
 sg13g2_decap_4 FILLER_9_367 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_fill_1 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_4 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_162 ();
 sg13g2_decap_4 FILLER_10_172 ();
 sg13g2_fill_1 FILLER_10_176 ();
 sg13g2_decap_4 FILLER_10_228 ();
 sg13g2_fill_1 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_fill_2 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_4 FILLER_10_289 ();
 sg13g2_fill_1 FILLER_10_293 ();
 sg13g2_decap_8 FILLER_10_311 ();
 sg13g2_fill_2 FILLER_10_318 ();
 sg13g2_fill_1 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_fill_1 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_4 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_37 ();
 sg13g2_decap_8 FILLER_11_44 ();
 sg13g2_decap_8 FILLER_11_51 ();
 sg13g2_decap_8 FILLER_11_58 ();
 sg13g2_decap_8 FILLER_11_65 ();
 sg13g2_decap_8 FILLER_11_72 ();
 sg13g2_decap_8 FILLER_11_79 ();
 sg13g2_decap_8 FILLER_11_86 ();
 sg13g2_decap_8 FILLER_11_93 ();
 sg13g2_decap_8 FILLER_11_100 ();
 sg13g2_decap_8 FILLER_11_107 ();
 sg13g2_decap_8 FILLER_11_114 ();
 sg13g2_decap_4 FILLER_11_121 ();
 sg13g2_fill_2 FILLER_11_142 ();
 sg13g2_fill_1 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_4 FILLER_11_186 ();
 sg13g2_fill_1 FILLER_11_190 ();
 sg13g2_fill_1 FILLER_11_231 ();
 sg13g2_decap_4 FILLER_11_249 ();
 sg13g2_fill_2 FILLER_11_253 ();
 sg13g2_decap_8 FILLER_11_272 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_4 FILLER_11_320 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_decap_4 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_356 ();
 sg13g2_fill_2 FILLER_11_363 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_4 FILLER_12_14 ();
 sg13g2_fill_2 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_37 ();
 sg13g2_decap_8 FILLER_12_44 ();
 sg13g2_decap_8 FILLER_12_51 ();
 sg13g2_decap_4 FILLER_12_58 ();
 sg13g2_decap_8 FILLER_12_79 ();
 sg13g2_decap_8 FILLER_12_86 ();
 sg13g2_decap_8 FILLER_12_93 ();
 sg13g2_decap_8 FILLER_12_100 ();
 sg13g2_decap_8 FILLER_12_107 ();
 sg13g2_decap_8 FILLER_12_114 ();
 sg13g2_decap_4 FILLER_12_121 ();
 sg13g2_fill_2 FILLER_12_142 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_fill_2 FILLER_12_179 ();
 sg13g2_fill_1 FILLER_12_181 ();
 sg13g2_decap_4 FILLER_12_228 ();
 sg13g2_fill_2 FILLER_12_249 ();
 sg13g2_fill_1 FILLER_12_251 ();
 sg13g2_decap_8 FILLER_12_272 ();
 sg13g2_fill_2 FILLER_12_323 ();
 sg13g2_fill_1 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_353 ();
 sg13g2_fill_2 FILLER_12_380 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_2 ();
 sg13g2_fill_2 FILLER_13_37 ();
 sg13g2_fill_1 FILLER_13_39 ();
 sg13g2_decap_4 FILLER_13_57 ();
 sg13g2_fill_1 FILLER_13_61 ();
 sg13g2_fill_1 FILLER_13_79 ();
 sg13g2_fill_2 FILLER_13_97 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_fill_1 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_162 ();
 sg13g2_fill_2 FILLER_13_169 ();
 sg13g2_fill_1 FILLER_13_181 ();
 sg13g2_decap_4 FILLER_13_205 ();
 sg13g2_fill_2 FILLER_13_209 ();
 sg13g2_decap_4 FILLER_13_228 ();
 sg13g2_decap_4 FILLER_13_249 ();
 sg13g2_fill_2 FILLER_13_253 ();
 sg13g2_decap_4 FILLER_13_272 ();
 sg13g2_fill_2 FILLER_13_313 ();
 sg13g2_fill_2 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_decap_4 FILLER_14_57 ();
 sg13g2_fill_1 FILLER_14_61 ();
 sg13g2_fill_1 FILLER_14_79 ();
 sg13g2_fill_2 FILLER_14_97 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_decap_8 FILLER_14_153 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_4 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_decap_8 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_14_206 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_decap_4 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_4 FILLER_14_249 ();
 sg13g2_fill_2 FILLER_14_253 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_fill_2 FILLER_14_307 ();
 sg13g2_fill_1 FILLER_14_309 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_4 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_324 ();
 sg13g2_fill_2 FILLER_14_360 ();
 sg13g2_fill_1 FILLER_14_362 ();
 sg13g2_fill_2 FILLER_14_380 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_32 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_fill_2 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_59 ();
 sg13g2_decap_8 FILLER_15_128 ();
 sg13g2_fill_2 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_154 ();
 sg13g2_fill_2 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_174 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_4 FILLER_15_216 ();
 sg13g2_decap_8 FILLER_15_254 ();
 sg13g2_decap_8 FILLER_15_261 ();
 sg13g2_decap_8 FILLER_15_285 ();
 sg13g2_decap_8 FILLER_15_292 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_4 FILLER_15_320 ();
 sg13g2_fill_2 FILLER_15_324 ();
 sg13g2_decap_8 FILLER_15_360 ();
 sg13g2_decap_8 FILLER_15_367 ();
 sg13g2_fill_2 FILLER_15_374 ();
 sg13g2_decap_8 FILLER_15_393 ();
 sg13g2_decap_8 FILLER_15_400 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_14 ();
 sg13g2_fill_1 FILLER_16_32 ();
 sg13g2_decap_4 FILLER_16_36 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_fill_2 FILLER_16_74 ();
 sg13g2_fill_1 FILLER_16_76 ();
 sg13g2_decap_8 FILLER_16_128 ();
 sg13g2_fill_1 FILLER_16_135 ();
 sg13g2_fill_2 FILLER_16_153 ();
 sg13g2_fill_2 FILLER_16_172 ();
 sg13g2_fill_1 FILLER_16_174 ();
 sg13g2_decap_8 FILLER_16_209 ();
 sg13g2_fill_1 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_fill_1 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_4 FILLER_16_334 ();
 sg13g2_fill_2 FILLER_16_338 ();
 sg13g2_fill_2 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_4 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_11 ();
 sg13g2_decap_8 FILLER_17_46 ();
 sg13g2_decap_8 FILLER_17_53 ();
 sg13g2_decap_8 FILLER_17_60 ();
 sg13g2_decap_4 FILLER_17_70 ();
 sg13g2_fill_1 FILLER_17_74 ();
 sg13g2_decap_8 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_85 ();
 sg13g2_fill_1 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_91 ();
 sg13g2_fill_1 FILLER_17_93 ();
 sg13g2_decap_4 FILLER_17_131 ();
 sg13g2_fill_1 FILLER_17_135 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_174 ();
 sg13g2_decap_8 FILLER_17_195 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_fill_2 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_341 ();
 sg13g2_fill_2 FILLER_17_359 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_34 ();
 sg13g2_decap_8 FILLER_18_41 ();
 sg13g2_decap_8 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_55 ();
 sg13g2_fill_1 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_92 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_decap_4 FILLER_18_106 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_decap_8 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_143 ();
 sg13g2_fill_2 FILLER_18_153 ();
 sg13g2_decap_8 FILLER_18_192 ();
 sg13g2_decap_8 FILLER_18_199 ();
 sg13g2_decap_8 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_213 ();
 sg13g2_decap_8 FILLER_18_234 ();
 sg13g2_decap_8 FILLER_18_241 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_255 ();
 sg13g2_decap_8 FILLER_18_262 ();
 sg13g2_fill_2 FILLER_18_269 ();
 sg13g2_decap_8 FILLER_18_288 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_decap_4 FILLER_18_359 ();
 sg13g2_fill_2 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_2 FILLER_19_34 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_decap_8 FILLER_19_43 ();
 sg13g2_decap_8 FILLER_19_50 ();
 sg13g2_fill_1 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_fill_2 FILLER_19_109 ();
 sg13g2_fill_1 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_129 ();
 sg13g2_decap_8 FILLER_19_136 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_decap_8 FILLER_19_150 ();
 sg13g2_decap_8 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_164 ();
 sg13g2_fill_1 FILLER_19_183 ();
 sg13g2_decap_4 FILLER_19_187 ();
 sg13g2_fill_2 FILLER_19_191 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_251 ();
 sg13g2_decap_8 FILLER_19_258 ();
 sg13g2_decap_4 FILLER_19_265 ();
 sg13g2_fill_2 FILLER_19_269 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_4 FILLER_19_295 ();
 sg13g2_fill_1 FILLER_19_299 ();
 sg13g2_decap_4 FILLER_19_337 ();
 sg13g2_fill_1 FILLER_19_341 ();
 sg13g2_decap_8 FILLER_19_362 ();
 sg13g2_decap_8 FILLER_19_369 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_decap_8 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_48 ();
 sg13g2_fill_2 FILLER_20_55 ();
 sg13g2_fill_1 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_92 ();
 sg13g2_decap_4 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_141 ();
 sg13g2_decap_4 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_164 ();
 sg13g2_decap_8 FILLER_20_183 ();
 sg13g2_decap_8 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_197 ();
 sg13g2_decap_4 FILLER_20_204 ();
 sg13g2_fill_2 FILLER_20_208 ();
 sg13g2_decap_4 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_251 ();
 sg13g2_decap_8 FILLER_20_258 ();
 sg13g2_decap_8 FILLER_20_265 ();
 sg13g2_decap_4 FILLER_20_289 ();
 sg13g2_fill_2 FILLER_20_293 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_fill_2 FILLER_20_305 ();
 sg13g2_fill_1 FILLER_20_311 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_decap_4 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_359 ();
 sg13g2_decap_8 FILLER_20_366 ();
 sg13g2_decap_4 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_20_377 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_fill_1 FILLER_21_16 ();
 sg13g2_decap_8 FILLER_21_37 ();
 sg13g2_decap_8 FILLER_21_44 ();
 sg13g2_decap_4 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_55 ();
 sg13g2_fill_1 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_92 ();
 sg13g2_decap_4 FILLER_21_99 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_fill_2 FILLER_21_138 ();
 sg13g2_fill_2 FILLER_21_163 ();
 sg13g2_fill_1 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_251 ();
 sg13g2_decap_8 FILLER_21_258 ();
 sg13g2_decap_8 FILLER_21_265 ();
 sg13g2_fill_2 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_4 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_93 ();
 sg13g2_decap_8 FILLER_22_100 ();
 sg13g2_decap_8 FILLER_22_107 ();
 sg13g2_decap_8 FILLER_22_114 ();
 sg13g2_fill_2 FILLER_22_138 ();
 sg13g2_fill_2 FILLER_22_160 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_4 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_258 ();
 sg13g2_decap_8 FILLER_22_265 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_325 ();
 sg13g2_decap_4 FILLER_22_344 ();
 sg13g2_decap_8 FILLER_22_365 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_69 ();
 sg13g2_decap_8 FILLER_23_90 ();
 sg13g2_fill_2 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_decap_4 FILLER_23_117 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_decap_8 FILLER_23_160 ();
 sg13g2_decap_8 FILLER_23_167 ();
 sg13g2_decap_4 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_decap_8 FILLER_23_241 ();
 sg13g2_decap_8 FILLER_23_248 ();
 sg13g2_decap_8 FILLER_23_255 ();
 sg13g2_decap_8 FILLER_23_262 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_fill_2 FILLER_23_306 ();
 sg13g2_fill_2 FILLER_23_325 ();
 sg13g2_fill_1 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_43 ();
 sg13g2_fill_2 FILLER_24_50 ();
 sg13g2_decap_4 FILLER_24_69 ();
 sg13g2_fill_2 FILLER_24_90 ();
 sg13g2_fill_1 FILLER_24_92 ();
 sg13g2_decap_4 FILLER_24_120 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_4 FILLER_24_173 ();
 sg13g2_fill_2 FILLER_24_177 ();
 sg13g2_decap_4 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_4 FILLER_24_241 ();
 sg13g2_fill_1 FILLER_24_245 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_4 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_fill_2 FILLER_24_325 ();
 sg13g2_decap_4 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_decap_4 FILLER_25_46 ();
 sg13g2_fill_2 FILLER_25_50 ();
 sg13g2_decap_8 FILLER_25_86 ();
 sg13g2_decap_4 FILLER_25_93 ();
 sg13g2_decap_8 FILLER_25_117 ();
 sg13g2_decap_8 FILLER_25_124 ();
 sg13g2_fill_1 FILLER_25_131 ();
 sg13g2_decap_8 FILLER_25_155 ();
 sg13g2_decap_8 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_fill_2 FILLER_25_176 ();
 sg13g2_fill_1 FILLER_25_178 ();
 sg13g2_decap_4 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_fill_2 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_297 ();
 sg13g2_decap_4 FILLER_25_304 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_decap_8 FILLER_25_351 ();
 sg13g2_decap_4 FILLER_25_358 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_40 ();
 sg13g2_decap_8 FILLER_26_47 ();
 sg13g2_decap_8 FILLER_26_54 ();
 sg13g2_decap_8 FILLER_26_61 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_decap_8 FILLER_26_86 ();
 sg13g2_decap_8 FILLER_26_93 ();
 sg13g2_fill_1 FILLER_26_117 ();
 sg13g2_fill_1 FILLER_26_152 ();
 sg13g2_fill_2 FILLER_26_170 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_decap_4 FILLER_26_220 ();
 sg13g2_fill_2 FILLER_26_224 ();
 sg13g2_fill_1 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_4 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_8 FILLER_26_401 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_decap_8 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_50 ();
 sg13g2_fill_2 FILLER_27_89 ();
 sg13g2_fill_1 FILLER_27_117 ();
 sg13g2_fill_1 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_216 ();
 sg13g2_fill_2 FILLER_27_223 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_decap_4 FILLER_27_260 ();
 sg13g2_decap_8 FILLER_27_298 ();
 sg13g2_decap_4 FILLER_27_305 ();
 sg13g2_fill_1 FILLER_27_309 ();
 sg13g2_decap_8 FILLER_27_344 ();
 sg13g2_decap_8 FILLER_27_351 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_57 ();
 sg13g2_decap_4 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_68 ();
 sg13g2_fill_2 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_145 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_2 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_decap_8 FILLER_28_211 ();
 sg13g2_decap_4 FILLER_28_218 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_263 ();
 sg13g2_decap_4 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_278 ();
 sg13g2_decap_8 FILLER_28_296 ();
 sg13g2_decap_8 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_4 FILLER_28_317 ();
 sg13g2_fill_1 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_11 ();
 sg13g2_decap_4 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_68 ();
 sg13g2_fill_2 FILLER_29_92 ();
 sg13g2_fill_1 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_decap_8 FILLER_29_223 ();
 sg13g2_fill_2 FILLER_29_230 ();
 sg13g2_decap_8 FILLER_29_252 ();
 sg13g2_decap_8 FILLER_29_259 ();
 sg13g2_decap_8 FILLER_29_266 ();
 sg13g2_decap_4 FILLER_29_273 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_321 ();
 sg13g2_fill_1 FILLER_29_342 ();
 sg13g2_fill_1 FILLER_29_377 ();
 sg13g2_decap_8 FILLER_29_395 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_7 ();
 sg13g2_fill_1 FILLER_30_9 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_decap_8 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_decap_8 FILLER_30_237 ();
 sg13g2_decap_8 FILLER_30_244 ();
 sg13g2_fill_1 FILLER_30_271 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_4 FILLER_30_322 ();
 sg13g2_fill_1 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_9 ();
 sg13g2_decap_4 FILLER_31_47 ();
 sg13g2_decap_4 FILLER_31_54 ();
 sg13g2_fill_2 FILLER_31_58 ();
 sg13g2_fill_1 FILLER_31_111 ();
 sg13g2_fill_1 FILLER_31_125 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_398 ();
 sg13g2_decap_4 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_decap_8 FILLER_32_61 ();
 sg13g2_decap_8 FILLER_32_68 ();
 sg13g2_fill_1 FILLER_32_75 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_256 ();
 sg13g2_decap_4 FILLER_32_308 ();
 sg13g2_fill_1 FILLER_32_343 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_fill_1 FILLER_33_64 ();
 sg13g2_fill_2 FILLER_33_125 ();
 sg13g2_fill_1 FILLER_33_177 ();
 sg13g2_fill_2 FILLER_33_225 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_decap_4 FILLER_33_405 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_131 ();
 sg13g2_decap_4 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_fill_2 FILLER_34_285 ();
 sg13g2_fill_1 FILLER_34_321 ();
 sg13g2_fill_1 FILLER_34_347 ();
 sg13g2_decap_4 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_27 ();
 sg13g2_fill_2 FILLER_35_57 ();
 sg13g2_decap_8 FILLER_35_236 ();
 sg13g2_decap_4 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_247 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_9 ();
 sg13g2_fill_1 FILLER_36_185 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_fill_1 FILLER_36_308 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_155 ();
 sg13g2_fill_2 FILLER_37_232 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_decap_4 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_decap_8 FILLER_37_289 ();
 sg13g2_decap_8 FILLER_37_401 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_fill_1 FILLER_38_34 ();
 sg13g2_fill_1 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_297 ();
 sg13g2_fill_1 FILLER_38_366 ();
 assign uio_oe[0] = net12;
 assign uio_oe[1] = net13;
 assign uio_oe[2] = net14;
 assign uio_oe[3] = net15;
 assign uio_oe[4] = net16;
 assign uio_oe[5] = net17;
 assign uio_oe[6] = net18;
 assign uio_oe[7] = net19;
endmodule
