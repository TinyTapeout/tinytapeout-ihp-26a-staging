module tt_um_embeddedinn_vga (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire \frame_cnt[0] ;
 wire \frame_cnt[1] ;
 wire \frame_cnt[2] ;
 wire \frame_cnt[3] ;
 wire \frame_cnt[4] ;
 wire \frame_cnt[5] ;
 wire \frame_cnt[6] ;
 wire \frame_cnt[7] ;
 wire \frame_cnt[8] ;
 wire \frame_cnt[9] ;
 wire hsync;
 wire \hvsync_gen.display_on ;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \tx[0] ;
 wire \tx[1] ;
 wire \tx[3] ;
 wire \tx[4] ;
 wire \tx[7] ;
 wire \tx[8] ;
 wire \ty[0] ;
 wire \ty[1] ;
 wire \ty[3] ;
 wire \ty[4] ;
 wire \ty[7] ;
 wire \ty[8] ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_0_clk;
 wire x_dir;
 wire y_dir;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net1;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;

 sg13g2_inv_1 _338_ (.Y(_023_),
    .A(\tx[0] ));
 sg13g2_inv_1 _339_ (.Y(_059_),
    .A(\ty[4] ));
 sg13g2_inv_1 _340_ (.Y(_029_),
    .A(\ty[0] ));
 sg13g2_inv_1 _341_ (.Y(_060_),
    .A(\tx[3] ));
 sg13g2_inv_1 _342_ (.Y(_061_),
    .A(\tx[4] ));
 sg13g2_inv_1 _343_ (.Y(_062_),
    .A(\tx[7] ));
 sg13g2_inv_1 _344_ (.Y(_063_),
    .A(\tx[8] ));
 sg13g2_inv_1 _345_ (.Y(_064_),
    .A(net69));
 sg13g2_inv_1 _346_ (.Y(_065_),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_inv_1 _347_ (.Y(_066_),
    .A(\hvsync_gen.hpos[2] ));
 sg13g2_inv_1 _348_ (.Y(_067_),
    .A(net53));
 sg13g2_inv_1 _349_ (.Y(_013_),
    .A(\frame_cnt[0] ));
 sg13g2_inv_1 _350_ (.Y(_068_),
    .A(\frame_cnt[7] ));
 sg13g2_inv_1 _351_ (.Y(_069_),
    .A(\frame_cnt[3] ));
 sg13g2_inv_1 _352_ (.Y(_070_),
    .A(net44));
 sg13g2_inv_1 _353_ (.Y(_071_),
    .A(net46));
 sg13g2_inv_1 _354_ (.Y(_072_),
    .A(_035_));
 sg13g2_inv_1 _355_ (.Y(_073_),
    .A(_036_));
 sg13g2_inv_1 _356_ (.Y(_074_),
    .A(_038_));
 sg13g2_nand2b_1 _357_ (.Y(_075_),
    .B(net44),
    .A_N(_040_));
 sg13g2_xnor2_1 _358_ (.Y(_076_),
    .A(net44),
    .B(_040_));
 sg13g2_a21oi_1 _359_ (.A1(_059_),
    .A2(_039_),
    .Y(_077_),
    .B1(_070_));
 sg13g2_xor2_1 _360_ (.B(_039_),
    .A(net44),
    .X(_078_));
 sg13g2_xnor2_1 _361_ (.Y(_079_),
    .A(\ty[4] ),
    .B(net45));
 sg13g2_nor2_1 _362_ (.A(\ty[3] ),
    .B(net45),
    .Y(_080_));
 sg13g2_nand2_1 _363_ (.Y(_081_),
    .A(\ty[3] ),
    .B(net45));
 sg13g2_nand2_1 _364_ (.Y(_082_),
    .A(\ty[1] ),
    .B(net45));
 sg13g2_xor2_1 _365_ (.B(net45),
    .A(\ty[1] ),
    .X(_083_));
 sg13g2_nand2_1 _366_ (.Y(_084_),
    .A(\ty[0] ),
    .B(_083_));
 sg13g2_xor2_1 _367_ (.B(_038_),
    .A(net45),
    .X(_085_));
 sg13g2_a21oi_1 _368_ (.A1(_082_),
    .A2(_084_),
    .Y(_086_),
    .B1(_085_));
 sg13g2_a21oi_1 _369_ (.A1(net45),
    .A2(_074_),
    .Y(_087_),
    .B1(_086_));
 sg13g2_o21ai_1 _370_ (.B1(_081_),
    .Y(_088_),
    .A1(_080_),
    .A2(_087_));
 sg13g2_nor2b_1 _371_ (.A(_079_),
    .B_N(_088_),
    .Y(_089_));
 sg13g2_nor2b_1 _372_ (.A(_078_),
    .B_N(_089_),
    .Y(_090_));
 sg13g2_o21ai_1 _373_ (.B1(_076_),
    .Y(_091_),
    .A1(_077_),
    .A2(_090_));
 sg13g2_or3_1 _374_ (.A(_076_),
    .B(_077_),
    .C(_090_),
    .X(_092_));
 sg13g2_nand2_1 _375_ (.Y(_046_),
    .A(_091_),
    .B(_092_));
 sg13g2_a21oi_1 _376_ (.A1(\ty[4] ),
    .A2(net44),
    .Y(_093_),
    .B1(_089_));
 sg13g2_xnor2_1 _377_ (.Y(_045_),
    .A(_078_),
    .B(_093_));
 sg13g2_nand3_1 _378_ (.B(_084_),
    .C(_085_),
    .A(_082_),
    .Y(_094_));
 sg13g2_nand2b_1 _379_ (.Y(_044_),
    .B(_094_),
    .A_N(_086_));
 sg13g2_nand2b_1 _380_ (.Y(_095_),
    .B(net46),
    .A_N(_037_));
 sg13g2_xor2_1 _381_ (.B(_037_),
    .A(net46),
    .X(_096_));
 sg13g2_a21oi_1 _382_ (.A1(_061_),
    .A2(_036_),
    .Y(_097_),
    .B1(_071_));
 sg13g2_xor2_1 _383_ (.B(_036_),
    .A(net46),
    .X(_098_));
 sg13g2_xnor2_1 _384_ (.Y(_099_),
    .A(\tx[4] ),
    .B(net46));
 sg13g2_nor2_1 _385_ (.A(\tx[3] ),
    .B(net47),
    .Y(_100_));
 sg13g2_nand2_1 _386_ (.Y(_101_),
    .A(\tx[3] ),
    .B(net47));
 sg13g2_nand2_1 _387_ (.Y(_102_),
    .A(\tx[1] ),
    .B(net47));
 sg13g2_xor2_1 _388_ (.B(net47),
    .A(\tx[1] ),
    .X(_103_));
 sg13g2_nand2_1 _389_ (.Y(_104_),
    .A(\tx[0] ),
    .B(_103_));
 sg13g2_xor2_1 _390_ (.B(_035_),
    .A(net47),
    .X(_105_));
 sg13g2_a21oi_1 _391_ (.A1(_102_),
    .A2(_104_),
    .Y(_106_),
    .B1(_105_));
 sg13g2_a21oi_1 _392_ (.A1(net47),
    .A2(_072_),
    .Y(_107_),
    .B1(_106_));
 sg13g2_o21ai_1 _393_ (.B1(_101_),
    .Y(_108_),
    .A1(_100_),
    .A2(_107_));
 sg13g2_nor2b_1 _394_ (.A(_099_),
    .B_N(_108_),
    .Y(_109_));
 sg13g2_nor2b_1 _395_ (.A(_098_),
    .B_N(_109_),
    .Y(_110_));
 sg13g2_nor2_1 _396_ (.A(_097_),
    .B(_110_),
    .Y(_111_));
 sg13g2_xnor2_1 _397_ (.Y(_043_),
    .A(_096_),
    .B(_111_));
 sg13g2_a21oi_1 _398_ (.A1(\tx[4] ),
    .A2(net46),
    .Y(_112_),
    .B1(_109_));
 sg13g2_xnor2_1 _399_ (.Y(_042_),
    .A(_098_),
    .B(_112_));
 sg13g2_nand3_1 _400_ (.B(_104_),
    .C(_105_),
    .A(_102_),
    .Y(_113_));
 sg13g2_nand2b_1 _401_ (.Y(_041_),
    .B(_113_),
    .A_N(_106_));
 sg13g2_a21o_1 _402_ (.A2(\hvsync_gen.vpos[3] ),
    .A1(\hvsync_gen.vpos[2] ),
    .B1(net70),
    .X(_114_));
 sg13g2_a21oi_1 _403_ (.A1(net27),
    .A2(net38),
    .Y(_115_),
    .B1(_114_));
 sg13g2_and2_1 _404_ (.A(net66),
    .B(_114_),
    .X(_116_));
 sg13g2_nand4_1 _405_ (.B(net69),
    .C(net36),
    .A(net66),
    .Y(_117_),
    .D(net24));
 sg13g2_or4_1 _406_ (.A(net33),
    .B(_115_),
    .C(_116_),
    .D(_117_),
    .X(_012_));
 sg13g2_nor3_1 _407_ (.A(\hvsync_gen.hpos[4] ),
    .B(\hvsync_gen.hpos[5] ),
    .C(\hvsync_gen.hpos[6] ),
    .Y(_118_));
 sg13g2_nand4_1 _408_ (.B(\hvsync_gen.hpos[5] ),
    .C(net53),
    .A(\hvsync_gen.hpos[4] ),
    .Y(_119_),
    .D(\hvsync_gen.hpos[6] ));
 sg13g2_nor2_1 _409_ (.A(net18),
    .B(_118_),
    .Y(_120_));
 sg13g2_nand4_1 _410_ (.B(net20),
    .C(_119_),
    .A(net53),
    .Y(_011_),
    .D(_120_));
 sg13g2_nand2_1 _411_ (.Y(_121_),
    .A(net20),
    .B(net18));
 sg13g2_a21oi_1 _412_ (.A1(net53),
    .A2(net20),
    .Y(_122_),
    .B1(net33));
 sg13g2_and3_1 _413_ (.X(_000_),
    .A(_117_),
    .B(_121_),
    .C(_122_));
 sg13g2_and3_1 _414_ (.X(_123_),
    .A(net41),
    .B(net17),
    .C(net30));
 sg13g2_and2_1 _415_ (.A(net68),
    .B(_123_),
    .X(_124_));
 sg13g2_and2_1 _416_ (.A(net74),
    .B(_124_),
    .X(_125_));
 sg13g2_nand2_1 _417_ (.Y(_126_),
    .A(\hvsync_gen.hpos[4] ),
    .B(_124_));
 sg13g2_nor3_1 _418_ (.A(\hvsync_gen.hpos[5] ),
    .B(net53),
    .C(\hvsync_gen.hpos[6] ),
    .Y(_127_));
 sg13g2_a21oi_1 _419_ (.A1(_126_),
    .A2(_127_),
    .Y(_128_),
    .B1(_121_));
 sg13g2_inv_1 _420_ (.Y(_129_),
    .A(net43));
 sg13g2_nor2_1 _421_ (.A(net17),
    .B(net42),
    .Y(_001_));
 sg13g2_xnor2_1 _422_ (.Y(_130_),
    .A(net41),
    .B(net17));
 sg13g2_nor2_1 _423_ (.A(net42),
    .B(_130_),
    .Y(_002_));
 sg13g2_a21oi_1 _424_ (.A1(\hvsync_gen.hpos[1] ),
    .A2(net17),
    .Y(_131_),
    .B1(net30));
 sg13g2_nor3_1 _425_ (.A(_123_),
    .B(net42),
    .C(net31),
    .Y(_003_));
 sg13g2_nor2_1 _426_ (.A(net68),
    .B(_123_),
    .Y(_132_));
 sg13g2_nor3_1 _427_ (.A(_124_),
    .B(net42),
    .C(_132_),
    .Y(_004_));
 sg13g2_nor2_1 _428_ (.A(net74),
    .B(_124_),
    .Y(_133_));
 sg13g2_nor3_1 _429_ (.A(_125_),
    .B(net42),
    .C(_133_),
    .Y(_005_));
 sg13g2_and2_1 _430_ (.A(net75),
    .B(_125_),
    .X(_134_));
 sg13g2_o21ai_1 _431_ (.B1(_121_),
    .Y(_135_),
    .A1(net75),
    .A2(_125_));
 sg13g2_nor2_1 _432_ (.A(_134_),
    .B(_135_),
    .Y(_006_));
 sg13g2_and2_1 _433_ (.A(net63),
    .B(_134_),
    .X(_136_));
 sg13g2_nor2_1 _434_ (.A(net63),
    .B(_134_),
    .Y(_137_));
 sg13g2_nor3_1 _435_ (.A(net42),
    .B(_136_),
    .C(net64),
    .Y(_007_));
 sg13g2_and2_1 _436_ (.A(net22),
    .B(_136_),
    .X(_138_));
 sg13g2_nor2_1 _437_ (.A(net53),
    .B(_136_),
    .Y(_139_));
 sg13g2_nor3_1 _438_ (.A(net43),
    .B(_138_),
    .C(_139_),
    .Y(_008_));
 sg13g2_o21ai_1 _439_ (.B1(_129_),
    .Y(_140_),
    .A1(net18),
    .A2(_138_));
 sg13g2_a21oi_1 _440_ (.A1(net18),
    .A2(_138_),
    .Y(_009_),
    .B1(_140_));
 sg13g2_a21oi_1 _441_ (.A1(net18),
    .A2(_138_),
    .Y(_141_),
    .B1(net20));
 sg13g2_nor2_1 _442_ (.A(net43),
    .B(net21),
    .Y(_010_));
 sg13g2_and2_1 _443_ (.A(\hvsync_gen.vpos[5] ),
    .B(_039_),
    .X(_142_));
 sg13g2_xor2_1 _444_ (.B(_039_),
    .A(\hvsync_gen.vpos[5] ),
    .X(_143_));
 sg13g2_nand2_1 _445_ (.Y(_144_),
    .A(_059_),
    .B(\hvsync_gen.vpos[4] ));
 sg13g2_nor2b_1 _446_ (.A(\ty[3] ),
    .B_N(\hvsync_gen.vpos[3] ),
    .Y(_145_));
 sg13g2_nand2_1 _447_ (.Y(_146_),
    .A(\hvsync_gen.vpos[2] ),
    .B(_038_));
 sg13g2_nor2_1 _448_ (.A(\hvsync_gen.vpos[2] ),
    .B(_038_),
    .Y(_147_));
 sg13g2_xor2_1 _449_ (.B(_038_),
    .A(\hvsync_gen.vpos[2] ),
    .X(_148_));
 sg13g2_nand2b_1 _450_ (.Y(_149_),
    .B(\ty[1] ),
    .A_N(\hvsync_gen.vpos[1] ));
 sg13g2_nor2b_1 _451_ (.A(\ty[1] ),
    .B_N(\hvsync_gen.vpos[1] ),
    .Y(_150_));
 sg13g2_nand2b_1 _452_ (.Y(_151_),
    .B(\ty[0] ),
    .A_N(\hvsync_gen.vpos[0] ));
 sg13g2_a21oi_1 _453_ (.A1(_149_),
    .A2(_151_),
    .Y(_152_),
    .B1(_150_));
 sg13g2_o21ai_1 _454_ (.B1(_146_),
    .Y(_153_),
    .A1(_147_),
    .A2(_152_));
 sg13g2_xnor2_1 _455_ (.Y(_154_),
    .A(\ty[3] ),
    .B(\hvsync_gen.vpos[3] ));
 sg13g2_a21oi_1 _456_ (.A1(_153_),
    .A2(_154_),
    .Y(_155_),
    .B1(_145_));
 sg13g2_nor2_1 _457_ (.A(_059_),
    .B(\hvsync_gen.vpos[4] ),
    .Y(_156_));
 sg13g2_xnor2_1 _458_ (.Y(_157_),
    .A(\ty[4] ),
    .B(\hvsync_gen.vpos[4] ));
 sg13g2_o21ai_1 _459_ (.B1(_144_),
    .Y(_158_),
    .A1(_155_),
    .A2(_156_));
 sg13g2_xnor2_1 _460_ (.Y(_159_),
    .A(_143_),
    .B(_158_));
 sg13g2_xnor2_1 _461_ (.Y(_160_),
    .A(_148_),
    .B(_152_));
 sg13g2_xnor2_1 _462_ (.Y(_161_),
    .A(_155_),
    .B(_157_));
 sg13g2_xor2_1 _463_ (.B(_154_),
    .A(_153_),
    .X(_162_));
 sg13g2_nand3b_1 _464_ (.B(_161_),
    .C(_160_),
    .Y(_163_),
    .A_N(_162_));
 sg13g2_nor2b_1 _465_ (.A(_163_),
    .B_N(_159_),
    .Y(_164_));
 sg13g2_xnor2_1 _466_ (.Y(_165_),
    .A(\tx[3] ),
    .B(\hvsync_gen.hpos[3] ));
 sg13g2_xor2_1 _467_ (.B(_035_),
    .A(\hvsync_gen.hpos[2] ),
    .X(_166_));
 sg13g2_nor2b_1 _468_ (.A(\hvsync_gen.hpos[1] ),
    .B_N(\tx[1] ),
    .Y(_167_));
 sg13g2_nand2b_1 _469_ (.Y(_168_),
    .B(\hvsync_gen.hpos[1] ),
    .A_N(\tx[1] ));
 sg13g2_nor2b_1 _470_ (.A(\hvsync_gen.hpos[0] ),
    .B_N(\tx[0] ),
    .Y(_169_));
 sg13g2_o21ai_1 _471_ (.B1(_168_),
    .Y(_170_),
    .A1(_167_),
    .A2(_169_));
 sg13g2_nand2_1 _472_ (.Y(_171_),
    .A(_166_),
    .B(_170_));
 sg13g2_o21ai_1 _473_ (.B1(_171_),
    .Y(_172_),
    .A1(_066_),
    .A2(_072_));
 sg13g2_xnor2_1 _474_ (.Y(_173_),
    .A(_165_),
    .B(_172_));
 sg13g2_xor2_1 _475_ (.B(_170_),
    .A(_166_),
    .X(_174_));
 sg13g2_nor2b_1 _476_ (.A(_174_),
    .B_N(_173_),
    .Y(_175_));
 sg13g2_nand2b_2 _477_ (.Y(_176_),
    .B(_173_),
    .A_N(_174_));
 sg13g2_or2_1 _478_ (.X(_177_),
    .B(_162_),
    .A(_161_));
 sg13g2_inv_1 _479_ (.Y(_178_),
    .A(_177_));
 sg13g2_xor2_1 _480_ (.B(_160_),
    .A(_159_),
    .X(_179_));
 sg13g2_xnor2_1 _481_ (.Y(_180_),
    .A(_159_),
    .B(_160_));
 sg13g2_o21ai_1 _482_ (.B1(_176_),
    .Y(_181_),
    .A1(_177_),
    .A2(_180_));
 sg13g2_nor2_1 _483_ (.A(_164_),
    .B(_181_),
    .Y(_182_));
 sg13g2_a22oi_1 _484_ (.Y(_183_),
    .B1(\hvsync_gen.hpos[2] ),
    .B2(_035_),
    .A2(\hvsync_gen.hpos[3] ),
    .A1(_060_));
 sg13g2_a22oi_1 _485_ (.Y(_184_),
    .B1(_171_),
    .B2(_183_),
    .A2(_065_),
    .A1(\tx[3] ));
 sg13g2_nor2b_1 _486_ (.A(\tx[4] ),
    .B_N(\hvsync_gen.hpos[4] ),
    .Y(_185_));
 sg13g2_xnor2_1 _487_ (.Y(_186_),
    .A(\tx[4] ),
    .B(\hvsync_gen.hpos[4] ));
 sg13g2_xor2_1 _488_ (.B(_036_),
    .A(\hvsync_gen.hpos[5] ),
    .X(_187_));
 sg13g2_and2_1 _489_ (.A(_186_),
    .B(_187_),
    .X(_188_));
 sg13g2_o21ai_1 _490_ (.B1(_185_),
    .Y(_189_),
    .A1(\hvsync_gen.hpos[5] ),
    .A2(_036_));
 sg13g2_inv_1 _491_ (.Y(_190_),
    .A(_189_));
 sg13g2_a221oi_1 _492_ (.B2(_188_),
    .C1(_190_),
    .B1(_184_),
    .A1(\hvsync_gen.hpos[5] ),
    .Y(_191_),
    .A2(_036_));
 sg13g2_nand2_1 _493_ (.Y(_192_),
    .A(\hvsync_gen.hpos[6] ),
    .B(_037_));
 sg13g2_xnor2_1 _494_ (.Y(_193_),
    .A(\hvsync_gen.hpos[6] ),
    .B(_037_));
 sg13g2_xor2_1 _495_ (.B(_193_),
    .A(_191_),
    .X(_194_));
 sg13g2_a21oi_1 _496_ (.A1(_184_),
    .A2(_186_),
    .Y(_195_),
    .B1(_185_));
 sg13g2_xnor2_1 _497_ (.Y(_196_),
    .A(_187_),
    .B(_195_));
 sg13g2_inv_1 _498_ (.Y(_197_),
    .A(_196_));
 sg13g2_nand2_1 _499_ (.Y(_198_),
    .A(_194_),
    .B(_197_));
 sg13g2_nor2b_1 _500_ (.A(\tx[8] ),
    .B_N(\hvsync_gen.hpos[8] ),
    .Y(_199_));
 sg13g2_xnor2_1 _501_ (.Y(_200_),
    .A(\tx[8] ),
    .B(\hvsync_gen.hpos[8] ));
 sg13g2_xnor2_1 _502_ (.Y(_201_),
    .A(\tx[7] ),
    .B(net53));
 sg13g2_nand2b_1 _503_ (.Y(_202_),
    .B(_201_),
    .A_N(_193_));
 sg13g2_a21oi_1 _504_ (.A1(\tx[7] ),
    .A2(_067_),
    .Y(_203_),
    .B1(_192_));
 sg13g2_a21oi_1 _505_ (.A1(_062_),
    .A2(net53),
    .Y(_204_),
    .B1(_203_));
 sg13g2_o21ai_1 _506_ (.B1(_204_),
    .Y(_205_),
    .A1(_191_),
    .A2(_202_));
 sg13g2_xnor2_1 _507_ (.Y(_206_),
    .A(_200_),
    .B(_205_));
 sg13g2_o21ai_1 _508_ (.B1(_192_),
    .Y(_207_),
    .A1(_191_),
    .A2(_193_));
 sg13g2_xor2_1 _509_ (.B(_207_),
    .A(_201_),
    .X(_208_));
 sg13g2_nand2b_1 _510_ (.Y(_209_),
    .B(_206_),
    .A_N(_208_));
 sg13g2_xnor2_1 _511_ (.Y(_210_),
    .A(_184_),
    .B(_186_));
 sg13g2_a221oi_1 _512_ (.B2(_175_),
    .C1(_164_),
    .B1(_210_),
    .A1(_178_),
    .Y(_211_),
    .A2(_179_));
 sg13g2_nor3_1 _513_ (.A(_176_),
    .B(_210_),
    .C(_211_),
    .Y(_212_));
 sg13g2_or4_1 _514_ (.A(_182_),
    .B(_198_),
    .C(_209_),
    .D(_212_),
    .X(_213_));
 sg13g2_nor3_1 _515_ (.A(_177_),
    .B(_180_),
    .C(_210_),
    .Y(_214_));
 sg13g2_nand4_1 _516_ (.B(_198_),
    .C(_206_),
    .A(_181_),
    .Y(_215_),
    .D(_208_));
 sg13g2_or2_1 _517_ (.X(_216_),
    .B(_215_),
    .A(_214_));
 sg13g2_xnor2_1 _518_ (.Y(_217_),
    .A(_194_),
    .B(_196_));
 sg13g2_nor3_2 _519_ (.A(_206_),
    .B(_208_),
    .C(_217_),
    .Y(_218_));
 sg13g2_nor3_1 _520_ (.A(_194_),
    .B(_197_),
    .C(_209_),
    .Y(_219_));
 sg13g2_nand2_1 _521_ (.Y(_220_),
    .A(_161_),
    .B(_162_));
 sg13g2_nand2b_1 _522_ (.Y(_221_),
    .B(_210_),
    .A_N(_173_));
 sg13g2_nor2_1 _523_ (.A(_174_),
    .B(_221_),
    .Y(_222_));
 sg13g2_nand3_1 _524_ (.B(_220_),
    .C(_222_),
    .A(_159_),
    .Y(_223_));
 sg13g2_o21ai_1 _525_ (.B1(_176_),
    .Y(_224_),
    .A1(_218_),
    .A2(_223_));
 sg13g2_o21ai_1 _526_ (.B1(_224_),
    .Y(_225_),
    .A1(_218_),
    .A2(_219_));
 sg13g2_nand4_1 _527_ (.B(_197_),
    .C(_206_),
    .A(_194_),
    .Y(_226_),
    .D(_208_));
 sg13g2_nand3b_1 _528_ (.B(_217_),
    .C(_206_),
    .Y(_227_),
    .A_N(_208_));
 sg13g2_a21oi_1 _529_ (.A1(_226_),
    .A2(_227_),
    .Y(_228_),
    .B1(_211_));
 sg13g2_nor4_1 _530_ (.A(_194_),
    .B(_196_),
    .C(_206_),
    .D(_208_),
    .Y(_229_));
 sg13g2_xnor2_1 _531_ (.Y(_230_),
    .A(_173_),
    .B(_210_));
 sg13g2_xor2_1 _532_ (.B(_174_),
    .A(_160_),
    .X(_231_));
 sg13g2_xor2_1 _533_ (.B(_173_),
    .A(_162_),
    .X(_232_));
 sg13g2_xnor2_1 _534_ (.Y(_233_),
    .A(_161_),
    .B(_230_));
 sg13g2_nor2_1 _535_ (.A(_159_),
    .B(_178_),
    .Y(_234_));
 sg13g2_xor2_1 _536_ (.B(_177_),
    .A(_159_),
    .X(_235_));
 sg13g2_nor4_1 _537_ (.A(_231_),
    .B(_232_),
    .C(_233_),
    .D(_235_),
    .Y(_236_));
 sg13g2_a221oi_1 _538_ (.B2(_218_),
    .C1(_228_),
    .B1(_236_),
    .A1(_222_),
    .Y(_237_),
    .A2(_229_));
 sg13g2_and4_1 _539_ (.A(_213_),
    .B(_216_),
    .C(_225_),
    .D(_237_),
    .X(_238_));
 sg13g2_nor2b_1 _540_ (.A(\ty[8] ),
    .B_N(\hvsync_gen.vpos[8] ),
    .Y(_239_));
 sg13g2_xor2_1 _541_ (.B(\hvsync_gen.vpos[8] ),
    .A(\ty[8] ),
    .X(_240_));
 sg13g2_nor2_1 _542_ (.A(\ty[7] ),
    .B(_064_),
    .Y(_241_));
 sg13g2_xnor2_1 _543_ (.Y(_242_),
    .A(\ty[7] ),
    .B(\hvsync_gen.vpos[7] ));
 sg13g2_nand2_1 _544_ (.Y(_243_),
    .A(\hvsync_gen.vpos[6] ),
    .B(_040_));
 sg13g2_xnor2_1 _545_ (.Y(_244_),
    .A(\hvsync_gen.vpos[6] ),
    .B(_040_));
 sg13g2_a21oi_1 _546_ (.A1(_143_),
    .A2(_158_),
    .Y(_245_),
    .B1(_142_));
 sg13g2_o21ai_1 _547_ (.B1(_243_),
    .Y(_246_),
    .A1(_244_),
    .A2(_245_));
 sg13g2_a21oi_1 _548_ (.A1(_242_),
    .A2(_246_),
    .Y(_247_),
    .B1(_241_));
 sg13g2_nor2_1 _549_ (.A(_240_),
    .B(_247_),
    .Y(_248_));
 sg13g2_o21ai_1 _550_ (.B1(\hvsync_gen.vpos[9] ),
    .Y(_249_),
    .A1(_239_),
    .A2(_248_));
 sg13g2_or3_1 _551_ (.A(\hvsync_gen.vpos[9] ),
    .B(_239_),
    .C(_248_),
    .X(_250_));
 sg13g2_xnor2_1 _552_ (.Y(_251_),
    .A(_240_),
    .B(_247_));
 sg13g2_nor3_1 _553_ (.A(_206_),
    .B(_218_),
    .C(_229_),
    .Y(_252_));
 sg13g2_xor2_1 _554_ (.B(_246_),
    .A(_242_),
    .X(_253_));
 sg13g2_xor2_1 _555_ (.B(_245_),
    .A(_244_),
    .X(_254_));
 sg13g2_o21ai_1 _556_ (.B1(\hvsync_gen.display_on ),
    .Y(_255_),
    .A1(_175_),
    .A2(_210_));
 sg13g2_a21oi_1 _557_ (.A1(_200_),
    .A2(_205_),
    .Y(_256_),
    .B1(_199_));
 sg13g2_xor2_1 _558_ (.B(_256_),
    .A(\hvsync_gen.hpos[9] ),
    .X(_257_));
 sg13g2_or4_1 _559_ (.A(_234_),
    .B(_254_),
    .C(_255_),
    .D(_257_),
    .X(_258_));
 sg13g2_nor3_1 _560_ (.A(_252_),
    .B(_253_),
    .C(_258_),
    .Y(_259_));
 sg13g2_nand4_1 _561_ (.B(_250_),
    .C(_251_),
    .A(_249_),
    .Y(_260_),
    .D(_259_));
 sg13g2_nor2_2 _562_ (.A(_238_),
    .B(_260_),
    .Y(uo_out[5]));
 sg13g2_xor2_1 _563_ (.B(\frame_cnt[9] ),
    .A(\frame_cnt[4] ),
    .X(_261_));
 sg13g2_xor2_1 _564_ (.B(\hvsync_gen.hpos[4] ),
    .A(\hvsync_gen.vpos[4] ),
    .X(_262_));
 sg13g2_xnor2_1 _565_ (.Y(_263_),
    .A(_261_),
    .B(_262_));
 sg13g2_xnor2_1 _566_ (.Y(_264_),
    .A(\frame_cnt[2] ),
    .B(\frame_cnt[7] ));
 sg13g2_xor2_1 _567_ (.B(\hvsync_gen.hpos[2] ),
    .A(\hvsync_gen.vpos[2] ),
    .X(_265_));
 sg13g2_xor2_1 _568_ (.B(\frame_cnt[8] ),
    .A(\frame_cnt[3] ),
    .X(_266_));
 sg13g2_xnor2_1 _569_ (.Y(_267_),
    .A(\hvsync_gen.vpos[3] ),
    .B(\hvsync_gen.hpos[3] ));
 sg13g2_xnor2_1 _570_ (.Y(_268_),
    .A(_266_),
    .B(_267_));
 sg13g2_xnor2_1 _571_ (.Y(_269_),
    .A(\frame_cnt[1] ),
    .B(\frame_cnt[6] ));
 sg13g2_xor2_1 _572_ (.B(\hvsync_gen.hpos[1] ),
    .A(\hvsync_gen.vpos[1] ),
    .X(_270_));
 sg13g2_xnor2_1 _573_ (.Y(_271_),
    .A(_269_),
    .B(_270_));
 sg13g2_xnor2_1 _574_ (.Y(_272_),
    .A(\frame_cnt[0] ),
    .B(\frame_cnt[5] ));
 sg13g2_xor2_1 _575_ (.B(\hvsync_gen.hpos[0] ),
    .A(\hvsync_gen.vpos[0] ),
    .X(_273_));
 sg13g2_xnor2_1 _576_ (.Y(_274_),
    .A(_272_),
    .B(_273_));
 sg13g2_a21oi_1 _577_ (.A1(_264_),
    .A2(_265_),
    .Y(_275_),
    .B1(_271_));
 sg13g2_o21ai_1 _578_ (.B1(\hvsync_gen.display_on ),
    .Y(_276_),
    .A1(_264_),
    .A2(_265_));
 sg13g2_nor3_1 _579_ (.A(_268_),
    .B(_274_),
    .C(_276_),
    .Y(_277_));
 sg13g2_nand3_1 _580_ (.B(_275_),
    .C(_277_),
    .A(_263_),
    .Y(_278_));
 sg13g2_o21ai_1 _581_ (.B1(_278_),
    .Y(uo_out[0]),
    .A1(_238_),
    .A2(_260_));
 sg13g2_nand2b_1 _582_ (.Y(_279_),
    .B(\hvsync_gen.display_on ),
    .A_N(\hvsync_gen.vpos[0] ));
 sg13g2_o21ai_1 _583_ (.B1(_279_),
    .Y(uo_out[6]),
    .A1(_238_),
    .A2(_260_));
 sg13g2_nand2_1 _584_ (.Y(_280_),
    .A(\hvsync_gen.vpos[0] ),
    .B(\hvsync_gen.display_on ));
 sg13g2_o21ai_1 _585_ (.B1(_280_),
    .Y(uo_out[2]),
    .A1(_238_),
    .A2(_260_));
 sg13g2_xnor2_1 _586_ (.Y(_030_),
    .A(_029_),
    .B(_083_));
 sg13g2_nor2b_1 _587_ (.A(_080_),
    .B_N(_081_),
    .Y(_281_));
 sg13g2_xnor2_1 _588_ (.Y(_031_),
    .A(_087_),
    .B(_281_));
 sg13g2_xnor2_1 _589_ (.Y(_032_),
    .A(_079_),
    .B(_088_));
 sg13g2_nand2_1 _590_ (.Y(_282_),
    .A(\ty[7] ),
    .B(net44));
 sg13g2_or2_1 _591_ (.X(_283_),
    .B(net44),
    .A(\ty[7] ));
 sg13g2_nand2_1 _592_ (.Y(_284_),
    .A(_282_),
    .B(_283_));
 sg13g2_nand2_1 _593_ (.Y(_285_),
    .A(_075_),
    .B(_091_));
 sg13g2_xnor2_1 _594_ (.Y(_033_),
    .A(_284_),
    .B(_285_));
 sg13g2_nand4_1 _595_ (.B(_090_),
    .C(_282_),
    .A(_076_),
    .Y(_286_),
    .D(_283_));
 sg13g2_nand3_1 _596_ (.B(_282_),
    .C(_286_),
    .A(_075_),
    .Y(_287_));
 sg13g2_nor2_1 _597_ (.A(_077_),
    .B(_287_),
    .Y(_288_));
 sg13g2_xor2_1 _598_ (.B(y_dir),
    .A(\ty[8] ),
    .X(_289_));
 sg13g2_xnor2_1 _599_ (.Y(_034_),
    .A(_288_),
    .B(_289_));
 sg13g2_xor2_1 _600_ (.B(\frame_cnt[1] ),
    .A(\frame_cnt[0] ),
    .X(_014_));
 sg13g2_nand3_1 _601_ (.B(\frame_cnt[1] ),
    .C(\frame_cnt[2] ),
    .A(\frame_cnt[0] ),
    .Y(_290_));
 sg13g2_a21o_1 _602_ (.A2(\frame_cnt[1] ),
    .A1(\frame_cnt[0] ),
    .B1(\frame_cnt[2] ),
    .X(_291_));
 sg13g2_and2_1 _603_ (.A(_290_),
    .B(_291_),
    .X(_015_));
 sg13g2_nor2_2 _604_ (.A(_069_),
    .B(_290_),
    .Y(_292_));
 sg13g2_xnor2_1 _605_ (.Y(_016_),
    .A(\frame_cnt[3] ),
    .B(_290_));
 sg13g2_xor2_1 _606_ (.B(_292_),
    .A(\frame_cnt[4] ),
    .X(_017_));
 sg13g2_nand3_1 _607_ (.B(\frame_cnt[4] ),
    .C(_292_),
    .A(\frame_cnt[5] ),
    .Y(_293_));
 sg13g2_a21o_1 _608_ (.A2(_292_),
    .A1(\frame_cnt[4] ),
    .B1(\frame_cnt[5] ),
    .X(_294_));
 sg13g2_and2_1 _609_ (.A(_293_),
    .B(_294_),
    .X(_018_));
 sg13g2_nand4_1 _610_ (.B(\frame_cnt[6] ),
    .C(\frame_cnt[4] ),
    .A(\frame_cnt[5] ),
    .Y(_295_),
    .D(_292_));
 sg13g2_xnor2_1 _611_ (.Y(_019_),
    .A(\frame_cnt[6] ),
    .B(_293_));
 sg13g2_nor2_1 _612_ (.A(_068_),
    .B(_295_),
    .Y(_296_));
 sg13g2_xnor2_1 _613_ (.Y(_020_),
    .A(\frame_cnt[7] ),
    .B(_295_));
 sg13g2_nand2_1 _614_ (.Y(_297_),
    .A(\frame_cnt[8] ),
    .B(_296_));
 sg13g2_xor2_1 _615_ (.B(_296_),
    .A(\frame_cnt[8] ),
    .X(_021_));
 sg13g2_xnor2_1 _616_ (.Y(_022_),
    .A(\frame_cnt[9] ),
    .B(_297_));
 sg13g2_xnor2_1 _617_ (.Y(_024_),
    .A(_023_),
    .B(_103_));
 sg13g2_nor2b_1 _618_ (.A(_100_),
    .B_N(_101_),
    .Y(_298_));
 sg13g2_xnor2_1 _619_ (.Y(_025_),
    .A(_107_),
    .B(_298_));
 sg13g2_xnor2_1 _620_ (.Y(_026_),
    .A(_099_),
    .B(_108_));
 sg13g2_xnor2_1 _621_ (.Y(_299_),
    .A(\tx[7] ),
    .B(net46));
 sg13g2_o21ai_1 _622_ (.B1(_095_),
    .Y(_300_),
    .A1(_096_),
    .A2(_111_));
 sg13g2_xnor2_1 _623_ (.Y(_027_),
    .A(_299_),
    .B(_300_));
 sg13g2_xor2_1 _624_ (.B(net47),
    .A(\tx[8] ),
    .X(_301_));
 sg13g2_nor2_1 _625_ (.A(_096_),
    .B(_299_),
    .Y(_302_));
 sg13g2_nand2b_1 _626_ (.Y(_303_),
    .B(_095_),
    .A_N(_097_));
 sg13g2_a221oi_1 _627_ (.B2(_302_),
    .C1(_303_),
    .B1(_110_),
    .A1(\tx[7] ),
    .Y(_304_),
    .A2(net46));
 sg13g2_xnor2_1 _628_ (.Y(_028_),
    .A(_301_),
    .B(_304_));
 sg13g2_or4_1 _629_ (.A(\hvsync_gen.vpos[5] ),
    .B(\hvsync_gen.vpos[7] ),
    .C(net71),
    .D(net24),
    .X(_305_));
 sg13g2_o21ai_1 _630_ (.B1(net33),
    .Y(_306_),
    .A1(_114_),
    .A2(net72));
 sg13g2_a21oi_1 _631_ (.A1(net43),
    .A2(_306_),
    .Y(_307_),
    .B1(net35));
 sg13g2_a21oi_1 _632_ (.A1(net35),
    .A2(net43),
    .Y(_047_),
    .B1(_307_));
 sg13g2_and3_2 _633_ (.X(_308_),
    .A(net35),
    .B(net27),
    .C(net42));
 sg13g2_nor2_2 _634_ (.A(_129_),
    .B(_306_),
    .Y(_309_));
 sg13g2_a21oi_1 _635_ (.A1(\hvsync_gen.vpos[0] ),
    .A2(net42),
    .Y(_310_),
    .B1(net27));
 sg13g2_nor3_1 _636_ (.A(_308_),
    .B(_309_),
    .C(net28),
    .Y(_048_));
 sg13g2_xnor2_1 _637_ (.Y(_311_),
    .A(net73),
    .B(_308_));
 sg13g2_nor2_1 _638_ (.A(_309_),
    .B(_311_),
    .Y(_049_));
 sg13g2_a21oi_1 _639_ (.A1(\hvsync_gen.vpos[2] ),
    .A2(_308_),
    .Y(_312_),
    .B1(net38));
 sg13g2_and3_1 _640_ (.X(_313_),
    .A(net73),
    .B(net38),
    .C(_308_));
 sg13g2_nor3_1 _641_ (.A(_309_),
    .B(net39),
    .C(_313_),
    .Y(_050_));
 sg13g2_nor2_1 _642_ (.A(net70),
    .B(_313_),
    .Y(_314_));
 sg13g2_and2_1 _643_ (.A(net70),
    .B(_313_),
    .X(_315_));
 sg13g2_nor3_1 _644_ (.A(_309_),
    .B(_314_),
    .C(_315_),
    .Y(_051_));
 sg13g2_and2_1 _645_ (.A(net66),
    .B(_315_),
    .X(_316_));
 sg13g2_nor2_1 _646_ (.A(net66),
    .B(_315_),
    .Y(_317_));
 sg13g2_nor3_1 _647_ (.A(_309_),
    .B(_316_),
    .C(net67),
    .Y(_052_));
 sg13g2_nand2_1 _648_ (.Y(_318_),
    .A(net36),
    .B(_316_));
 sg13g2_inv_1 _649_ (.Y(_319_),
    .A(_318_));
 sg13g2_nand2b_1 _650_ (.Y(_320_),
    .B(_318_),
    .A_N(_309_));
 sg13g2_nor2_1 _651_ (.A(net36),
    .B(_316_),
    .Y(_321_));
 sg13g2_nor2_1 _652_ (.A(_320_),
    .B(net37),
    .Y(_053_));
 sg13g2_nand2_1 _653_ (.Y(_322_),
    .A(_064_),
    .B(_306_));
 sg13g2_a22oi_1 _654_ (.Y(_054_),
    .B1(_320_),
    .B2(_322_),
    .A2(_318_),
    .A1(_064_));
 sg13g2_a21oi_1 _655_ (.A1(\hvsync_gen.vpos[7] ),
    .A2(_319_),
    .Y(_323_),
    .B1(net24));
 sg13g2_nor2b_1 _656_ (.A(_117_),
    .B_N(_315_),
    .Y(_324_));
 sg13g2_nor3_1 _657_ (.A(_309_),
    .B(net25),
    .C(_324_),
    .Y(_055_));
 sg13g2_nor2_1 _658_ (.A(net33),
    .B(_324_),
    .Y(_325_));
 sg13g2_nor2_1 _659_ (.A(_309_),
    .B(net34),
    .Y(_056_));
 sg13g2_and2_1 _660_ (.A(\tx[0] ),
    .B(\tx[1] ),
    .X(_326_));
 sg13g2_o21ai_1 _661_ (.B1(\tx[3] ),
    .Y(_327_),
    .A1(_072_),
    .A2(_326_));
 sg13g2_nor2_1 _662_ (.A(\tx[4] ),
    .B(\tx[8] ),
    .Y(_328_));
 sg13g2_a221oi_1 _663_ (.B2(_328_),
    .C1(_100_),
    .B1(_327_),
    .A1(_061_),
    .Y(_329_),
    .A2(_071_));
 sg13g2_nor3_1 _664_ (.A(\tx[7] ),
    .B(_073_),
    .C(_329_),
    .Y(_330_));
 sg13g2_a22oi_1 _665_ (.Y(_057_),
    .B1(_037_),
    .B2(_330_),
    .A2(_071_),
    .A1(_063_));
 sg13g2_nor3_1 _666_ (.A(\ty[3] ),
    .B(\ty[4] ),
    .C(_074_),
    .Y(_331_));
 sg13g2_o21ai_1 _667_ (.B1(_040_),
    .Y(_332_),
    .A1(_039_),
    .A2(_331_));
 sg13g2_and2_1 _668_ (.A(\ty[8] ),
    .B(\ty[7] ),
    .X(_333_));
 sg13g2_a21oi_1 _669_ (.A1(\ty[1] ),
    .A2(\ty[0] ),
    .Y(_334_),
    .B1(_074_));
 sg13g2_nor3_1 _670_ (.A(\ty[4] ),
    .B(\ty[8] ),
    .C(\ty[7] ),
    .Y(_335_));
 sg13g2_nand3_1 _671_ (.B(_040_),
    .C(_335_),
    .A(_039_),
    .Y(_336_));
 sg13g2_a22oi_1 _672_ (.Y(_337_),
    .B1(_336_),
    .B2(net44),
    .A2(_333_),
    .A1(_332_));
 sg13g2_o21ai_1 _673_ (.B1(_337_),
    .Y(_058_),
    .A1(_081_),
    .A2(_334_));
 sg13g2_dfrbpq_2 _674_ (.RESET_B(net59),
    .D(_013_),
    .Q(\frame_cnt[0] ),
    .CLK(net51));
 sg13g2_dfrbpq_2 _675_ (.RESET_B(net59),
    .D(_014_),
    .Q(\frame_cnt[1] ),
    .CLK(net51));
 sg13g2_dfrbpq_2 _676_ (.RESET_B(net59),
    .D(_015_),
    .Q(\frame_cnt[2] ),
    .CLK(net51));
 sg13g2_dfrbpq_2 _677_ (.RESET_B(net54),
    .D(_016_),
    .Q(\frame_cnt[3] ),
    .CLK(net48));
 sg13g2_dfrbpq_2 _678_ (.RESET_B(net54),
    .D(_017_),
    .Q(\frame_cnt[4] ),
    .CLK(net49));
 sg13g2_dfrbpq_2 _679_ (.RESET_B(net54),
    .D(_018_),
    .Q(\frame_cnt[5] ),
    .CLK(net49));
 sg13g2_dfrbpq_2 _680_ (.RESET_B(net54),
    .D(_019_),
    .Q(\frame_cnt[6] ),
    .CLK(net48));
 sg13g2_dfrbpq_2 _681_ (.RESET_B(net54),
    .D(_020_),
    .Q(\frame_cnt[7] ),
    .CLK(net49));
 sg13g2_dfrbpq_2 _682_ (.RESET_B(net54),
    .D(_021_),
    .Q(\frame_cnt[8] ),
    .CLK(net49));
 sg13g2_dfrbpq_1 _683_ (.RESET_B(net54),
    .D(_022_),
    .Q(\frame_cnt[9] ),
    .CLK(net49));
 sg13g2_dfrbpq_1 _684_ (.RESET_B(net62),
    .D(_023_),
    .Q(\tx[0] ),
    .CLK(net51));
 sg13g2_dfrbpq_2 _685_ (.RESET_B(net62),
    .D(_024_),
    .Q(\tx[1] ),
    .CLK(net51));
 sg13g2_dfrbpq_2 _686_ (.RESET_B(net62),
    .D(_041_),
    .Q(_035_),
    .CLK(net51));
 sg13g2_dfrbpq_2 _687_ (.RESET_B(net59),
    .D(_025_),
    .Q(\tx[3] ),
    .CLK(net51));
 sg13g2_dfrbpq_2 _688_ (.RESET_B(net60),
    .D(_026_),
    .Q(\tx[4] ),
    .CLK(net51));
 sg13g2_dfrbpq_2 _689_ (.RESET_B(net60),
    .D(_042_),
    .Q(_036_),
    .CLK(net52));
 sg13g2_dfrbpq_2 _690_ (.RESET_B(net61),
    .D(_043_),
    .Q(_037_),
    .CLK(net52));
 sg13g2_dfrbpq_2 _691_ (.RESET_B(net61),
    .D(_027_),
    .Q(\tx[7] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _692_ (.RESET_B(net61),
    .D(_028_),
    .Q(\tx[8] ),
    .CLK(net52));
 sg13g2_dfrbpq_2 _693_ (.RESET_B(net55),
    .D(_029_),
    .Q(\ty[0] ),
    .CLK(net48));
 sg13g2_dfrbpq_2 _694_ (.RESET_B(net55),
    .D(_030_),
    .Q(\ty[1] ),
    .CLK(net48));
 sg13g2_dfrbpq_2 _695_ (.RESET_B(net55),
    .D(_044_),
    .Q(_038_),
    .CLK(net48));
 sg13g2_dfrbpq_2 _696_ (.RESET_B(net55),
    .D(_031_),
    .Q(\ty[3] ),
    .CLK(net48));
 sg13g2_dfrbpq_2 _697_ (.RESET_B(net55),
    .D(_032_),
    .Q(\ty[4] ),
    .CLK(net48));
 sg13g2_dfrbpq_2 _698_ (.RESET_B(net56),
    .D(_045_),
    .Q(_039_),
    .CLK(net50));
 sg13g2_dfrbpq_2 _699_ (.RESET_B(net56),
    .D(_046_),
    .Q(_040_),
    .CLK(net50));
 sg13g2_dfrbpq_2 _700_ (.RESET_B(net56),
    .D(_033_),
    .Q(\ty[7] ),
    .CLK(net50));
 sg13g2_dfrbpq_2 _701_ (.RESET_B(net56),
    .D(_034_),
    .Q(\ty[8] ),
    .CLK(net50));
 sg13g2_dfrbpq_2 _702_ (.RESET_B(net57),
    .D(_047_),
    .Q(\hvsync_gen.vpos[0] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _703_ (.RESET_B(net54),
    .D(net29),
    .Q(\hvsync_gen.vpos[1] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _704_ (.RESET_B(net58),
    .D(_049_),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _705_ (.RESET_B(net55),
    .D(net40),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _706_ (.RESET_B(net57),
    .D(_051_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _707_ (.RESET_B(net56),
    .D(_052_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _708_ (.RESET_B(net56),
    .D(_053_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _709_ (.RESET_B(net56),
    .D(_054_),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _710_ (.RESET_B(net56),
    .D(net26),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _711_ (.RESET_B(net57),
    .D(_056_),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _712_ (.RESET_B(net61),
    .D(_057_),
    .Q(x_dir),
    .CLK(net52));
 sg13g2_dfrbpq_2 _713_ (.RESET_B(net59),
    .D(_001_),
    .Q(\hvsync_gen.hpos[0] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _714_ (.RESET_B(net59),
    .D(_002_),
    .Q(\hvsync_gen.hpos[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _715_ (.RESET_B(net59),
    .D(net32),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _716_ (.RESET_B(net59),
    .D(_004_),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _717_ (.RESET_B(net60),
    .D(_005_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _718_ (.RESET_B(net60),
    .D(_006_),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _719_ (.RESET_B(net60),
    .D(net65),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _720_ (.RESET_B(net60),
    .D(_008_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _721_ (.RESET_B(net60),
    .D(net19),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _722_ (.RESET_B(net57),
    .D(_010_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _723_ (.RESET_B(net57),
    .D(_012_),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _724_ (.RESET_B(net57),
    .D(_000_),
    .Q(\hvsync_gen.display_on ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _725_ (.RESET_B(net60),
    .D(net23),
    .Q(hsync),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _726_ (.RESET_B(net55),
    .D(_058_),
    .Q(y_dir),
    .CLK(net48));
 sg13g2_tielo tt_um_embeddedinn_vga_2 (.L_LO(net2));
 sg13g2_tielo tt_um_embeddedinn_vga_3 (.L_LO(net3));
 sg13g2_tielo tt_um_embeddedinn_vga_4 (.L_LO(net4));
 sg13g2_tielo tt_um_embeddedinn_vga_5 (.L_LO(net5));
 sg13g2_tielo tt_um_embeddedinn_vga_6 (.L_LO(net6));
 sg13g2_tielo tt_um_embeddedinn_vga_7 (.L_LO(net7));
 sg13g2_tielo tt_um_embeddedinn_vga_8 (.L_LO(net8));
 sg13g2_tielo tt_um_embeddedinn_vga_9 (.L_LO(net9));
 sg13g2_tielo tt_um_embeddedinn_vga_10 (.L_LO(net10));
 sg13g2_tielo tt_um_embeddedinn_vga_11 (.L_LO(net11));
 sg13g2_tielo tt_um_embeddedinn_vga_12 (.L_LO(net12));
 sg13g2_tielo tt_um_embeddedinn_vga_13 (.L_LO(net13));
 sg13g2_tielo tt_um_embeddedinn_vga_14 (.L_LO(net14));
 sg13g2_tielo tt_um_embeddedinn_vga_15 (.L_LO(net15));
 sg13g2_tielo tt_um_embeddedinn_vga_16 (.L_LO(net16));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _743_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _744_ (.A(net50),
    .X(uo_out[3]));
 sg13g2_buf_1 _745_ (.A(uo_out[5]),
    .X(uo_out[4]));
 sg13g2_buf_1 _746_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout42 (.A(_128_),
    .X(net42));
 sg13g2_buf_1 fanout43 (.A(_128_),
    .X(net43));
 sg13g2_buf_8 fanout44 (.A(net45),
    .X(net44));
 sg13g2_buf_8 fanout45 (.A(y_dir),
    .X(net45));
 sg13g2_buf_8 fanout46 (.A(net47),
    .X(net46));
 sg13g2_buf_8 fanout47 (.A(x_dir),
    .X(net47));
 sg13g2_buf_8 fanout48 (.A(net50),
    .X(net48));
 sg13g2_buf_1 fanout49 (.A(net50),
    .X(net49));
 sg13g2_buf_8 fanout50 (.A(\hvsync_gen.vsync ),
    .X(net50));
 sg13g2_buf_8 fanout51 (.A(\hvsync_gen.vsync ),
    .X(net51));
 sg13g2_buf_1 fanout52 (.A(\hvsync_gen.vsync ),
    .X(net52));
 sg13g2_buf_8 fanout53 (.A(net22),
    .X(net53));
 sg13g2_buf_8 fanout54 (.A(net55),
    .X(net54));
 sg13g2_buf_8 fanout55 (.A(net58),
    .X(net55));
 sg13g2_buf_8 fanout56 (.A(net58),
    .X(net56));
 sg13g2_buf_8 fanout57 (.A(net58),
    .X(net57));
 sg13g2_buf_8 fanout58 (.A(rst_n),
    .X(net58));
 sg13g2_buf_8 fanout59 (.A(net62),
    .X(net59));
 sg13g2_buf_8 fanout60 (.A(net62),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(net62),
    .X(net61));
 sg13g2_buf_8 fanout62 (.A(rst_n),
    .X(net62));
 sg13g2_tielo tt_um_embeddedinn_vga_1 (.L_LO(net1));
 sg13g2_buf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hvsync_gen.hpos[0] ),
    .X(net17));
 sg13g2_dlygate4sd3_1 hold2 (.A(\hvsync_gen.hpos[8] ),
    .X(net18));
 sg13g2_dlygate4sd3_1 hold3 (.A(_009_),
    .X(net19));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.hpos[9] ),
    .X(net20));
 sg13g2_dlygate4sd3_1 hold5 (.A(_141_),
    .X(net21));
 sg13g2_dlygate4sd3_1 hold6 (.A(\hvsync_gen.hpos[7] ),
    .X(net22));
 sg13g2_dlygate4sd3_1 hold7 (.A(_011_),
    .X(net23));
 sg13g2_dlygate4sd3_1 hold8 (.A(\hvsync_gen.vpos[8] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold9 (.A(_323_),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold10 (.A(_055_),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold11 (.A(\hvsync_gen.vpos[1] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold12 (.A(_310_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold13 (.A(_048_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold14 (.A(\hvsync_gen.hpos[2] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold15 (.A(_131_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold16 (.A(_003_),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold17 (.A(\hvsync_gen.vpos[9] ),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold18 (.A(_325_),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold19 (.A(\hvsync_gen.vpos[0] ),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold20 (.A(\hvsync_gen.vpos[6] ),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold21 (.A(_321_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hvsync_gen.vpos[3] ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold23 (.A(_312_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold24 (.A(_050_),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hvsync_gen.hpos[1] ),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hvsync_gen.hpos[6] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold27 (.A(_137_),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold28 (.A(_007_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hvsync_gen.vpos[5] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold30 (.A(_317_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold31 (.A(\hvsync_gen.hpos[3] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold32 (.A(\hvsync_gen.vpos[7] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hvsync_gen.vpos[4] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hvsync_gen.vpos[6] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold35 (.A(_305_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold36 (.A(\hvsync_gen.vpos[2] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold37 (.A(\hvsync_gen.hpos[4] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold38 (.A(\hvsync_gen.hpos[5] ),
    .X(net75));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_fill_1 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_247 ();
 sg13g2_decap_8 FILLER_16_254 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_decap_8 FILLER_16_275 ();
 sg13g2_decap_8 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_289 ();
 sg13g2_decap_8 FILLER_16_296 ();
 sg13g2_decap_8 FILLER_16_303 ();
 sg13g2_decap_8 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_317 ();
 sg13g2_decap_8 FILLER_16_324 ();
 sg13g2_decap_8 FILLER_16_331 ();
 sg13g2_decap_8 FILLER_16_338 ();
 sg13g2_decap_8 FILLER_16_345 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_373 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_decap_8 FILLER_16_387 ();
 sg13g2_decap_8 FILLER_16_394 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_184 ();
 sg13g2_decap_8 FILLER_17_191 ();
 sg13g2_decap_8 FILLER_17_198 ();
 sg13g2_decap_8 FILLER_17_205 ();
 sg13g2_decap_8 FILLER_17_212 ();
 sg13g2_decap_8 FILLER_17_219 ();
 sg13g2_fill_2 FILLER_17_226 ();
 sg13g2_fill_2 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_4 FILLER_17_403 ();
 sg13g2_fill_2 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_168 ();
 sg13g2_fill_2 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_fill_2 FILLER_18_230 ();
 sg13g2_fill_1 FILLER_18_232 ();
 sg13g2_decap_8 FILLER_18_244 ();
 sg13g2_decap_8 FILLER_18_251 ();
 sg13g2_decap_8 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_265 ();
 sg13g2_decap_8 FILLER_18_272 ();
 sg13g2_decap_8 FILLER_18_279 ();
 sg13g2_decap_8 FILLER_18_286 ();
 sg13g2_decap_8 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_8 FILLER_18_349 ();
 sg13g2_decap_8 FILLER_18_356 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_370 ();
 sg13g2_decap_8 FILLER_18_377 ();
 sg13g2_decap_8 FILLER_18_384 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_153 ();
 sg13g2_decap_8 FILLER_19_160 ();
 sg13g2_fill_1 FILLER_19_167 ();
 sg13g2_decap_8 FILLER_19_183 ();
 sg13g2_fill_2 FILLER_19_190 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_210 ();
 sg13g2_fill_2 FILLER_19_264 ();
 sg13g2_decap_8 FILLER_19_279 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_fill_1 FILLER_20_91 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_decap_8 FILLER_20_131 ();
 sg13g2_decap_4 FILLER_20_138 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_decap_4 FILLER_20_171 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_2 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_fill_2 FILLER_20_252 ();
 sg13g2_fill_1 FILLER_20_254 ();
 sg13g2_decap_4 FILLER_20_263 ();
 sg13g2_fill_2 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_304 ();
 sg13g2_decap_4 FILLER_20_311 ();
 sg13g2_fill_2 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_decap_8 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_383 ();
 sg13g2_decap_8 FILLER_20_390 ();
 sg13g2_decap_8 FILLER_20_397 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_77 ();
 sg13g2_decap_4 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_110 ();
 sg13g2_decap_8 FILLER_21_129 ();
 sg13g2_decap_8 FILLER_21_136 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_8 FILLER_21_150 ();
 sg13g2_decap_8 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_fill_1 FILLER_21_176 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_decap_8 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_213 ();
 sg13g2_decap_8 FILLER_21_222 ();
 sg13g2_decap_4 FILLER_21_229 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_244 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_4 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_316 ();
 sg13g2_decap_8 FILLER_21_323 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_decap_8 FILLER_21_337 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_8 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_358 ();
 sg13g2_decap_8 FILLER_21_365 ();
 sg13g2_decap_8 FILLER_21_372 ();
 sg13g2_decap_8 FILLER_21_379 ();
 sg13g2_decap_8 FILLER_21_386 ();
 sg13g2_decap_8 FILLER_21_393 ();
 sg13g2_decap_8 FILLER_21_400 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_fill_2 FILLER_22_70 ();
 sg13g2_fill_1 FILLER_22_72 ();
 sg13g2_decap_8 FILLER_22_90 ();
 sg13g2_decap_4 FILLER_22_97 ();
 sg13g2_fill_1 FILLER_22_101 ();
 sg13g2_decap_4 FILLER_22_115 ();
 sg13g2_decap_4 FILLER_22_124 ();
 sg13g2_decap_4 FILLER_22_156 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_1 FILLER_22_220 ();
 sg13g2_fill_2 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_257 ();
 sg13g2_fill_1 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_fill_1 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_4 FILLER_22_354 ();
 sg13g2_fill_1 FILLER_22_358 ();
 sg13g2_decap_8 FILLER_22_367 ();
 sg13g2_decap_8 FILLER_22_374 ();
 sg13g2_decap_8 FILLER_22_381 ();
 sg13g2_decap_8 FILLER_22_388 ();
 sg13g2_decap_8 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_fill_1 FILLER_23_72 ();
 sg13g2_decap_8 FILLER_23_90 ();
 sg13g2_decap_8 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_104 ();
 sg13g2_fill_1 FILLER_23_106 ();
 sg13g2_decap_4 FILLER_23_120 ();
 sg13g2_decap_4 FILLER_23_137 ();
 sg13g2_fill_1 FILLER_23_141 ();
 sg13g2_decap_8 FILLER_23_166 ();
 sg13g2_decap_8 FILLER_23_201 ();
 sg13g2_fill_1 FILLER_23_208 ();
 sg13g2_decap_8 FILLER_23_226 ();
 sg13g2_decap_4 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_1 FILLER_23_265 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_fill_2 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_4 FILLER_24_63 ();
 sg13g2_fill_2 FILLER_24_136 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_decap_8 FILLER_24_163 ();
 sg13g2_fill_2 FILLER_24_170 ();
 sg13g2_fill_1 FILLER_24_172 ();
 sg13g2_decap_4 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_decap_4 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_255 ();
 sg13g2_fill_1 FILLER_24_257 ();
 sg13g2_decap_4 FILLER_24_296 ();
 sg13g2_fill_1 FILLER_24_300 ();
 sg13g2_fill_2 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_decap_4 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_349 ();
 sg13g2_decap_8 FILLER_24_356 ();
 sg13g2_decap_8 FILLER_24_363 ();
 sg13g2_decap_8 FILLER_24_370 ();
 sg13g2_decap_8 FILLER_24_377 ();
 sg13g2_decap_8 FILLER_24_384 ();
 sg13g2_decap_8 FILLER_24_391 ();
 sg13g2_decap_8 FILLER_24_398 ();
 sg13g2_decap_4 FILLER_24_405 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_4 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_87 ();
 sg13g2_decap_8 FILLER_25_94 ();
 sg13g2_decap_8 FILLER_25_101 ();
 sg13g2_decap_8 FILLER_25_113 ();
 sg13g2_decap_8 FILLER_25_120 ();
 sg13g2_decap_8 FILLER_25_127 ();
 sg13g2_decap_8 FILLER_25_134 ();
 sg13g2_decap_8 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_161 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_2 FILLER_25_211 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_decap_4 FILLER_25_302 ();
 sg13g2_fill_1 FILLER_25_306 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_decap_8 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_351 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_4 FILLER_26_63 ();
 sg13g2_fill_1 FILLER_26_67 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_fill_1 FILLER_26_110 ();
 sg13g2_decap_8 FILLER_26_122 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_1 FILLER_26_135 ();
 sg13g2_decap_8 FILLER_26_152 ();
 sg13g2_decap_4 FILLER_26_159 ();
 sg13g2_fill_2 FILLER_26_163 ();
 sg13g2_fill_1 FILLER_26_177 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_1 FILLER_26_198 ();
 sg13g2_fill_1 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_230 ();
 sg13g2_fill_1 FILLER_26_237 ();
 sg13g2_decap_4 FILLER_26_251 ();
 sg13g2_fill_1 FILLER_26_255 ();
 sg13g2_fill_1 FILLER_26_278 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_317 ();
 sg13g2_decap_4 FILLER_26_324 ();
 sg13g2_fill_1 FILLER_26_328 ();
 sg13g2_decap_4 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_fill_2 FILLER_27_70 ();
 sg13g2_fill_1 FILLER_27_72 ();
 sg13g2_decap_8 FILLER_27_86 ();
 sg13g2_decap_4 FILLER_27_93 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_decap_8 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_137 ();
 sg13g2_decap_4 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_156 ();
 sg13g2_fill_1 FILLER_27_166 ();
 sg13g2_fill_2 FILLER_27_180 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_2 FILLER_27_211 ();
 sg13g2_fill_2 FILLER_27_220 ();
 sg13g2_fill_1 FILLER_27_222 ();
 sg13g2_decap_4 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_255 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_fill_2 FILLER_27_280 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_291 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_fill_2 FILLER_27_326 ();
 sg13g2_fill_1 FILLER_27_328 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_fill_1 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_4 FILLER_28_70 ();
 sg13g2_fill_1 FILLER_28_74 ();
 sg13g2_decap_4 FILLER_28_95 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_decap_8 FILLER_28_113 ();
 sg13g2_decap_8 FILLER_28_120 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_134 ();
 sg13g2_fill_2 FILLER_28_141 ();
 sg13g2_fill_1 FILLER_28_143 ();
 sg13g2_decap_4 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_166 ();
 sg13g2_fill_1 FILLER_28_186 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_215 ();
 sg13g2_fill_2 FILLER_28_226 ();
 sg13g2_fill_2 FILLER_28_240 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_4 FILLER_28_259 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_8 FILLER_28_325 ();
 sg13g2_fill_2 FILLER_28_332 ();
 sg13g2_fill_1 FILLER_28_334 ();
 sg13g2_decap_8 FILLER_28_348 ();
 sg13g2_decap_8 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_362 ();
 sg13g2_decap_8 FILLER_28_369 ();
 sg13g2_decap_8 FILLER_28_376 ();
 sg13g2_decap_8 FILLER_28_383 ();
 sg13g2_decap_8 FILLER_28_390 ();
 sg13g2_decap_8 FILLER_28_397 ();
 sg13g2_decap_4 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_fill_2 FILLER_29_70 ();
 sg13g2_fill_1 FILLER_29_72 ();
 sg13g2_decap_8 FILLER_29_93 ();
 sg13g2_decap_8 FILLER_29_100 ();
 sg13g2_decap_8 FILLER_29_107 ();
 sg13g2_fill_2 FILLER_29_150 ();
 sg13g2_decap_8 FILLER_29_160 ();
 sg13g2_fill_2 FILLER_29_167 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_279 ();
 sg13g2_decap_8 FILLER_29_290 ();
 sg13g2_decap_4 FILLER_29_297 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_fill_2 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_fill_2 FILLER_30_70 ();
 sg13g2_fill_1 FILLER_30_72 ();
 sg13g2_decap_8 FILLER_30_90 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_128 ();
 sg13g2_fill_2 FILLER_30_142 ();
 sg13g2_fill_1 FILLER_30_144 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_fill_2 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_199 ();
 sg13g2_fill_1 FILLER_30_213 ();
 sg13g2_decap_8 FILLER_30_232 ();
 sg13g2_decap_4 FILLER_30_257 ();
 sg13g2_fill_2 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_fill_2 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_313 ();
 sg13g2_decap_8 FILLER_30_320 ();
 sg13g2_decap_4 FILLER_30_327 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_355 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_70 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_163 ();
 sg13g2_fill_2 FILLER_31_183 ();
 sg13g2_fill_2 FILLER_31_213 ();
 sg13g2_decap_4 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_247 ();
 sg13g2_fill_2 FILLER_31_254 ();
 sg13g2_fill_1 FILLER_31_265 ();
 sg13g2_decap_4 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_282 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_decap_8 FILLER_31_295 ();
 sg13g2_decap_4 FILLER_31_320 ();
 sg13g2_decap_8 FILLER_31_345 ();
 sg13g2_decap_4 FILLER_31_352 ();
 sg13g2_fill_1 FILLER_31_356 ();
 sg13g2_decap_8 FILLER_31_368 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_4 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_4 FILLER_32_105 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_133 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_4 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_233 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_258 ();
 sg13g2_fill_1 FILLER_32_260 ();
 sg13g2_decap_4 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_decap_4 FILLER_32_295 ();
 sg13g2_fill_1 FILLER_32_304 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_decap_4 FILLER_32_327 ();
 sg13g2_fill_1 FILLER_32_331 ();
 sg13g2_fill_1 FILLER_32_365 ();
 sg13g2_fill_1 FILLER_32_371 ();
 sg13g2_fill_1 FILLER_32_378 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_98 ();
 sg13g2_fill_1 FILLER_33_102 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_4 FILLER_33_226 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_decap_8 FILLER_33_235 ();
 sg13g2_fill_1 FILLER_33_242 ();
 sg13g2_decap_4 FILLER_33_271 ();
 sg13g2_fill_2 FILLER_33_275 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_decap_8 FILLER_33_314 ();
 sg13g2_decap_4 FILLER_33_321 ();
 sg13g2_fill_2 FILLER_33_334 ();
 sg13g2_decap_8 FILLER_33_349 ();
 sg13g2_decap_4 FILLER_33_356 ();
 sg13g2_decap_4 FILLER_33_373 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_247 ();
 sg13g2_fill_2 FILLER_34_261 ();
 sg13g2_decap_8 FILLER_34_289 ();
 sg13g2_fill_1 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_309 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_decap_4 FILLER_35_149 ();
 sg13g2_fill_2 FILLER_35_153 ();
 sg13g2_decap_4 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_173 ();
 sg13g2_decap_4 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_fill_1 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_216 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_4 FILLER_35_228 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_decap_4 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_247 ();
 sg13g2_fill_1 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_316 ();
 sg13g2_decap_8 FILLER_35_323 ();
 sg13g2_decap_8 FILLER_35_342 ();
 sg13g2_decap_8 FILLER_35_349 ();
 sg13g2_decap_8 FILLER_35_356 ();
 sg13g2_decap_8 FILLER_35_363 ();
 sg13g2_decap_8 FILLER_35_370 ();
 sg13g2_fill_2 FILLER_35_377 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_fill_2 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_decap_4 FILLER_36_241 ();
 sg13g2_fill_1 FILLER_36_245 ();
 sg13g2_fill_1 FILLER_36_265 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_316 ();
 sg13g2_decap_8 FILLER_36_323 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_decap_8 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_344 ();
 sg13g2_decap_8 FILLER_36_374 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_8 FILLER_36_388 ();
 sg13g2_decap_8 FILLER_36_395 ();
 sg13g2_decap_8 FILLER_36_402 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_203 ();
 sg13g2_decap_4 FILLER_37_219 ();
 sg13g2_decap_8 FILLER_37_232 ();
 sg13g2_decap_4 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_249 ();
 sg13g2_fill_2 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_4 FILLER_38_201 ();
 sg13g2_fill_2 FILLER_38_205 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_1 FILLER_38_264 ();
 sg13g2_fill_2 FILLER_38_293 ();
 sg13g2_fill_1 FILLER_38_295 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net11;
 assign uio_out[3] = net12;
 assign uio_out[4] = net13;
 assign uio_out[5] = net14;
 assign uio_out[6] = net15;
 assign uio_out[7] = net16;
endmodule
