module tt_um_arthfink_ddmtd (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire clk_fb;
 wire clk_helper;
 wire \ctrl[10] ;
 wire \ctrl[11] ;
 wire \ctrl[12] ;
 wire \ctrl[13] ;
 wire \ctrl[14] ;
 wire \ctrl[15] ;
 wire \ctrl[16] ;
 wire \ctrl[17] ;
 wire \ctrl[18] ;
 wire \ctrl[19] ;
 wire \ctrl[20] ;
 wire \ctrl[21] ;
 wire \ctrl[22] ;
 wire \ctrl[23] ;
 wire \ctrl[8] ;
 wire \ctrl[9] ;
 wire fb_samp;
 wire helper_msb_d;
 wire \nco_phase_acc[0] ;
 wire \nco_phase_acc[10] ;
 wire \nco_phase_acc[11] ;
 wire \nco_phase_acc[12] ;
 wire \nco_phase_acc[13] ;
 wire \nco_phase_acc[14] ;
 wire \nco_phase_acc[15] ;
 wire \nco_phase_acc[16] ;
 wire \nco_phase_acc[17] ;
 wire \nco_phase_acc[18] ;
 wire \nco_phase_acc[19] ;
 wire \nco_phase_acc[1] ;
 wire \nco_phase_acc[20] ;
 wire \nco_phase_acc[21] ;
 wire \nco_phase_acc[22] ;
 wire \nco_phase_acc[2] ;
 wire \nco_phase_acc[3] ;
 wire \nco_phase_acc[4] ;
 wire \nco_phase_acc[5] ;
 wire \nco_phase_acc[6] ;
 wire \nco_phase_acc[7] ;
 wire \nco_phase_acc[8] ;
 wire \nco_phase_acc[9] ;
 wire \phase_err_beat[10] ;
 wire \phase_err_beat[11] ;
 wire \phase_err_beat[12] ;
 wire \phase_err_beat[13] ;
 wire \phase_err_beat[14] ;
 wire \phase_err_beat[15] ;
 wire \phase_err_beat[3] ;
 wire \phase_err_beat[4] ;
 wire \phase_err_beat[5] ;
 wire \phase_err_beat[6] ;
 wire \phase_err_beat[7] ;
 wire \phase_err_beat[8] ;
 wire \phase_err_beat[9] ;
 wire phase_valid;
 wire ref_samp;
 wire \u_core.beat_cnt[0] ;
 wire \u_core.beat_cnt[10] ;
 wire \u_core.beat_cnt[11] ;
 wire \u_core.beat_cnt[12] ;
 wire \u_core.beat_cnt[13] ;
 wire \u_core.beat_cnt[14] ;
 wire \u_core.beat_cnt[15] ;
 wire \u_core.beat_cnt[1] ;
 wire \u_core.beat_cnt[2] ;
 wire \u_core.beat_cnt[3] ;
 wire \u_core.beat_cnt[4] ;
 wire \u_core.beat_cnt[5] ;
 wire \u_core.beat_cnt[6] ;
 wire \u_core.beat_cnt[7] ;
 wire \u_core.beat_cnt[8] ;
 wire \u_core.beat_cnt[9] ;
 wire \u_core.fb_samp_d ;
 wire \u_core.fb_sync[0] ;
 wire \u_core.fb_sync[1] ;
 wire \u_core.have_fb ;
 wire \u_core.have_ref ;
 wire \u_core.ref_samp_d ;
 wire \u_core.ref_sync[0] ;
 wire \u_core.ref_sync[1] ;
 wire \u_core.t_fb[0] ;
 wire \u_core.t_fb[10] ;
 wire \u_core.t_fb[11] ;
 wire \u_core.t_fb[12] ;
 wire \u_core.t_fb[13] ;
 wire \u_core.t_fb[14] ;
 wire \u_core.t_fb[15] ;
 wire \u_core.t_fb[1] ;
 wire \u_core.t_fb[2] ;
 wire \u_core.t_fb[3] ;
 wire \u_core.t_fb[4] ;
 wire \u_core.t_fb[5] ;
 wire \u_core.t_fb[6] ;
 wire \u_core.t_fb[7] ;
 wire \u_core.t_fb[8] ;
 wire \u_core.t_fb[9] ;
 wire \u_core.t_ref[0] ;
 wire \u_core.t_ref[10] ;
 wire \u_core.t_ref[11] ;
 wire \u_core.t_ref[12] ;
 wire \u_core.t_ref[13] ;
 wire \u_core.t_ref[14] ;
 wire \u_core.t_ref[15] ;
 wire \u_core.t_ref[1] ;
 wire \u_core.t_ref[2] ;
 wire \u_core.t_ref[3] ;
 wire \u_core.t_ref[4] ;
 wire \u_core.t_ref[5] ;
 wire \u_core.t_ref[6] ;
 wire \u_core.t_ref[7] ;
 wire \u_core.t_ref[8] ;
 wire \u_core.t_ref[9] ;
 wire \u_lf.i_acc[0] ;
 wire \u_lf.i_acc[10] ;
 wire \u_lf.i_acc[11] ;
 wire \u_lf.i_acc[12] ;
 wire \u_lf.i_acc[13] ;
 wire \u_lf.i_acc[14] ;
 wire \u_lf.i_acc[15] ;
 wire \u_lf.i_acc[16] ;
 wire \u_lf.i_acc[17] ;
 wire \u_lf.i_acc[18] ;
 wire \u_lf.i_acc[19] ;
 wire \u_lf.i_acc[1] ;
 wire \u_lf.i_acc[20] ;
 wire \u_lf.i_acc[21] ;
 wire \u_lf.i_acc[22] ;
 wire \u_lf.i_acc[23] ;
 wire \u_lf.i_acc[24] ;
 wire \u_lf.i_acc[25] ;
 wire \u_lf.i_acc[26] ;
 wire \u_lf.i_acc[27] ;
 wire \u_lf.i_acc[28] ;
 wire \u_lf.i_acc[29] ;
 wire \u_lf.i_acc[2] ;
 wire \u_lf.i_acc[3] ;
 wire \u_lf.i_acc[4] ;
 wire \u_lf.i_acc[5] ;
 wire \u_lf.i_acc[6] ;
 wire \u_lf.i_acc[7] ;
 wire \u_lf.i_acc[8] ;
 wire \u_lf.i_acc[9] ;
 wire \u_lf.ki_sel_latched[0] ;
 wire \u_lf.kp_sel_latched[0] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire clknet_0_clk;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;

 sg13g2_inv_1 _0718_ (.Y(_0153_),
    .A(net205));
 sg13g2_inv_1 _0719_ (.Y(_0154_),
    .A(net113));
 sg13g2_inv_1 _0720_ (.Y(_0155_),
    .A(net56));
 sg13g2_inv_2 _0721_ (.Y(_0156_),
    .A(net199));
 sg13g2_inv_1 _0722_ (.Y(_0157_),
    .A(net206));
 sg13g2_inv_1 _0723_ (.Y(_0158_),
    .A(net325));
 sg13g2_inv_1 _0724_ (.Y(_0159_),
    .A(net246));
 sg13g2_inv_1 _0725_ (.Y(_0160_),
    .A(net280));
 sg13g2_inv_1 _0726_ (.Y(_0161_),
    .A(net155));
 sg13g2_inv_1 _0727_ (.Y(_0162_),
    .A(net150));
 sg13g2_inv_1 _0728_ (.Y(_0163_),
    .A(net46));
 sg13g2_inv_1 _0729_ (.Y(_0164_),
    .A(net44));
 sg13g2_inv_1 _0730_ (.Y(_0165_),
    .A(net129));
 sg13g2_inv_1 _0731_ (.Y(_0166_),
    .A(net87));
 sg13g2_inv_1 _0732_ (.Y(_0167_),
    .A(net123));
 sg13g2_inv_1 _0733_ (.Y(_0168_),
    .A(net127));
 sg13g2_inv_1 _0734_ (.Y(_0169_),
    .A(net77));
 sg13g2_inv_1 _0735_ (.Y(_0170_),
    .A(net138));
 sg13g2_inv_1 _0736_ (.Y(_0171_),
    .A(net268));
 sg13g2_inv_1 _0737_ (.Y(_0172_),
    .A(net110));
 sg13g2_inv_1 _0738_ (.Y(_0173_),
    .A(net135));
 sg13g2_inv_1 _0739_ (.Y(_0174_),
    .A(net102));
 sg13g2_inv_1 _0740_ (.Y(_0175_),
    .A(net318));
 sg13g2_inv_1 _0741_ (.Y(_0176_),
    .A(net287));
 sg13g2_inv_1 _0742_ (.Y(_0177_),
    .A(net324));
 sg13g2_inv_1 _0743_ (.Y(_0178_),
    .A(\nco_phase_acc[9] ));
 sg13g2_inv_1 _0744_ (.Y(_0179_),
    .A(net260));
 sg13g2_inv_1 _0745_ (.Y(_0180_),
    .A(net96));
 sg13g2_inv_1 _0746_ (.Y(_0181_),
    .A(net115));
 sg13g2_inv_1 _0747_ (.Y(_0182_),
    .A(net316));
 sg13g2_inv_1 _0748_ (.Y(_0183_),
    .A(\nco_phase_acc[13] ));
 sg13g2_inv_1 _0749_ (.Y(_0184_),
    .A(net152));
 sg13g2_o21ai_1 _0750_ (.B1(net240),
    .Y(_0185_),
    .A1(helper_msb_d),
    .A2(net26));
 sg13g2_a21oi_2 _0751_ (.B1(_0185_),
    .Y(_0186_),
    .A2(net26),
    .A1(helper_msb_d));
 sg13g2_inv_2 _0752_ (.Y(_0187_),
    .A(net186));
 sg13g2_nand3_1 _0753_ (.B(net261),
    .C(net186),
    .A(net300),
    .Y(_0188_));
 sg13g2_inv_1 _0754_ (.Y(_0000_),
    .A(net176));
 sg13g2_nand2_1 _0755_ (.Y(_0189_),
    .A(net239),
    .B(net271));
 sg13g2_inv_1 _0756_ (.Y(net184),
    .A(net188));
 sg13g2_mux2_1 _0757_ (.A0(net2),
    .A1(net26),
    .S(net3),
    .X(clk_fb));
 sg13g2_and2_1 _0758_ (.A(net239),
    .B(net200),
    .X(uo_out[1]));
 sg13g2_and2_1 _0759_ (.A(net239),
    .B(\phase_err_beat[6] ),
    .X(uo_out[2]));
 sg13g2_and2_1 _0760_ (.A(net239),
    .B(\phase_err_beat[7] ),
    .X(uo_out[3]));
 sg13g2_and2_1 _0761_ (.A(net239),
    .B(\phase_err_beat[8] ),
    .X(uo_out[4]));
 sg13g2_and2_1 _0762_ (.A(net239),
    .B(\phase_err_beat[9] ),
    .X(uo_out[5]));
 sg13g2_and2_1 _0763_ (.A(net239),
    .B(\phase_err_beat[10] ),
    .X(uo_out[6]));
 sg13g2_and2_1 _0764_ (.A(net242),
    .B(net203),
    .X(uo_out[7]));
 sg13g2_nand2_1 _0765_ (.Y(_0190_),
    .A(net240),
    .B(\ctrl[8] ));
 sg13g2_xnor2_1 _0766_ (.Y(_0003_),
    .A(net32),
    .B(_0190_));
 sg13g2_nor2_1 _0767_ (.A(net240),
    .B(net121),
    .Y(_0191_));
 sg13g2_nand2_1 _0768_ (.Y(_0192_),
    .A(net87),
    .B(net32));
 sg13g2_nand2_1 _0769_ (.Y(_0193_),
    .A(\ctrl[9] ),
    .B(\nco_phase_acc[1] ));
 sg13g2_xnor2_1 _0770_ (.Y(_0194_),
    .A(\ctrl[9] ),
    .B(net121));
 sg13g2_xnor2_1 _0771_ (.Y(_0195_),
    .A(_0192_),
    .B(_0194_));
 sg13g2_a21oi_1 _0772_ (.A1(net240),
    .A2(_0195_),
    .Y(_0004_),
    .B1(_0191_));
 sg13g2_nor2_1 _0773_ (.A(net240),
    .B(net79),
    .Y(_0196_));
 sg13g2_and2_1 _0774_ (.A(\ctrl[10] ),
    .B(net79),
    .X(_0197_));
 sg13g2_xor2_1 _0775_ (.B(net79),
    .A(\ctrl[10] ),
    .X(_0198_));
 sg13g2_o21ai_1 _0776_ (.B1(_0193_),
    .Y(_0199_),
    .A1(_0192_),
    .A2(_0194_));
 sg13g2_xnor2_1 _0777_ (.Y(_0200_),
    .A(_0198_),
    .B(_0199_));
 sg13g2_a21oi_1 _0778_ (.A1(net240),
    .A2(_0200_),
    .Y(_0005_),
    .B1(_0196_));
 sg13g2_nor2_1 _0779_ (.A(net237),
    .B(net100),
    .Y(_0201_));
 sg13g2_nand2_1 _0780_ (.Y(_0202_),
    .A(\ctrl[11] ),
    .B(\nco_phase_acc[3] ));
 sg13g2_xnor2_1 _0781_ (.Y(_0203_),
    .A(\ctrl[11] ),
    .B(net100));
 sg13g2_a21oi_1 _0782_ (.A1(_0198_),
    .A2(_0199_),
    .Y(_0204_),
    .B1(_0197_));
 sg13g2_xnor2_1 _0783_ (.Y(_0205_),
    .A(_0203_),
    .B(_0204_));
 sg13g2_a21oi_1 _0784_ (.A1(net237),
    .A2(_0205_),
    .Y(_0006_),
    .B1(_0201_));
 sg13g2_and2_1 _0785_ (.A(net77),
    .B(net94),
    .X(_0206_));
 sg13g2_or2_1 _0786_ (.X(_0207_),
    .B(net94),
    .A(net77));
 sg13g2_nor2b_1 _0787_ (.A(_0206_),
    .B_N(_0207_),
    .Y(_0208_));
 sg13g2_o21ai_1 _0788_ (.B1(_0202_),
    .Y(_0209_),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_xnor2_1 _0789_ (.Y(_0210_),
    .A(_0208_),
    .B(_0209_));
 sg13g2_nor2_1 _0790_ (.A(net237),
    .B(net94),
    .Y(_0211_));
 sg13g2_a21oi_1 _0791_ (.A1(net238),
    .A2(_0210_),
    .Y(_0007_),
    .B1(_0211_));
 sg13g2_nor2_1 _0792_ (.A(net238),
    .B(net117),
    .Y(_0212_));
 sg13g2_a21oi_1 _0793_ (.A1(_0207_),
    .A2(_0209_),
    .Y(_0213_),
    .B1(_0206_));
 sg13g2_nor2_1 _0794_ (.A(\ctrl[13] ),
    .B(\nco_phase_acc[5] ),
    .Y(_0214_));
 sg13g2_xnor2_1 _0795_ (.Y(_0215_),
    .A(\ctrl[13] ),
    .B(net117));
 sg13g2_xnor2_1 _0796_ (.Y(_0216_),
    .A(_0213_),
    .B(_0215_));
 sg13g2_a21oi_1 _0797_ (.A1(net238),
    .A2(_0216_),
    .Y(_0008_),
    .B1(_0212_));
 sg13g2_nand2_1 _0798_ (.Y(_0217_),
    .A(\ctrl[14] ),
    .B(\nco_phase_acc[6] ));
 sg13g2_xnor2_1 _0799_ (.Y(_0218_),
    .A(\ctrl[14] ),
    .B(net110));
 sg13g2_a221oi_1 _0800_ (.B2(_0209_),
    .C1(_0206_),
    .B1(_0208_),
    .A1(\ctrl[13] ),
    .Y(_0219_),
    .A2(\nco_phase_acc[5] ));
 sg13g2_or3_1 _0801_ (.A(_0214_),
    .B(_0218_),
    .C(_0219_),
    .X(_0220_));
 sg13g2_o21ai_1 _0802_ (.B1(_0218_),
    .Y(_0221_),
    .A1(_0214_),
    .A2(_0219_));
 sg13g2_nand3_1 _0803_ (.B(_0220_),
    .C(_0221_),
    .A(net237),
    .Y(_0222_));
 sg13g2_o21ai_1 _0804_ (.B1(_0222_),
    .Y(_0009_),
    .A1(net237),
    .A2(_0172_));
 sg13g2_nand2_1 _0805_ (.Y(_0223_),
    .A(net135),
    .B(net102));
 sg13g2_xnor2_1 _0806_ (.Y(_0224_),
    .A(\ctrl[15] ),
    .B(net102));
 sg13g2_a21o_1 _0807_ (.A2(_0220_),
    .A1(_0217_),
    .B1(_0224_),
    .X(_0225_));
 sg13g2_nand3_1 _0808_ (.B(_0220_),
    .C(_0224_),
    .A(_0217_),
    .Y(_0226_));
 sg13g2_nand3_1 _0809_ (.B(_0225_),
    .C(_0226_),
    .A(net237),
    .Y(_0227_));
 sg13g2_o21ai_1 _0810_ (.B1(_0227_),
    .Y(_0010_),
    .A1(net237),
    .A2(_0174_));
 sg13g2_xnor2_1 _0811_ (.Y(_0228_),
    .A(\ctrl[16] ),
    .B(net287));
 sg13g2_a21o_2 _0812_ (.A2(_0225_),
    .A1(_0223_),
    .B1(_0228_),
    .X(_0229_));
 sg13g2_nand3_1 _0813_ (.B(_0225_),
    .C(_0228_),
    .A(_0223_),
    .Y(_0230_));
 sg13g2_nand3_1 _0814_ (.B(_0229_),
    .C(_0230_),
    .A(net235),
    .Y(_0231_));
 sg13g2_o21ai_1 _0815_ (.B1(_0231_),
    .Y(_0011_),
    .A1(net235),
    .A2(_0176_));
 sg13g2_nor2_1 _0816_ (.A(net235),
    .B(net251),
    .Y(_0232_));
 sg13g2_xor2_1 _0817_ (.B(net251),
    .A(\ctrl[17] ),
    .X(_0233_));
 sg13g2_o21ai_1 _0818_ (.B1(_0229_),
    .Y(_0234_),
    .A1(_0175_),
    .A2(_0176_));
 sg13g2_xnor2_1 _0819_ (.Y(_0235_),
    .A(_0233_),
    .B(_0234_));
 sg13g2_a21oi_1 _0820_ (.A1(net235),
    .A2(_0235_),
    .Y(_0012_),
    .B1(_0232_));
 sg13g2_nand2_1 _0821_ (.Y(_0236_),
    .A(\ctrl[18] ),
    .B(net83));
 sg13g2_xor2_1 _0822_ (.B(net83),
    .A(\ctrl[18] ),
    .X(_0237_));
 sg13g2_a22oi_1 _0823_ (.Y(_0238_),
    .B1(\ctrl[17] ),
    .B2(\nco_phase_acc[9] ),
    .A2(\nco_phase_acc[8] ),
    .A1(\ctrl[16] ));
 sg13g2_a22oi_1 _0824_ (.Y(_0239_),
    .B1(_0229_),
    .B2(_0238_),
    .A2(_0178_),
    .A1(_0177_));
 sg13g2_nand2_1 _0825_ (.Y(_0240_),
    .A(_0237_),
    .B(_0239_));
 sg13g2_xnor2_1 _0826_ (.Y(_0241_),
    .A(_0237_),
    .B(_0239_));
 sg13g2_nor2_1 _0827_ (.A(net234),
    .B(net83),
    .Y(_0242_));
 sg13g2_a21oi_1 _0828_ (.A1(net234),
    .A2(_0241_),
    .Y(_0013_),
    .B1(_0242_));
 sg13g2_nor2_1 _0829_ (.A(net96),
    .B(net133),
    .Y(_0243_));
 sg13g2_nand2_1 _0830_ (.Y(_0244_),
    .A(net96),
    .B(\nco_phase_acc[11] ));
 sg13g2_nor2b_1 _0831_ (.A(_0243_),
    .B_N(_0244_),
    .Y(_0245_));
 sg13g2_nand2_1 _0832_ (.Y(_0246_),
    .A(_0236_),
    .B(_0240_));
 sg13g2_xnor2_1 _0833_ (.Y(_0247_),
    .A(_0245_),
    .B(_0246_));
 sg13g2_nor2_1 _0834_ (.A(net234),
    .B(net133),
    .Y(_0248_));
 sg13g2_a21oi_1 _0835_ (.A1(net234),
    .A2(_0247_),
    .Y(_0014_),
    .B1(_0248_));
 sg13g2_nor2_1 _0836_ (.A(net234),
    .B(net92),
    .Y(_0249_));
 sg13g2_nand2_1 _0837_ (.Y(_0250_),
    .A(_0237_),
    .B(_0245_));
 sg13g2_a221oi_1 _0838_ (.B2(_0238_),
    .C1(_0250_),
    .B1(_0229_),
    .A1(_0177_),
    .Y(_0251_),
    .A2(_0178_));
 sg13g2_o21ai_1 _0839_ (.B1(_0244_),
    .Y(_0252_),
    .A1(_0236_),
    .A2(_0243_));
 sg13g2_nor2_1 _0840_ (.A(_0251_),
    .B(_0252_),
    .Y(_0253_));
 sg13g2_nand2_1 _0841_ (.Y(_0254_),
    .A(net115),
    .B(net92));
 sg13g2_xnor2_1 _0842_ (.Y(_0255_),
    .A(\ctrl[20] ),
    .B(net92));
 sg13g2_xnor2_1 _0843_ (.Y(_0256_),
    .A(_0253_),
    .B(_0255_));
 sg13g2_a21oi_1 _0844_ (.A1(net234),
    .A2(_0256_),
    .Y(_0015_),
    .B1(_0249_));
 sg13g2_xor2_1 _0845_ (.B(net144),
    .A(\ctrl[21] ),
    .X(_0257_));
 sg13g2_o21ai_1 _0846_ (.B1(_0254_),
    .Y(_0258_),
    .A1(_0253_),
    .A2(_0255_));
 sg13g2_o21ai_1 _0847_ (.B1(net234),
    .Y(_0259_),
    .A1(_0257_),
    .A2(_0258_));
 sg13g2_a21oi_1 _0848_ (.A1(_0257_),
    .A2(_0258_),
    .Y(_0260_),
    .B1(_0259_));
 sg13g2_nand2b_1 _0849_ (.Y(_0261_),
    .B(net144),
    .A_N(net234));
 sg13g2_nand2b_1 _0850_ (.Y(_0016_),
    .B(_0261_),
    .A_N(_0260_));
 sg13g2_nor2_1 _0851_ (.A(net236),
    .B(net90),
    .Y(_0262_));
 sg13g2_nor2b_1 _0852_ (.A(_0255_),
    .B_N(_0257_),
    .Y(_0263_));
 sg13g2_o21ai_1 _0853_ (.B1(_0263_),
    .Y(_0264_),
    .A1(_0251_),
    .A2(_0252_));
 sg13g2_a21oi_1 _0854_ (.A1(_0182_),
    .A2(_0183_),
    .Y(_0265_),
    .B1(_0254_));
 sg13g2_a21oi_1 _0855_ (.A1(\ctrl[21] ),
    .A2(\nco_phase_acc[13] ),
    .Y(_0266_),
    .B1(_0265_));
 sg13g2_nand2_1 _0856_ (.Y(_0267_),
    .A(_0264_),
    .B(_0266_));
 sg13g2_nand2_1 _0857_ (.Y(_0268_),
    .A(\ctrl[22] ),
    .B(\nco_phase_acc[14] ));
 sg13g2_xor2_1 _0858_ (.B(net90),
    .A(\ctrl[22] ),
    .X(_0269_));
 sg13g2_nand2_1 _0859_ (.Y(_0270_),
    .A(_0267_),
    .B(_0269_));
 sg13g2_xnor2_1 _0860_ (.Y(_0271_),
    .A(_0267_),
    .B(_0269_));
 sg13g2_a21oi_1 _0861_ (.A1(net236),
    .A2(_0271_),
    .Y(_0017_),
    .B1(_0262_));
 sg13g2_and2_1 _0862_ (.A(_0268_),
    .B(_0270_),
    .X(_0272_));
 sg13g2_nor2_1 _0863_ (.A(\ctrl[23] ),
    .B(net73),
    .Y(_0273_));
 sg13g2_nand2_1 _0864_ (.Y(_0274_),
    .A(\ctrl[23] ),
    .B(net73));
 sg13g2_nor2b_1 _0865_ (.A(_0273_),
    .B_N(_0274_),
    .Y(_0275_));
 sg13g2_xor2_1 _0866_ (.B(_0275_),
    .A(_0272_),
    .X(_0276_));
 sg13g2_nor2_1 _0867_ (.A(net236),
    .B(net73),
    .Y(_0277_));
 sg13g2_a21oi_1 _0868_ (.A1(net236),
    .A2(_0276_),
    .Y(_0018_),
    .B1(_0277_));
 sg13g2_nand2_1 _0869_ (.Y(_0278_),
    .A(_0269_),
    .B(_0275_));
 sg13g2_a21oi_1 _0870_ (.A1(_0264_),
    .A2(_0266_),
    .Y(_0279_),
    .B1(_0278_));
 sg13g2_o21ai_1 _0871_ (.B1(_0274_),
    .Y(_0280_),
    .A1(_0268_),
    .A2(_0273_));
 sg13g2_nor2_1 _0872_ (.A(_0279_),
    .B(_0280_),
    .Y(_0281_));
 sg13g2_nand2_1 _0873_ (.Y(_0282_),
    .A(net235),
    .B(_0281_));
 sg13g2_nor3_2 _0874_ (.A(net85),
    .B(_0279_),
    .C(_0280_),
    .Y(_0283_));
 sg13g2_a22oi_1 _0875_ (.Y(_0284_),
    .B1(net86),
    .B2(net237),
    .A2(_0282_),
    .A1(net85));
 sg13g2_inv_1 _0876_ (.Y(_0019_),
    .A(_0284_));
 sg13g2_nor2b_1 _0877_ (.A(_0283_),
    .B_N(net240),
    .Y(_0285_));
 sg13g2_xor2_1 _0878_ (.B(_0285_),
    .A(net40),
    .X(_0020_));
 sg13g2_nand3_1 _0879_ (.B(net40),
    .C(net37),
    .A(net240),
    .Y(_0286_));
 sg13g2_nor2_2 _0880_ (.A(_0283_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_a21oi_1 _0881_ (.A1(\nco_phase_acc[17] ),
    .A2(_0285_),
    .Y(_0288_),
    .B1(net37));
 sg13g2_nor2_1 _0882_ (.A(_0287_),
    .B(net38),
    .Y(_0021_));
 sg13g2_xor2_1 _0883_ (.B(_0287_),
    .A(net42),
    .X(_0022_));
 sg13g2_and2_1 _0884_ (.A(net42),
    .B(net27),
    .X(_0289_));
 sg13g2_a21oi_1 _0885_ (.A1(\nco_phase_acc[19] ),
    .A2(_0287_),
    .Y(_0290_),
    .B1(net27));
 sg13g2_a21oi_1 _0886_ (.A1(_0287_),
    .A2(_0289_),
    .Y(_0023_),
    .B1(net28));
 sg13g2_a21oi_1 _0887_ (.A1(_0287_),
    .A2(_0289_),
    .Y(_0291_),
    .B1(net70));
 sg13g2_nand3_1 _0888_ (.B(_0287_),
    .C(_0289_),
    .A(net70),
    .Y(_0292_));
 sg13g2_nor2b_1 _0889_ (.A(_0291_),
    .B_N(_0292_),
    .Y(_0024_));
 sg13g2_nand4_1 _0890_ (.B(net30),
    .C(_0287_),
    .A(net70),
    .Y(_0293_),
    .D(_0289_));
 sg13g2_xnor2_1 _0891_ (.Y(_0025_),
    .A(net30),
    .B(_0292_));
 sg13g2_xnor2_1 _0892_ (.Y(_0026_),
    .A(net26),
    .B(_0293_));
 sg13g2_nor2_1 _0893_ (.A(net241),
    .B(net4),
    .Y(_0294_));
 sg13g2_a21oi_1 _0894_ (.A1(net239),
    .A2(_0157_),
    .Y(_0027_),
    .B1(_0294_));
 sg13g2_nand2_1 _0895_ (.Y(_0295_),
    .A(net205),
    .B(net241));
 sg13g2_o21ai_1 _0896_ (.B1(_0295_),
    .Y(_0028_),
    .A1(net5),
    .A2(net241));
 sg13g2_nor2b_1 _0897_ (.A(\u_lf.ki_sel_latched[0] ),
    .B_N(_0002_),
    .Y(_0296_));
 sg13g2_nand2b_1 _0898_ (.Y(_0297_),
    .B(\u_lf.ki_sel_latched[0] ),
    .A_N(_0002_));
 sg13g2_mux4_1 _0899_ (.S0(\u_lf.ki_sel_latched[0] ),
    .A0(net201),
    .A1(\phase_err_beat[13] ),
    .A2(\phase_err_beat[12] ),
    .A3(net200),
    .S1(_0002_),
    .X(_0298_));
 sg13g2_mux4_1 _0900_ (.S0(\u_lf.ki_sel_latched[0] ),
    .A0(\phase_err_beat[10] ),
    .A1(\phase_err_beat[9] ),
    .A2(net202),
    .A3(\phase_err_beat[11] ),
    .S1(_0002_),
    .X(_0299_));
 sg13g2_nand2_1 _0901_ (.Y(_0300_),
    .A(net183),
    .B(_0299_));
 sg13g2_nand2_1 _0902_ (.Y(_0301_),
    .A(net52),
    .B(_0299_));
 sg13g2_xnor2_1 _0903_ (.Y(_0029_),
    .A(net52),
    .B(_0300_));
 sg13g2_mux4_1 _0904_ (.S0(\u_lf.ki_sel_latched[0] ),
    .A0(net203),
    .A1(\phase_err_beat[10] ),
    .A2(\phase_err_beat[13] ),
    .A3(net202),
    .S1(_0002_),
    .X(_0302_));
 sg13g2_nand2_1 _0905_ (.Y(_0303_),
    .A(\u_lf.i_acc[1] ),
    .B(_0302_));
 sg13g2_xnor2_1 _0906_ (.Y(_0304_),
    .A(net298),
    .B(_0302_));
 sg13g2_o21ai_1 _0907_ (.B1(net183),
    .Y(_0305_),
    .A1(_0301_),
    .A2(_0304_));
 sg13g2_a21oi_1 _0908_ (.A1(_0301_),
    .A2(_0304_),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_a21o_1 _0909_ (.A2(net190),
    .A1(net298),
    .B1(_0306_),
    .X(_0030_));
 sg13g2_nor2_1 _0910_ (.A(net153),
    .B(net183),
    .Y(_0307_));
 sg13g2_o21ai_1 _0911_ (.B1(_0303_),
    .Y(_0308_),
    .A1(_0301_),
    .A2(_0304_));
 sg13g2_mux4_1 _0912_ (.S0(\u_lf.ki_sel_latched[0] ),
    .A0(net202),
    .A1(net203),
    .A2(net201),
    .A3(\phase_err_beat[13] ),
    .S1(_0002_),
    .X(_0309_));
 sg13g2_nand2_1 _0913_ (.Y(_0310_),
    .A(net153),
    .B(_0309_));
 sg13g2_inv_1 _0914_ (.Y(_0311_),
    .A(_0310_));
 sg13g2_or2_1 _0915_ (.X(_0312_),
    .B(_0309_),
    .A(net153));
 sg13g2_nand2_1 _0916_ (.Y(_0313_),
    .A(_0310_),
    .B(_0312_));
 sg13g2_xor2_1 _0917_ (.B(_0313_),
    .A(_0308_),
    .X(_0314_));
 sg13g2_a21oi_1 _0918_ (.A1(net183),
    .A2(_0314_),
    .Y(_0031_),
    .B1(_0307_));
 sg13g2_nor2_1 _0919_ (.A(net278),
    .B(net183),
    .Y(_0315_));
 sg13g2_mux4_1 _0920_ (.S0(\u_lf.ki_sel_latched[0] ),
    .A0(\phase_err_beat[13] ),
    .A1(net202),
    .A2(net200),
    .A3(net201),
    .S1(_0002_),
    .X(_0316_));
 sg13g2_nand2_1 _0921_ (.Y(_0317_),
    .A(net278),
    .B(_0316_));
 sg13g2_xnor2_1 _0922_ (.Y(_0318_),
    .A(net278),
    .B(_0316_));
 sg13g2_a21oi_1 _0923_ (.A1(_0308_),
    .A2(_0312_),
    .Y(_0319_),
    .B1(_0311_));
 sg13g2_xnor2_1 _0924_ (.Y(_0320_),
    .A(_0318_),
    .B(_0319_));
 sg13g2_a21oi_1 _0925_ (.A1(net183),
    .A2(_0320_),
    .Y(_0032_),
    .B1(_0315_));
 sg13g2_nor2_1 _0926_ (.A(net282),
    .B(net183),
    .Y(_0321_));
 sg13g2_o21ai_1 _0927_ (.B1(_0317_),
    .Y(_0322_),
    .A1(_0318_),
    .A2(_0319_));
 sg13g2_nor2_1 _0928_ (.A(_0296_),
    .B(_0298_),
    .Y(_0323_));
 sg13g2_a21oi_1 _0929_ (.A1(_0156_),
    .A2(_0296_),
    .Y(_0324_),
    .B1(_0323_));
 sg13g2_and2_1 _0930_ (.A(net282),
    .B(_0324_),
    .X(_0325_));
 sg13g2_xnor2_1 _0931_ (.Y(_0326_),
    .A(net282),
    .B(_0324_));
 sg13g2_inv_1 _0932_ (.Y(_0327_),
    .A(_0326_));
 sg13g2_xnor2_1 _0933_ (.Y(_0328_),
    .A(_0322_),
    .B(_0327_));
 sg13g2_a21oi_1 _0934_ (.A1(net183),
    .A2(_0328_),
    .Y(_0033_),
    .B1(_0321_));
 sg13g2_nor2_1 _0935_ (.A(net306),
    .B(uo_out[0]),
    .Y(_0329_));
 sg13g2_a21oi_1 _0936_ (.A1(_0322_),
    .A2(_0327_),
    .Y(_0330_),
    .B1(_0325_));
 sg13g2_nor2_1 _0937_ (.A(net201),
    .B(_0297_),
    .Y(_0331_));
 sg13g2_a21oi_1 _0938_ (.A1(_0156_),
    .A2(_0297_),
    .Y(_0332_),
    .B1(_0331_));
 sg13g2_nor2_1 _0939_ (.A(\u_lf.i_acc[5] ),
    .B(_0332_),
    .Y(_0333_));
 sg13g2_xnor2_1 _0940_ (.Y(_0334_),
    .A(net306),
    .B(_0332_));
 sg13g2_xnor2_1 _0941_ (.Y(_0335_),
    .A(_0330_),
    .B(_0334_));
 sg13g2_a21oi_1 _0942_ (.A1(uo_out[0]),
    .A2(_0335_),
    .Y(_0034_),
    .B1(_0329_));
 sg13g2_xnor2_1 _0943_ (.Y(_0336_),
    .A(net200),
    .B(net275));
 sg13g2_a221oi_1 _0944_ (.B2(\u_lf.i_acc[5] ),
    .C1(_0325_),
    .B1(_0332_),
    .A1(_0322_),
    .Y(_0337_),
    .A2(_0327_));
 sg13g2_nor3_1 _0945_ (.A(_0333_),
    .B(_0336_),
    .C(_0337_),
    .Y(_0338_));
 sg13g2_o21ai_1 _0946_ (.B1(_0336_),
    .Y(_0339_),
    .A1(_0333_),
    .A2(_0337_));
 sg13g2_nand2_1 _0947_ (.Y(_0340_),
    .A(net275),
    .B(net190));
 sg13g2_nand2_1 _0948_ (.Y(_0341_),
    .A(net185),
    .B(_0339_));
 sg13g2_o21ai_1 _0949_ (.B1(_0340_),
    .Y(_0035_),
    .A1(_0338_),
    .A2(_0341_));
 sg13g2_xor2_1 _0950_ (.B(net248),
    .A(net199),
    .X(_0342_));
 sg13g2_a21oi_1 _0951_ (.A1(net199),
    .A2(\u_lf.i_acc[6] ),
    .Y(_0343_),
    .B1(_0338_));
 sg13g2_xor2_1 _0952_ (.B(_0343_),
    .A(_0342_),
    .X(_0344_));
 sg13g2_nand2_1 _0953_ (.Y(_0345_),
    .A(net248),
    .B(net190));
 sg13g2_o21ai_1 _0954_ (.B1(_0345_),
    .Y(_0036_),
    .A1(net189),
    .A2(_0344_));
 sg13g2_o21ai_1 _0955_ (.B1(net199),
    .Y(_0346_),
    .A1(\u_lf.i_acc[7] ),
    .A2(\u_lf.i_acc[6] ));
 sg13g2_inv_1 _0956_ (.Y(_0347_),
    .A(_0346_));
 sg13g2_a21o_2 _0957_ (.A2(_0342_),
    .A1(_0338_),
    .B1(_0347_),
    .X(_0348_));
 sg13g2_xor2_1 _0958_ (.B(net279),
    .A(net198),
    .X(_0349_));
 sg13g2_and2_1 _0959_ (.A(_0348_),
    .B(_0349_),
    .X(_0350_));
 sg13g2_nand2_1 _0960_ (.Y(_0351_),
    .A(net279),
    .B(net189));
 sg13g2_o21ai_1 _0961_ (.B1(net181),
    .Y(_0352_),
    .A1(_0348_),
    .A2(_0349_));
 sg13g2_o21ai_1 _0962_ (.B1(_0351_),
    .Y(_0037_),
    .A1(_0350_),
    .A2(_0352_));
 sg13g2_nor2_1 _0963_ (.A(net312),
    .B(net185),
    .Y(_0353_));
 sg13g2_xor2_1 _0964_ (.B(net312),
    .A(net198),
    .X(_0354_));
 sg13g2_a21oi_1 _0965_ (.A1(net198),
    .A2(net279),
    .Y(_0355_),
    .B1(_0350_));
 sg13g2_xor2_1 _0966_ (.B(_0355_),
    .A(_0354_),
    .X(_0356_));
 sg13g2_a21oi_1 _0967_ (.A1(net185),
    .A2(_0356_),
    .Y(_0038_),
    .B1(_0353_));
 sg13g2_xnor2_1 _0968_ (.Y(_0357_),
    .A(net198),
    .B(net263));
 sg13g2_o21ai_1 _0969_ (.B1(net198),
    .Y(_0358_),
    .A1(\u_lf.i_acc[9] ),
    .A2(\u_lf.i_acc[8] ));
 sg13g2_nand2_1 _0970_ (.Y(_0359_),
    .A(_0350_),
    .B(_0354_));
 sg13g2_a21oi_1 _0971_ (.A1(_0358_),
    .A2(_0359_),
    .Y(_0360_),
    .B1(_0357_));
 sg13g2_nand3_1 _0972_ (.B(_0358_),
    .C(_0359_),
    .A(_0357_),
    .Y(_0361_));
 sg13g2_nand2_1 _0973_ (.Y(_0362_),
    .A(net263),
    .B(net189));
 sg13g2_nand2_1 _0974_ (.Y(_0363_),
    .A(net181),
    .B(_0361_));
 sg13g2_o21ai_1 _0975_ (.B1(net264),
    .Y(_0039_),
    .A1(_0360_),
    .A2(_0363_));
 sg13g2_nor2_1 _0976_ (.A(net305),
    .B(net185),
    .Y(_0364_));
 sg13g2_xnor2_1 _0977_ (.Y(_0365_),
    .A(net198),
    .B(net305));
 sg13g2_a21oi_1 _0978_ (.A1(net198),
    .A2(net263),
    .Y(_0366_),
    .B1(_0360_));
 sg13g2_xnor2_1 _0979_ (.Y(_0367_),
    .A(_0365_),
    .B(_0366_));
 sg13g2_a21oi_1 _0980_ (.A1(net185),
    .A2(_0367_),
    .Y(_0040_),
    .B1(_0364_));
 sg13g2_xor2_1 _0981_ (.B(\u_lf.i_acc[12] ),
    .A(net196),
    .X(_0368_));
 sg13g2_inv_1 _0982_ (.Y(_0369_),
    .A(_0368_));
 sg13g2_o21ai_1 _0983_ (.B1(net198),
    .Y(_0370_),
    .A1(\u_lf.i_acc[11] ),
    .A2(\u_lf.i_acc[10] ));
 sg13g2_and2_1 _0984_ (.A(_0358_),
    .B(_0370_),
    .X(_0371_));
 sg13g2_nor2_1 _0985_ (.A(_0357_),
    .B(_0365_),
    .Y(_0372_));
 sg13g2_nand3_1 _0986_ (.B(_0354_),
    .C(_0372_),
    .A(_0349_),
    .Y(_0373_));
 sg13g2_nand2b_1 _0987_ (.Y(_0374_),
    .B(_0348_),
    .A_N(_0373_));
 sg13g2_a21oi_1 _0988_ (.A1(_0371_),
    .A2(_0374_),
    .Y(_0375_),
    .B1(_0369_));
 sg13g2_inv_1 _0989_ (.Y(_0376_),
    .A(_0375_));
 sg13g2_nand3_1 _0990_ (.B(_0371_),
    .C(_0374_),
    .A(_0369_),
    .Y(_0377_));
 sg13g2_nand3_1 _0991_ (.B(_0376_),
    .C(_0377_),
    .A(net181),
    .Y(_0378_));
 sg13g2_o21ai_1 _0992_ (.B1(_0378_),
    .Y(_0041_),
    .A1(_0158_),
    .A2(net182));
 sg13g2_nor2_1 _0993_ (.A(net243),
    .B(net181),
    .Y(_0379_));
 sg13g2_xnor2_1 _0994_ (.Y(_0380_),
    .A(net196),
    .B(\u_lf.i_acc[13] ));
 sg13g2_a21oi_1 _0995_ (.A1(net196),
    .A2(\u_lf.i_acc[12] ),
    .Y(_0381_),
    .B1(_0375_));
 sg13g2_xnor2_1 _0996_ (.Y(_0382_),
    .A(_0380_),
    .B(_0381_));
 sg13g2_a21oi_1 _0997_ (.A1(net181),
    .A2(_0382_),
    .Y(_0042_),
    .B1(_0379_));
 sg13g2_o21ai_1 _0998_ (.B1(net196),
    .Y(_0383_),
    .A1(\u_lf.i_acc[13] ),
    .A2(\u_lf.i_acc[12] ));
 sg13g2_o21ai_1 _0999_ (.B1(_0383_),
    .Y(_0384_),
    .A1(_0376_),
    .A2(_0380_));
 sg13g2_and2_1 _1000_ (.A(net197),
    .B(\u_lf.i_acc[14] ),
    .X(_0385_));
 sg13g2_xor2_1 _1001_ (.B(\u_lf.i_acc[14] ),
    .A(net196),
    .X(_0386_));
 sg13g2_inv_1 _1002_ (.Y(_0387_),
    .A(_0386_));
 sg13g2_o21ai_1 _1003_ (.B1(net181),
    .Y(_0388_),
    .A1(_0384_),
    .A2(_0386_));
 sg13g2_a21oi_1 _1004_ (.A1(_0384_),
    .A2(_0386_),
    .Y(_0389_),
    .B1(_0388_));
 sg13g2_a21o_1 _1005_ (.A2(net188),
    .A1(net272),
    .B1(_0389_),
    .X(_0043_));
 sg13g2_nor2_1 _1006_ (.A(net266),
    .B(net181),
    .Y(_0390_));
 sg13g2_xnor2_1 _1007_ (.Y(_0391_),
    .A(net196),
    .B(net266));
 sg13g2_a21oi_1 _1008_ (.A1(_0384_),
    .A2(_0386_),
    .Y(_0392_),
    .B1(_0385_));
 sg13g2_xnor2_1 _1009_ (.Y(_0393_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_a21oi_1 _1010_ (.A1(net181),
    .A2(_0393_),
    .Y(_0044_),
    .B1(_0390_));
 sg13g2_nand2_1 _1011_ (.Y(_0394_),
    .A(net125),
    .B(net187));
 sg13g2_xor2_1 _1012_ (.B(net338),
    .A(net195),
    .X(_0395_));
 sg13g2_or4_1 _1013_ (.A(_0369_),
    .B(_0380_),
    .C(_0387_),
    .D(_0391_),
    .X(_0396_));
 sg13g2_nor2_1 _1014_ (.A(_0373_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_o21ai_1 _1015_ (.B1(net196),
    .Y(_0398_),
    .A1(\u_lf.i_acc[15] ),
    .A2(\u_lf.i_acc[14] ));
 sg13g2_and2_1 _1016_ (.A(_0383_),
    .B(_0398_),
    .X(_0399_));
 sg13g2_nand2_1 _1017_ (.Y(_0400_),
    .A(_0371_),
    .B(_0399_));
 sg13g2_a21oi_2 _1018_ (.B1(_0400_),
    .Y(_0401_),
    .A2(_0397_),
    .A1(_0348_));
 sg13g2_nor2b_1 _1019_ (.A(_0401_),
    .B_N(_0395_),
    .Y(_0402_));
 sg13g2_xor2_1 _1020_ (.B(_0401_),
    .A(_0395_),
    .X(_0403_));
 sg13g2_o21ai_1 _1021_ (.B1(_0394_),
    .Y(_0045_),
    .A1(net187),
    .A2(_0403_));
 sg13g2_nor2_1 _1022_ (.A(net160),
    .B(net179),
    .Y(_0404_));
 sg13g2_xor2_1 _1023_ (.B(\u_lf.i_acc[17] ),
    .A(net195),
    .X(_0405_));
 sg13g2_a21oi_1 _1024_ (.A1(net195),
    .A2(net125),
    .Y(_0406_),
    .B1(_0402_));
 sg13g2_xor2_1 _1025_ (.B(_0406_),
    .A(_0405_),
    .X(_0407_));
 sg13g2_a21oi_1 _1026_ (.A1(net179),
    .A2(_0407_),
    .Y(_0046_),
    .B1(_0404_));
 sg13g2_o21ai_1 _1027_ (.B1(net195),
    .Y(_0408_),
    .A1(\u_lf.i_acc[17] ),
    .A2(net337));
 sg13g2_inv_1 _1028_ (.Y(_0409_),
    .A(_0408_));
 sg13g2_nand2_1 _1029_ (.Y(_0410_),
    .A(_0402_),
    .B(_0405_));
 sg13g2_nand2_1 _1030_ (.Y(_0411_),
    .A(net194),
    .B(\u_lf.i_acc[18] ));
 sg13g2_xnor2_1 _1031_ (.Y(_0412_),
    .A(net194),
    .B(\u_lf.i_acc[18] ));
 sg13g2_a21oi_1 _1032_ (.A1(_0408_),
    .A2(_0410_),
    .Y(_0413_),
    .B1(_0412_));
 sg13g2_nand3_1 _1033_ (.B(_0410_),
    .C(_0412_),
    .A(_0408_),
    .Y(_0414_));
 sg13g2_nand2_1 _1034_ (.Y(_0415_),
    .A(net112),
    .B(net187));
 sg13g2_nand2_1 _1035_ (.Y(_0416_),
    .A(net179),
    .B(_0414_));
 sg13g2_o21ai_1 _1036_ (.B1(_0415_),
    .Y(_0047_),
    .A1(_0413_),
    .A2(_0416_));
 sg13g2_nor2_1 _1037_ (.A(net140),
    .B(net179),
    .Y(_0417_));
 sg13g2_xnor2_1 _1038_ (.Y(_0418_),
    .A(net194),
    .B(net140));
 sg13g2_a21oi_1 _1039_ (.A1(net195),
    .A2(net112),
    .Y(_0419_),
    .B1(_0413_));
 sg13g2_xnor2_1 _1040_ (.Y(_0420_),
    .A(_0418_),
    .B(_0419_));
 sg13g2_a21oi_1 _1041_ (.A1(net179),
    .A2(_0420_),
    .Y(_0048_),
    .B1(_0417_));
 sg13g2_o21ai_1 _1042_ (.B1(net194),
    .Y(_0421_),
    .A1(\u_lf.i_acc[19] ),
    .A2(\u_lf.i_acc[18] ));
 sg13g2_and2_1 _1043_ (.A(_0408_),
    .B(_0421_),
    .X(_0422_));
 sg13g2_nand2_1 _1044_ (.Y(_0423_),
    .A(_0408_),
    .B(_0421_));
 sg13g2_nor2_1 _1045_ (.A(_0412_),
    .B(_0418_),
    .Y(_0424_));
 sg13g2_nand3_1 _1046_ (.B(_0405_),
    .C(_0424_),
    .A(_0395_),
    .Y(_0425_));
 sg13g2_inv_1 _1047_ (.Y(_0426_),
    .A(_0425_));
 sg13g2_o21ai_1 _1048_ (.B1(_0422_),
    .Y(_0427_),
    .A1(_0401_),
    .A2(_0425_));
 sg13g2_and2_1 _1049_ (.A(net194),
    .B(\u_lf.i_acc[20] ),
    .X(_0428_));
 sg13g2_xor2_1 _1050_ (.B(\u_lf.i_acc[20] ),
    .A(net194),
    .X(_0429_));
 sg13g2_o21ai_1 _1051_ (.B1(net179),
    .Y(_0430_),
    .A1(_0427_),
    .A2(_0429_));
 sg13g2_a21oi_1 _1052_ (.A1(_0427_),
    .A2(_0429_),
    .Y(_0431_),
    .B1(_0430_));
 sg13g2_a21o_1 _1053_ (.A2(net187),
    .A1(net256),
    .B1(_0431_),
    .X(_0049_));
 sg13g2_nor2_1 _1054_ (.A(net141),
    .B(net179),
    .Y(_0432_));
 sg13g2_xor2_1 _1055_ (.B(net141),
    .A(net194),
    .X(_0433_));
 sg13g2_a21oi_1 _1056_ (.A1(_0427_),
    .A2(_0429_),
    .Y(_0434_),
    .B1(_0428_));
 sg13g2_xor2_1 _1057_ (.B(_0434_),
    .A(_0433_),
    .X(_0435_));
 sg13g2_a21oi_1 _1058_ (.A1(net179),
    .A2(_0435_),
    .Y(_0050_),
    .B1(_0432_));
 sg13g2_nor2_1 _1059_ (.A(net296),
    .B(net177),
    .Y(_0436_));
 sg13g2_o21ai_1 _1060_ (.B1(net194),
    .Y(_0437_),
    .A1(\u_lf.i_acc[21] ),
    .A2(\u_lf.i_acc[20] ));
 sg13g2_nand2_1 _1061_ (.Y(_0438_),
    .A(_0429_),
    .B(_0433_));
 sg13g2_nor2b_1 _1062_ (.A(_0438_),
    .B_N(_0427_),
    .Y(_0439_));
 sg13g2_nor2b_1 _1063_ (.A(_0439_),
    .B_N(_0437_),
    .Y(_0440_));
 sg13g2_and2_1 _1064_ (.A(net192),
    .B(\u_lf.i_acc[22] ),
    .X(_0441_));
 sg13g2_nand2_1 _1065_ (.Y(_0442_),
    .A(net192),
    .B(net296));
 sg13g2_or2_1 _1066_ (.X(_0443_),
    .B(\u_lf.i_acc[22] ),
    .A(net192));
 sg13g2_nand2_2 _1067_ (.Y(_0444_),
    .A(_0442_),
    .B(_0443_));
 sg13g2_xnor2_1 _1068_ (.Y(_0445_),
    .A(_0440_),
    .B(_0444_));
 sg13g2_a21oi_1 _1069_ (.A1(net177),
    .A2(_0445_),
    .Y(_0051_),
    .B1(_0436_));
 sg13g2_nor2_1 _1070_ (.A(net157),
    .B(net177),
    .Y(_0446_));
 sg13g2_xnor2_1 _1071_ (.Y(_0447_),
    .A(net192),
    .B(net157));
 sg13g2_o21ai_1 _1072_ (.B1(_0442_),
    .Y(_0448_),
    .A1(_0440_),
    .A2(_0444_));
 sg13g2_xor2_1 _1073_ (.B(_0448_),
    .A(_0447_),
    .X(_0449_));
 sg13g2_a21oi_1 _1074_ (.A1(net177),
    .A2(_0449_),
    .Y(_0052_),
    .B1(_0446_));
 sg13g2_nor2_1 _1075_ (.A(net273),
    .B(net177),
    .Y(_0450_));
 sg13g2_o21ai_1 _1076_ (.B1(net193),
    .Y(_0451_),
    .A1(\u_lf.i_acc[23] ),
    .A2(\u_lf.i_acc[22] ));
 sg13g2_nand3_1 _1077_ (.B(_0437_),
    .C(_0451_),
    .A(_0422_),
    .Y(_0452_));
 sg13g2_inv_1 _1078_ (.Y(_0453_),
    .A(_0452_));
 sg13g2_nor4_1 _1079_ (.A(_0425_),
    .B(_0438_),
    .C(_0444_),
    .D(_0447_),
    .Y(_0454_));
 sg13g2_inv_1 _1080_ (.Y(_0455_),
    .A(_0454_));
 sg13g2_o21ai_1 _1081_ (.B1(_0453_),
    .Y(_0456_),
    .A1(_0401_),
    .A2(_0455_));
 sg13g2_nand2_1 _1082_ (.Y(_0457_),
    .A(net192),
    .B(\u_lf.i_acc[24] ));
 sg13g2_xnor2_1 _1083_ (.Y(_0458_),
    .A(net192),
    .B(\u_lf.i_acc[24] ));
 sg13g2_nand2b_1 _1084_ (.Y(_0459_),
    .B(_0456_),
    .A_N(_0458_));
 sg13g2_xor2_1 _1085_ (.B(_0458_),
    .A(_0456_),
    .X(_0460_));
 sg13g2_a21oi_1 _1086_ (.A1(net177),
    .A2(_0460_),
    .Y(_0053_),
    .B1(_0450_));
 sg13g2_nor2_1 _1087_ (.A(net147),
    .B(net177),
    .Y(_0461_));
 sg13g2_xor2_1 _1088_ (.B(net147),
    .A(net192),
    .X(_0462_));
 sg13g2_nand2_1 _1089_ (.Y(_0463_),
    .A(_0457_),
    .B(_0459_));
 sg13g2_xnor2_1 _1090_ (.Y(_0464_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_a21oi_1 _1091_ (.A1(net177),
    .A2(_0464_),
    .Y(_0054_),
    .B1(_0461_));
 sg13g2_nor2_1 _1092_ (.A(net270),
    .B(net178),
    .Y(_0465_));
 sg13g2_o21ai_1 _1093_ (.B1(net192),
    .Y(_0466_),
    .A1(\u_lf.i_acc[25] ),
    .A2(\u_lf.i_acc[24] ));
 sg13g2_inv_1 _1094_ (.Y(_0467_),
    .A(_0466_));
 sg13g2_nor2b_1 _1095_ (.A(_0458_),
    .B_N(_0462_),
    .Y(_0468_));
 sg13g2_nand2b_1 _1096_ (.Y(_0469_),
    .B(_0462_),
    .A_N(_0458_));
 sg13g2_a21oi_1 _1097_ (.A1(_0456_),
    .A2(_0468_),
    .Y(_0470_),
    .B1(_0467_));
 sg13g2_and2_1 _1098_ (.A(net193),
    .B(\u_lf.i_acc[26] ),
    .X(_0471_));
 sg13g2_xor2_1 _1099_ (.B(\u_lf.i_acc[26] ),
    .A(net197),
    .X(_0472_));
 sg13g2_xnor2_1 _1100_ (.Y(_0473_),
    .A(net193),
    .B(net270));
 sg13g2_nor2_1 _1101_ (.A(_0470_),
    .B(_0473_),
    .Y(_0474_));
 sg13g2_xnor2_1 _1102_ (.Y(_0475_),
    .A(_0470_),
    .B(_0473_));
 sg13g2_a21oi_1 _1103_ (.A1(net178),
    .A2(_0475_),
    .Y(_0055_),
    .B1(_0465_));
 sg13g2_nor2_1 _1104_ (.A(net253),
    .B(net178),
    .Y(_0476_));
 sg13g2_xnor2_1 _1105_ (.Y(_0477_),
    .A(net193),
    .B(net253));
 sg13g2_nor2_1 _1106_ (.A(_0471_),
    .B(_0474_),
    .Y(_0478_));
 sg13g2_xnor2_1 _1107_ (.Y(_0479_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_a21oi_1 _1108_ (.A1(net178),
    .A2(_0479_),
    .Y(_0056_),
    .B1(_0476_));
 sg13g2_nor2_1 _1109_ (.A(net146),
    .B(net178),
    .Y(_0480_));
 sg13g2_nand2_1 _1110_ (.Y(_0481_),
    .A(net193),
    .B(\u_lf.i_acc[28] ));
 sg13g2_xnor2_1 _1111_ (.Y(_0482_),
    .A(net193),
    .B(net146));
 sg13g2_o21ai_1 _1112_ (.B1(net193),
    .Y(_0483_),
    .A1(net335),
    .A2(\u_lf.i_acc[26] ));
 sg13g2_nand2_1 _1113_ (.Y(_0484_),
    .A(_0466_),
    .B(net336));
 sg13g2_nor3_1 _1114_ (.A(_0469_),
    .B(_0473_),
    .C(_0477_),
    .Y(_0485_));
 sg13g2_a21oi_1 _1115_ (.A1(_0456_),
    .A2(_0485_),
    .Y(_0486_),
    .B1(_0484_));
 sg13g2_xnor2_1 _1116_ (.Y(_0487_),
    .A(_0482_),
    .B(_0486_));
 sg13g2_a21oi_1 _1117_ (.A1(net178),
    .A2(_0487_),
    .Y(_0057_),
    .B1(_0480_));
 sg13g2_nor2_1 _1118_ (.A(net106),
    .B(net182),
    .Y(_0488_));
 sg13g2_o21ai_1 _1119_ (.B1(_0481_),
    .Y(_0489_),
    .A1(_0482_),
    .A2(_0486_));
 sg13g2_xor2_1 _1120_ (.B(net196),
    .A(net106),
    .X(_0490_));
 sg13g2_xnor2_1 _1121_ (.Y(_0491_),
    .A(_0489_),
    .B(_0490_));
 sg13g2_a21oi_1 _1122_ (.A1(net178),
    .A2(_0491_),
    .Y(_0058_),
    .B1(_0488_));
 sg13g2_nor2b_1 _1123_ (.A(net205),
    .B_N(net207),
    .Y(_0492_));
 sg13g2_nor2b_1 _1124_ (.A(net207),
    .B_N(net205),
    .Y(_0493_));
 sg13g2_mux4_1 _1125_ (.S0(net206),
    .A0(\phase_err_beat[5] ),
    .A1(\phase_err_beat[4] ),
    .A2(\phase_err_beat[7] ),
    .A3(\phase_err_beat[6] ),
    .S1(net204),
    .X(_0494_));
 sg13g2_mux4_1 _1126_ (.S0(net206),
    .A0(\phase_err_beat[4] ),
    .A1(\phase_err_beat[3] ),
    .A2(\phase_err_beat[6] ),
    .A3(\phase_err_beat[5] ),
    .S1(net204),
    .X(_0495_));
 sg13g2_a22oi_1 _1127_ (.Y(_0496_),
    .B1(_0495_),
    .B2(\u_lf.i_acc[0] ),
    .A2(_0494_),
    .A1(\u_lf.i_acc[1] ));
 sg13g2_mux4_1 _1128_ (.S0(net206),
    .A0(\phase_err_beat[6] ),
    .A1(\phase_err_beat[5] ),
    .A2(\phase_err_beat[8] ),
    .A3(\phase_err_beat[7] ),
    .S1(net204),
    .X(_0497_));
 sg13g2_nor2_1 _1129_ (.A(\u_lf.i_acc[2] ),
    .B(_0497_),
    .Y(_0498_));
 sg13g2_nor2_1 _1130_ (.A(\u_lf.i_acc[1] ),
    .B(_0494_),
    .Y(_0499_));
 sg13g2_nor3_1 _1131_ (.A(_0496_),
    .B(_0498_),
    .C(_0499_),
    .Y(_0500_));
 sg13g2_mux4_1 _1132_ (.S0(net206),
    .A0(\phase_err_beat[7] ),
    .A1(\phase_err_beat[6] ),
    .A2(\phase_err_beat[9] ),
    .A3(\phase_err_beat[8] ),
    .S1(net204),
    .X(_0501_));
 sg13g2_a221oi_1 _1133_ (.B2(\u_lf.i_acc[3] ),
    .C1(_0500_),
    .B1(_0501_),
    .A1(\u_lf.i_acc[2] ),
    .Y(_0502_),
    .A2(_0497_));
 sg13g2_mux4_1 _1134_ (.S0(net207),
    .A0(net203),
    .A1(\phase_err_beat[10] ),
    .A2(\phase_err_beat[13] ),
    .A3(\phase_err_beat[12] ),
    .S1(net204),
    .X(_0503_));
 sg13g2_nand2_1 _1135_ (.Y(_0504_),
    .A(\u_lf.i_acc[7] ),
    .B(_0503_));
 sg13g2_or2_1 _1136_ (.X(_0505_),
    .B(_0503_),
    .A(\u_lf.i_acc[7] ));
 sg13g2_mux2_1 _1137_ (.A0(net202),
    .A1(\phase_err_beat[13] ),
    .S(net207),
    .X(_0506_));
 sg13g2_mux4_1 _1138_ (.S0(net206),
    .A0(\phase_err_beat[10] ),
    .A1(\phase_err_beat[9] ),
    .A2(net202),
    .A3(net203),
    .S1(net204),
    .X(_0507_));
 sg13g2_xor2_1 _1139_ (.B(_0507_),
    .A(\u_lf.i_acc[6] ),
    .X(_0508_));
 sg13g2_and3_1 _1140_ (.X(_0509_),
    .A(_0504_),
    .B(_0505_),
    .C(_0508_));
 sg13g2_mux4_1 _1141_ (.S0(net206),
    .A0(\phase_err_beat[9] ),
    .A1(\phase_err_beat[8] ),
    .A2(net203),
    .A3(\phase_err_beat[10] ),
    .S1(net205),
    .X(_0510_));
 sg13g2_nor2_1 _1142_ (.A(\u_lf.i_acc[5] ),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_nand2_1 _1143_ (.Y(_0512_),
    .A(\u_lf.i_acc[5] ),
    .B(_0510_));
 sg13g2_mux4_1 _1144_ (.S0(net206),
    .A0(\phase_err_beat[8] ),
    .A1(\phase_err_beat[7] ),
    .A2(\phase_err_beat[10] ),
    .A3(\phase_err_beat[9] ),
    .S1(net204),
    .X(_0513_));
 sg13g2_nand2_1 _1145_ (.Y(_0514_),
    .A(\u_lf.i_acc[4] ),
    .B(_0513_));
 sg13g2_nor2_1 _1146_ (.A(\u_lf.i_acc[3] ),
    .B(_0501_),
    .Y(_0515_));
 sg13g2_xor2_1 _1147_ (.B(_0513_),
    .A(\u_lf.i_acc[4] ),
    .X(_0516_));
 sg13g2_nor2_1 _1148_ (.A(_0511_),
    .B(_0515_),
    .Y(_0517_));
 sg13g2_nand4_1 _1149_ (.B(_0512_),
    .C(_0516_),
    .A(_0509_),
    .Y(_0518_),
    .D(_0517_));
 sg13g2_o21ai_1 _1150_ (.B1(_0512_),
    .Y(_0519_),
    .A1(_0511_),
    .A2(_0514_));
 sg13g2_and3_1 _1151_ (.X(_0520_),
    .A(\u_lf.i_acc[6] ),
    .B(_0505_),
    .C(_0507_));
 sg13g2_a221oi_1 _1152_ (.B2(_0519_),
    .C1(_0520_),
    .B1(_0509_),
    .A1(\u_lf.i_acc[7] ),
    .Y(_0521_),
    .A2(_0503_));
 sg13g2_o21ai_1 _1153_ (.B1(_0521_),
    .Y(_0522_),
    .A1(_0502_),
    .A2(_0518_));
 sg13g2_nor3_1 _1154_ (.A(net205),
    .B(_0157_),
    .C(net203),
    .Y(_0523_));
 sg13g2_nor3_1 _1155_ (.A(_0492_),
    .B(_0493_),
    .C(_0506_),
    .Y(_0524_));
 sg13g2_nor2b_1 _1156_ (.A(net201),
    .B_N(_0493_),
    .Y(_0525_));
 sg13g2_nor2b_1 _1157_ (.A(net207),
    .B_N(net201),
    .Y(_0526_));
 sg13g2_nor3_1 _1158_ (.A(_0523_),
    .B(_0524_),
    .C(_0525_),
    .Y(_0527_));
 sg13g2_nand2_1 _1159_ (.Y(_0528_),
    .A(\u_lf.i_acc[8] ),
    .B(_0527_));
 sg13g2_xnor2_1 _1160_ (.Y(_0529_),
    .A(\u_lf.i_acc[8] ),
    .B(_0527_));
 sg13g2_nand2b_1 _1161_ (.Y(_0530_),
    .B(_0522_),
    .A_N(_0529_));
 sg13g2_and2_1 _1162_ (.A(net204),
    .B(net199),
    .X(_0531_));
 sg13g2_mux4_1 _1163_ (.S0(net207),
    .A0(\phase_err_beat[13] ),
    .A1(net202),
    .A2(net199),
    .A3(net201),
    .S1(_0001_),
    .X(_0532_));
 sg13g2_nand2_1 _1164_ (.Y(_0533_),
    .A(\u_lf.i_acc[9] ),
    .B(_0532_));
 sg13g2_a221oi_1 _1165_ (.B2(_0153_),
    .C1(_0531_),
    .B1(_0526_),
    .A1(_0492_),
    .Y(_0534_),
    .A2(_0506_));
 sg13g2_nand2b_1 _1166_ (.Y(_0535_),
    .B(\u_lf.i_acc[10] ),
    .A_N(_0534_));
 sg13g2_xnor2_1 _1167_ (.Y(_0536_),
    .A(\u_lf.i_acc[10] ),
    .B(_0534_));
 sg13g2_nand3b_1 _1168_ (.B(net207),
    .C(\phase_err_beat[14] ),
    .Y(_0537_),
    .A_N(net205));
 sg13g2_o21ai_1 _1169_ (.B1(_0537_),
    .Y(_0538_),
    .A1(_0156_),
    .A2(_0492_));
 sg13g2_nand2_1 _1170_ (.Y(_0539_),
    .A(\u_lf.i_acc[11] ),
    .B(_0538_));
 sg13g2_nor2_1 _1171_ (.A(\u_lf.i_acc[11] ),
    .B(_0538_),
    .Y(_0540_));
 sg13g2_xor2_1 _1172_ (.B(_0538_),
    .A(\u_lf.i_acc[11] ),
    .X(_0541_));
 sg13g2_nor2_1 _1173_ (.A(\u_lf.i_acc[9] ),
    .B(_0532_),
    .Y(_0542_));
 sg13g2_nand2_1 _1174_ (.Y(_0543_),
    .A(_0536_),
    .B(_0541_));
 sg13g2_nor2_1 _1175_ (.A(_0542_),
    .B(_0543_),
    .Y(_0544_));
 sg13g2_xnor2_1 _1176_ (.Y(_0545_),
    .A(\u_lf.i_acc[9] ),
    .B(_0532_));
 sg13g2_nor3_1 _1177_ (.A(_0529_),
    .B(_0543_),
    .C(_0545_),
    .Y(_0546_));
 sg13g2_nand2_1 _1178_ (.Y(_0547_),
    .A(_0528_),
    .B(_0533_));
 sg13g2_o21ai_1 _1179_ (.B1(_0539_),
    .Y(_0548_),
    .A1(_0535_),
    .A2(_0540_));
 sg13g2_a221oi_1 _1180_ (.B2(_0544_),
    .C1(_0548_),
    .B1(_0547_),
    .A1(_0522_),
    .Y(_0549_),
    .A2(_0546_));
 sg13g2_o21ai_1 _1181_ (.B1(_0399_),
    .Y(_0550_),
    .A1(_0396_),
    .A2(_0549_));
 sg13g2_a21oi_2 _1182_ (.B1(_0452_),
    .Y(_0551_),
    .A2(_0550_),
    .A1(_0454_));
 sg13g2_a21o_1 _1183_ (.A2(_0550_),
    .A1(_0454_),
    .B1(_0452_),
    .X(_0552_));
 sg13g2_o21ai_1 _1184_ (.B1(_0466_),
    .Y(_0553_),
    .A1(_0469_),
    .A2(_0551_));
 sg13g2_a21oi_1 _1185_ (.A1(_0472_),
    .A2(_0553_),
    .Y(_0554_),
    .B1(_0471_));
 sg13g2_xor2_1 _1186_ (.B(_0554_),
    .A(_0477_),
    .X(_0555_));
 sg13g2_a21oi_1 _1187_ (.A1(_0426_),
    .A2(_0550_),
    .Y(_0556_),
    .B1(_0423_));
 sg13g2_o21ai_1 _1188_ (.B1(_0437_),
    .Y(_0557_),
    .A1(_0438_),
    .A2(_0556_));
 sg13g2_a21oi_1 _1189_ (.A1(_0443_),
    .A2(_0557_),
    .Y(_0558_),
    .B1(_0441_));
 sg13g2_xor2_1 _1190_ (.B(_0558_),
    .A(_0447_),
    .X(_0559_));
 sg13g2_xnor2_1 _1191_ (.Y(_0560_),
    .A(_0472_),
    .B(_0553_));
 sg13g2_xnor2_1 _1192_ (.Y(_0561_),
    .A(_0458_),
    .B(_0551_));
 sg13g2_o21ai_1 _1193_ (.B1(_0457_),
    .Y(_0562_),
    .A1(_0458_),
    .A2(_0551_));
 sg13g2_xnor2_1 _1194_ (.Y(_0563_),
    .A(_0462_),
    .B(_0562_));
 sg13g2_a21oi_1 _1195_ (.A1(_0485_),
    .A2(_0552_),
    .Y(_0564_),
    .B1(_0484_));
 sg13g2_xnor2_1 _1196_ (.Y(_0565_),
    .A(_0482_),
    .B(_0564_));
 sg13g2_nor4_1 _1197_ (.A(_0560_),
    .B(_0561_),
    .C(_0563_),
    .D(_0565_),
    .Y(_0566_));
 sg13g2_nand3_1 _1198_ (.B(_0559_),
    .C(_0566_),
    .A(_0555_),
    .Y(_0567_));
 sg13g2_o21ai_1 _1199_ (.B1(_0481_),
    .Y(_0568_),
    .A1(_0482_),
    .A2(_0564_));
 sg13g2_xor2_1 _1200_ (.B(_0568_),
    .A(_0490_),
    .X(_0569_));
 sg13g2_nand2_2 _1201_ (.Y(_0570_),
    .A(_0567_),
    .B(_0569_));
 sg13g2_nand2b_1 _1202_ (.Y(_0571_),
    .B(_0529_),
    .A_N(_0522_));
 sg13g2_nand3_1 _1203_ (.B(net165),
    .C(_0571_),
    .A(_0530_),
    .Y(_0572_));
 sg13g2_and2_1 _1204_ (.A(net180),
    .B(_0569_),
    .X(_0573_));
 sg13g2_nand3_1 _1205_ (.B(_0560_),
    .C(_0561_),
    .A(net178),
    .Y(_0574_));
 sg13g2_nand2_1 _1206_ (.Y(_0575_),
    .A(_0563_),
    .B(_0565_));
 sg13g2_nor4_1 _1207_ (.A(_0555_),
    .B(_0559_),
    .C(_0574_),
    .D(_0575_),
    .Y(_0576_));
 sg13g2_or2_1 _1208_ (.X(_0577_),
    .B(_0576_),
    .A(_0573_));
 sg13g2_a22oi_1 _1209_ (.Y(_0059_),
    .B1(_0572_),
    .B2(net164),
    .A2(net189),
    .A1(_0166_));
 sg13g2_and2_1 _1210_ (.A(_0528_),
    .B(_0530_),
    .X(_0578_));
 sg13g2_xor2_1 _1211_ (.B(_0578_),
    .A(_0545_),
    .X(_0579_));
 sg13g2_nand2_1 _1212_ (.Y(_0580_),
    .A(net166),
    .B(_0579_));
 sg13g2_a22oi_1 _1213_ (.Y(_0060_),
    .B1(net164),
    .B2(_0580_),
    .A2(net190),
    .A1(_0165_));
 sg13g2_o21ai_1 _1214_ (.B1(_0533_),
    .Y(_0581_),
    .A1(_0542_),
    .A2(_0578_));
 sg13g2_nand2_1 _1215_ (.Y(_0582_),
    .A(_0536_),
    .B(_0581_));
 sg13g2_xor2_1 _1216_ (.B(_0581_),
    .A(_0536_),
    .X(_0583_));
 sg13g2_nand2_1 _1217_ (.Y(_0584_),
    .A(net166),
    .B(_0583_));
 sg13g2_a22oi_1 _1218_ (.Y(_0061_),
    .B1(net164),
    .B2(_0584_),
    .A2(net189),
    .A1(_0167_));
 sg13g2_nand2_1 _1219_ (.Y(_0585_),
    .A(_0535_),
    .B(_0582_));
 sg13g2_xor2_1 _1220_ (.B(_0585_),
    .A(_0541_),
    .X(_0586_));
 sg13g2_nand2_1 _1221_ (.Y(_0587_),
    .A(net166),
    .B(_0586_));
 sg13g2_a22oi_1 _1222_ (.Y(_0062_),
    .B1(net164),
    .B2(_0587_),
    .A2(net189),
    .A1(_0168_));
 sg13g2_nand2b_1 _1223_ (.Y(_0588_),
    .B(_0368_),
    .A_N(_0549_));
 sg13g2_nand2_1 _1224_ (.Y(_0589_),
    .A(_0369_),
    .B(_0549_));
 sg13g2_nand3_1 _1225_ (.B(_0588_),
    .C(_0589_),
    .A(net166),
    .Y(_0590_));
 sg13g2_a22oi_1 _1226_ (.Y(_0063_),
    .B1(net164),
    .B2(_0590_),
    .A2(net189),
    .A1(_0169_));
 sg13g2_o21ai_1 _1227_ (.B1(_0588_),
    .Y(_0591_),
    .A1(_0156_),
    .A2(_0158_));
 sg13g2_xnor2_1 _1228_ (.Y(_0592_),
    .A(_0380_),
    .B(_0591_));
 sg13g2_nand2_1 _1229_ (.Y(_0593_),
    .A(net166),
    .B(_0592_));
 sg13g2_a22oi_1 _1230_ (.Y(_0064_),
    .B1(net164),
    .B2(_0593_),
    .A2(net189),
    .A1(_0170_));
 sg13g2_o21ai_1 _1231_ (.B1(_0383_),
    .Y(_0594_),
    .A1(_0380_),
    .A2(_0588_));
 sg13g2_xnor2_1 _1232_ (.Y(_0595_),
    .A(_0387_),
    .B(_0594_));
 sg13g2_nand2_1 _1233_ (.Y(_0596_),
    .A(net166),
    .B(_0595_));
 sg13g2_a22oi_1 _1234_ (.Y(_0065_),
    .B1(net164),
    .B2(_0596_),
    .A2(net188),
    .A1(_0171_));
 sg13g2_a21oi_1 _1235_ (.A1(_0386_),
    .A2(_0594_),
    .Y(_0597_),
    .B1(_0385_));
 sg13g2_xnor2_1 _1236_ (.Y(_0598_),
    .A(_0391_),
    .B(_0597_));
 sg13g2_nand2b_1 _1237_ (.Y(_0599_),
    .B(net166),
    .A_N(_0598_));
 sg13g2_a22oi_1 _1238_ (.Y(_0066_),
    .B1(net163),
    .B2(_0599_),
    .A2(net188),
    .A1(_0173_));
 sg13g2_and2_1 _1239_ (.A(_0395_),
    .B(_0550_),
    .X(_0600_));
 sg13g2_xor2_1 _1240_ (.B(_0550_),
    .A(_0395_),
    .X(_0601_));
 sg13g2_nand2_1 _1241_ (.Y(_0602_),
    .A(net165),
    .B(_0601_));
 sg13g2_a22oi_1 _1242_ (.Y(_0067_),
    .B1(net163),
    .B2(_0602_),
    .A2(net187),
    .A1(_0175_));
 sg13g2_a21oi_1 _1243_ (.A1(net195),
    .A2(net125),
    .Y(_0603_),
    .B1(_0600_));
 sg13g2_xnor2_1 _1244_ (.Y(_0604_),
    .A(_0405_),
    .B(_0603_));
 sg13g2_nand2_1 _1245_ (.Y(_0605_),
    .A(net165),
    .B(_0604_));
 sg13g2_a22oi_1 _1246_ (.Y(_0068_),
    .B1(net163),
    .B2(_0605_),
    .A2(net187),
    .A1(_0177_));
 sg13g2_a21oi_1 _1247_ (.A1(_0405_),
    .A2(_0600_),
    .Y(_0606_),
    .B1(_0409_));
 sg13g2_xor2_1 _1248_ (.B(_0606_),
    .A(_0412_),
    .X(_0607_));
 sg13g2_nand2_1 _1249_ (.Y(_0608_),
    .A(net165),
    .B(_0607_));
 sg13g2_a22oi_1 _1250_ (.Y(_0069_),
    .B1(net163),
    .B2(_0608_),
    .A2(net187),
    .A1(_0179_));
 sg13g2_o21ai_1 _1251_ (.B1(_0411_),
    .Y(_0609_),
    .A1(_0412_),
    .A2(_0606_));
 sg13g2_xnor2_1 _1252_ (.Y(_0610_),
    .A(_0418_),
    .B(_0609_));
 sg13g2_nand2_1 _1253_ (.Y(_0611_),
    .A(net165),
    .B(_0610_));
 sg13g2_a22oi_1 _1254_ (.Y(_0070_),
    .B1(net163),
    .B2(_0611_),
    .A2(net188),
    .A1(_0180_));
 sg13g2_nor2b_1 _1255_ (.A(_0556_),
    .B_N(_0429_),
    .Y(_0612_));
 sg13g2_xnor2_1 _1256_ (.Y(_0613_),
    .A(_0429_),
    .B(_0556_));
 sg13g2_nand2_1 _1257_ (.Y(_0614_),
    .A(net165),
    .B(_0613_));
 sg13g2_a22oi_1 _1258_ (.Y(_0071_),
    .B1(net163),
    .B2(_0614_),
    .A2(net188),
    .A1(_0181_));
 sg13g2_nor2_1 _1259_ (.A(_0428_),
    .B(_0612_),
    .Y(_0615_));
 sg13g2_xnor2_1 _1260_ (.Y(_0616_),
    .A(_0433_),
    .B(_0615_));
 sg13g2_nand2_1 _1261_ (.Y(_0617_),
    .A(net165),
    .B(_0616_));
 sg13g2_a22oi_1 _1262_ (.Y(_0072_),
    .B1(net163),
    .B2(_0617_),
    .A2(net188),
    .A1(_0182_));
 sg13g2_xnor2_1 _1263_ (.Y(_0618_),
    .A(_0444_),
    .B(_0557_));
 sg13g2_nand2_1 _1264_ (.Y(_0619_),
    .A(net165),
    .B(_0618_));
 sg13g2_a22oi_1 _1265_ (.Y(_0073_),
    .B1(net163),
    .B2(_0619_),
    .A2(net187),
    .A1(_0184_));
 sg13g2_a21o_1 _1266_ (.A2(net191),
    .A1(net149),
    .B1(_0573_),
    .X(_0074_));
 sg13g2_nand2_1 _1267_ (.Y(_0620_),
    .A(fb_samp),
    .B(_0186_));
 sg13g2_nor2_1 _1268_ (.A(net56),
    .B(_0620_),
    .Y(_0621_));
 sg13g2_o21ai_1 _1269_ (.B1(net176),
    .Y(_0622_),
    .A1(net300),
    .A2(net172));
 sg13g2_inv_1 _1270_ (.Y(_0075_),
    .A(net301));
 sg13g2_mux2_1 _1271_ (.A0(net6),
    .A1(net329),
    .S(net241),
    .X(_0076_));
 sg13g2_nand2_1 _1272_ (.Y(_0623_),
    .A(net319),
    .B(net241));
 sg13g2_o21ai_1 _1273_ (.B1(_0623_),
    .Y(_0077_),
    .A1(net7),
    .A2(net241));
 sg13g2_mux2_1 _1274_ (.A0(\u_core.ref_samp_d ),
    .A1(net113),
    .S(net186),
    .X(_0078_));
 sg13g2_xor2_1 _1275_ (.B(net186),
    .A(net60),
    .X(_0079_));
 sg13g2_and3_2 _1276_ (.X(_0624_),
    .A(net60),
    .B(net89),
    .C(net186));
 sg13g2_a21oi_1 _1277_ (.A1(net60),
    .A2(net186),
    .Y(_0625_),
    .B1(net89));
 sg13g2_nor2_1 _1278_ (.A(_0624_),
    .B(_0625_),
    .Y(_0080_));
 sg13g2_xor2_1 _1279_ (.B(_0624_),
    .A(net71),
    .X(_0081_));
 sg13g2_nand3_1 _1280_ (.B(net326),
    .C(_0624_),
    .A(net71),
    .Y(_0626_));
 sg13g2_a21o_1 _1281_ (.A2(_0624_),
    .A1(net71),
    .B1(net326),
    .X(_0627_));
 sg13g2_and2_1 _1282_ (.A(_0626_),
    .B(_0627_),
    .X(_0082_));
 sg13g2_nor2_1 _1283_ (.A(_0163_),
    .B(_0626_),
    .Y(_0628_));
 sg13g2_xnor2_1 _1284_ (.Y(_0083_),
    .A(net46),
    .B(_0626_));
 sg13g2_nand4_1 _1285_ (.B(\u_core.beat_cnt[3] ),
    .C(net46),
    .A(net71),
    .Y(_0629_),
    .D(net64));
 sg13g2_xor2_1 _1286_ (.B(_0628_),
    .A(net64),
    .X(_0084_));
 sg13g2_a21oi_1 _1287_ (.A1(net64),
    .A2(_0628_),
    .Y(_0630_),
    .B1(net75));
 sg13g2_nand3_1 _1288_ (.B(net75),
    .C(_0628_),
    .A(net64),
    .Y(_0631_));
 sg13g2_nor2b_1 _1289_ (.A(net76),
    .B_N(_0631_),
    .Y(_0085_));
 sg13g2_nor2_1 _1290_ (.A(_0164_),
    .B(_0631_),
    .Y(_0632_));
 sg13g2_xnor2_1 _1291_ (.Y(_0086_),
    .A(net44),
    .B(_0631_));
 sg13g2_and2_1 _1292_ (.A(net48),
    .B(_0632_),
    .X(_0633_));
 sg13g2_xor2_1 _1293_ (.B(_0632_),
    .A(net48),
    .X(_0087_));
 sg13g2_xor2_1 _1294_ (.B(_0633_),
    .A(net62),
    .X(_0088_));
 sg13g2_nand3_1 _1295_ (.B(net44),
    .C(net48),
    .A(net75),
    .Y(_0634_));
 sg13g2_nand3_1 _1296_ (.B(net89),
    .C(net62),
    .A(net60),
    .Y(_0635_));
 sg13g2_nor4_2 _1297_ (.A(_0187_),
    .B(_0629_),
    .C(_0634_),
    .Y(_0636_),
    .D(_0635_));
 sg13g2_xor2_1 _1298_ (.B(_0636_),
    .A(net58),
    .X(_0089_));
 sg13g2_a21oi_1 _1299_ (.A1(net58),
    .A2(_0636_),
    .Y(_0637_),
    .B1(net104));
 sg13g2_nand4_1 _1300_ (.B(net58),
    .C(net104),
    .A(net62),
    .Y(_0638_),
    .D(_0633_));
 sg13g2_nor2b_1 _1301_ (.A(net105),
    .B_N(_0638_),
    .Y(_0090_));
 sg13g2_and4_1 _1302_ (.A(net58),
    .B(net334),
    .C(net66),
    .D(_0636_),
    .X(_0639_));
 sg13g2_xnor2_1 _1303_ (.Y(_0091_),
    .A(net66),
    .B(_0638_));
 sg13g2_xor2_1 _1304_ (.B(_0639_),
    .A(net54),
    .X(_0092_));
 sg13g2_a21oi_1 _1305_ (.A1(net54),
    .A2(_0639_),
    .Y(_0640_),
    .B1(net98));
 sg13g2_nand3_1 _1306_ (.B(net98),
    .C(_0639_),
    .A(net54),
    .Y(_0641_));
 sg13g2_nor2b_1 _1307_ (.A(net99),
    .B_N(_0641_),
    .Y(_0093_));
 sg13g2_xnor2_1 _1308_ (.Y(_0094_),
    .A(net50),
    .B(_0641_));
 sg13g2_nand2b_1 _1309_ (.Y(_0642_),
    .B(\u_core.t_ref[0] ),
    .A_N(\u_core.t_fb[0] ));
 sg13g2_nor2b_1 _1310_ (.A(\u_core.t_ref[1] ),
    .B_N(\u_core.t_fb[1] ),
    .Y(_0643_));
 sg13g2_xnor2_1 _1311_ (.Y(_0644_),
    .A(\u_core.t_fb[1] ),
    .B(\u_core.t_ref[1] ));
 sg13g2_nor2b_1 _1312_ (.A(\u_core.t_ref[2] ),
    .B_N(\u_core.t_fb[2] ),
    .Y(_0645_));
 sg13g2_nand2b_1 _1313_ (.Y(_0646_),
    .B(\u_core.t_ref[2] ),
    .A_N(\u_core.t_fb[2] ));
 sg13g2_a21o_1 _1314_ (.A2(_0644_),
    .A1(_0642_),
    .B1(_0643_),
    .X(_0647_));
 sg13g2_nor2_1 _1315_ (.A(net81),
    .B(net175),
    .Y(_0648_));
 sg13g2_nand2b_1 _1316_ (.Y(_0649_),
    .B(\u_core.t_fb[3] ),
    .A_N(\u_core.t_ref[3] ));
 sg13g2_xor2_1 _1317_ (.B(\u_core.t_ref[3] ),
    .A(\u_core.t_fb[3] ),
    .X(_0650_));
 sg13g2_a21oi_1 _1318_ (.A1(_0646_),
    .A2(_0647_),
    .Y(_0651_),
    .B1(_0645_));
 sg13g2_xnor2_1 _1319_ (.Y(_0652_),
    .A(_0650_),
    .B(_0651_));
 sg13g2_a21oi_1 _1320_ (.A1(net175),
    .A2(_0652_),
    .Y(_0095_),
    .B1(_0648_));
 sg13g2_nor2b_1 _1321_ (.A(net108),
    .B_N(net137),
    .Y(_0653_));
 sg13g2_nand2b_1 _1322_ (.Y(_0654_),
    .B(net108),
    .A_N(net137));
 sg13g2_nand2b_1 _1323_ (.Y(_0655_),
    .B(_0654_),
    .A_N(_0653_));
 sg13g2_o21ai_1 _1324_ (.B1(_0649_),
    .Y(_0656_),
    .A1(_0650_),
    .A2(_0651_));
 sg13g2_xnor2_1 _1325_ (.Y(_0657_),
    .A(_0655_),
    .B(_0656_));
 sg13g2_mux2_1 _1326_ (.A0(net245),
    .A1(_0657_),
    .S(net175),
    .X(_0096_));
 sg13g2_nor2_1 _1327_ (.A(net285),
    .B(net175),
    .Y(_0658_));
 sg13g2_a21oi_1 _1328_ (.A1(_0654_),
    .A2(_0656_),
    .Y(_0659_),
    .B1(_0653_));
 sg13g2_nor2_1 _1329_ (.A(\u_core.t_fb[5] ),
    .B(_0160_),
    .Y(_0660_));
 sg13g2_xor2_1 _1330_ (.B(net280),
    .A(\u_core.t_fb[5] ),
    .X(_0661_));
 sg13g2_xnor2_1 _1331_ (.Y(_0662_),
    .A(_0659_),
    .B(_0661_));
 sg13g2_a21oi_1 _1332_ (.A1(net175),
    .A2(_0662_),
    .Y(_0097_),
    .B1(_0658_));
 sg13g2_nand2b_1 _1333_ (.Y(_0663_),
    .B(net289),
    .A_N(\u_core.t_ref[6] ));
 sg13g2_xor2_1 _1334_ (.B(\u_core.t_ref[6] ),
    .A(\u_core.t_fb[6] ),
    .X(_0664_));
 sg13g2_a221oi_1 _1335_ (.B2(_0656_),
    .C1(_0653_),
    .B1(_0654_),
    .A1(\u_core.t_fb[5] ),
    .Y(_0665_),
    .A2(_0160_));
 sg13g2_or3_1 _1336_ (.A(_0660_),
    .B(_0664_),
    .C(_0665_),
    .X(_0666_));
 sg13g2_o21ai_1 _1337_ (.B1(_0664_),
    .Y(_0667_),
    .A1(_0660_),
    .A2(_0665_));
 sg13g2_and2_1 _1338_ (.A(_0666_),
    .B(_0667_),
    .X(_0668_));
 sg13g2_mux2_1 _1339_ (.A0(net317),
    .A1(_0668_),
    .S(net175),
    .X(_0098_));
 sg13g2_nand2b_1 _1340_ (.Y(_0669_),
    .B(net162),
    .A_N(net131));
 sg13g2_xnor2_1 _1341_ (.Y(_0670_),
    .A(\u_core.t_fb[7] ),
    .B(\u_core.t_ref[7] ));
 sg13g2_inv_1 _1342_ (.Y(_0671_),
    .A(_0670_));
 sg13g2_a21o_1 _1343_ (.A2(_0666_),
    .A1(_0663_),
    .B1(_0671_),
    .X(_0672_));
 sg13g2_nand3_1 _1344_ (.B(_0666_),
    .C(_0671_),
    .A(_0663_),
    .Y(_0673_));
 sg13g2_and3_1 _1345_ (.X(_0674_),
    .A(net174),
    .B(_0672_),
    .C(_0673_));
 sg13g2_a21o_1 _1346_ (.A2(net176),
    .A1(net307),
    .B1(_0674_),
    .X(_0099_));
 sg13g2_nor2b_1 _1347_ (.A(net292),
    .B_N(net311),
    .Y(_0675_));
 sg13g2_xor2_1 _1348_ (.B(\u_core.t_ref[8] ),
    .A(\u_core.t_fb[8] ),
    .X(_0676_));
 sg13g2_a21o_1 _1349_ (.A2(_0672_),
    .A1(_0669_),
    .B1(_0676_),
    .X(_0677_));
 sg13g2_nand3_1 _1350_ (.B(_0672_),
    .C(_0676_),
    .A(_0669_),
    .Y(_0678_));
 sg13g2_a21oi_1 _1351_ (.A1(_0677_),
    .A2(_0678_),
    .Y(_0679_),
    .B1(net176));
 sg13g2_a21oi_1 _1352_ (.A1(_0159_),
    .A2(net176),
    .Y(_0100_),
    .B1(_0679_));
 sg13g2_nor2_1 _1353_ (.A(net313),
    .B(net175),
    .Y(_0680_));
 sg13g2_xor2_1 _1354_ (.B(net150),
    .A(net155),
    .X(_0681_));
 sg13g2_nor2b_1 _1355_ (.A(_0675_),
    .B_N(_0677_),
    .Y(_0682_));
 sg13g2_xnor2_1 _1356_ (.Y(_0683_),
    .A(_0681_),
    .B(_0682_));
 sg13g2_a21oi_1 _1357_ (.A1(net174),
    .A2(_0683_),
    .Y(_0101_),
    .B1(_0680_));
 sg13g2_nor2b_1 _1358_ (.A(net299),
    .B_N(net310),
    .Y(_0684_));
 sg13g2_xnor2_1 _1359_ (.Y(_0685_),
    .A(net310),
    .B(net299));
 sg13g2_a21oi_1 _1360_ (.A1(\u_core.t_fb[9] ),
    .A2(_0162_),
    .Y(_0686_),
    .B1(_0675_));
 sg13g2_a22oi_1 _1361_ (.Y(_0687_),
    .B1(_0677_),
    .B2(_0686_),
    .A2(\u_core.t_ref[9] ),
    .A1(_0161_));
 sg13g2_o21ai_1 _1362_ (.B1(net174),
    .Y(_0688_),
    .A1(_0685_),
    .A2(_0687_));
 sg13g2_a21oi_1 _1363_ (.A1(_0685_),
    .A2(_0687_),
    .Y(_0689_),
    .B1(_0688_));
 sg13g2_a21o_1 _1364_ (.A2(_0188_),
    .A1(net320),
    .B1(_0689_),
    .X(_0102_));
 sg13g2_nor2_1 _1365_ (.A(net203),
    .B(net173),
    .Y(_0690_));
 sg13g2_nor2b_1 _1366_ (.A(net258),
    .B_N(\u_core.t_fb[11] ),
    .Y(_0691_));
 sg13g2_nand2b_1 _1367_ (.Y(_0692_),
    .B(\u_core.t_ref[11] ),
    .A_N(\u_core.t_fb[11] ));
 sg13g2_nor2b_1 _1368_ (.A(_0691_),
    .B_N(_0692_),
    .Y(_0693_));
 sg13g2_a21oi_1 _1369_ (.A1(_0685_),
    .A2(_0687_),
    .Y(_0694_),
    .B1(_0684_));
 sg13g2_xor2_1 _1370_ (.B(_0694_),
    .A(_0693_),
    .X(_0695_));
 sg13g2_a21oi_1 _1371_ (.A1(net173),
    .A2(_0695_),
    .Y(_0103_),
    .B1(_0690_));
 sg13g2_nand2b_1 _1372_ (.Y(_0696_),
    .B(net294),
    .A_N(\u_core.t_ref[12] ));
 sg13g2_nor2b_1 _1373_ (.A(\u_core.t_fb[12] ),
    .B_N(\u_core.t_ref[12] ),
    .Y(_0697_));
 sg13g2_xnor2_1 _1374_ (.Y(_0698_),
    .A(net294),
    .B(net314));
 sg13g2_and2_1 _1375_ (.A(_0685_),
    .B(_0693_),
    .X(_0699_));
 sg13g2_a221oi_1 _1376_ (.B2(_0687_),
    .C1(_0691_),
    .B1(_0699_),
    .A1(_0684_),
    .Y(_0700_),
    .A2(_0692_));
 sg13g2_xnor2_1 _1377_ (.Y(_0701_),
    .A(_0698_),
    .B(_0700_));
 sg13g2_mux2_1 _1378_ (.A0(net202),
    .A1(_0701_),
    .S(net173),
    .X(_0104_));
 sg13g2_nor2_1 _1379_ (.A(net322),
    .B(net173),
    .Y(_0702_));
 sg13g2_o21ai_1 _1380_ (.B1(_0696_),
    .Y(_0703_),
    .A1(_0697_),
    .A2(_0700_));
 sg13g2_nor2b_1 _1381_ (.A(net284),
    .B_N(net255),
    .Y(_0704_));
 sg13g2_nand2b_1 _1382_ (.Y(_0705_),
    .B(net284),
    .A_N(net255));
 sg13g2_nor2b_1 _1383_ (.A(_0704_),
    .B_N(_0705_),
    .Y(_0706_));
 sg13g2_xnor2_1 _1384_ (.Y(_0707_),
    .A(_0703_),
    .B(_0706_));
 sg13g2_a21oi_1 _1385_ (.A1(net173),
    .A2(_0707_),
    .Y(_0105_),
    .B1(_0702_));
 sg13g2_nor2_1 _1386_ (.A(net201),
    .B(net173),
    .Y(_0708_));
 sg13g2_nand2b_1 _1387_ (.Y(_0709_),
    .B(net302),
    .A_N(net277));
 sg13g2_xor2_1 _1388_ (.B(net277),
    .A(net302),
    .X(_0710_));
 sg13g2_a21oi_1 _1389_ (.A1(_0703_),
    .A2(_0705_),
    .Y(_0711_),
    .B1(_0704_));
 sg13g2_xnor2_1 _1390_ (.Y(_0712_),
    .A(_0710_),
    .B(_0711_));
 sg13g2_a21oi_1 _1391_ (.A1(net173),
    .A2(_0712_),
    .Y(_0106_),
    .B1(_0708_));
 sg13g2_o21ai_1 _1392_ (.B1(_0709_),
    .Y(_0713_),
    .A1(_0710_),
    .A2(_0711_));
 sg13g2_xnor2_1 _1393_ (.Y(_0714_),
    .A(net250),
    .B(net143));
 sg13g2_nand2_1 _1394_ (.Y(_0715_),
    .A(net200),
    .B(net176));
 sg13g2_xnor2_1 _1395_ (.Y(_0716_),
    .A(_0713_),
    .B(_0714_));
 sg13g2_o21ai_1 _1396_ (.B1(_0715_),
    .Y(_0107_),
    .A1(net176),
    .A2(_0716_));
 sg13g2_nor3_1 _1397_ (.A(_0154_),
    .B(\u_core.ref_samp_d ),
    .C(_0187_),
    .Y(_0717_));
 sg13g2_mux2_1 _1398_ (.A0(net119),
    .A1(net60),
    .S(net168),
    .X(_0108_));
 sg13g2_mux2_1 _1399_ (.A0(net304),
    .A1(net89),
    .S(net168),
    .X(_0109_));
 sg13g2_mux2_1 _1400_ (.A0(net257),
    .A1(net71),
    .S(net168),
    .X(_0110_));
 sg13g2_mux2_1 _1401_ (.A0(net290),
    .A1(\u_core.beat_cnt[3] ),
    .S(net168),
    .X(_0111_));
 sg13g2_nor2_1 _1402_ (.A(net108),
    .B(net168),
    .Y(_0144_));
 sg13g2_a21oi_1 _1403_ (.A1(_0163_),
    .A2(net168),
    .Y(_0112_),
    .B1(net109));
 sg13g2_nand2_1 _1404_ (.Y(_0145_),
    .A(net64),
    .B(net168));
 sg13g2_o21ai_1 _1405_ (.B1(_0145_),
    .Y(_0113_),
    .A1(_0160_),
    .A2(net169));
 sg13g2_mux2_1 _1406_ (.A0(net283),
    .A1(net75),
    .S(net168),
    .X(_0114_));
 sg13g2_nor2_1 _1407_ (.A(net131),
    .B(net167),
    .Y(_0146_));
 sg13g2_a21oi_1 _1408_ (.A1(_0164_),
    .A2(net167),
    .Y(_0115_),
    .B1(net132));
 sg13g2_mux2_1 _1409_ (.A0(net292),
    .A1(net48),
    .S(net167),
    .X(_0116_));
 sg13g2_nand2_1 _1410_ (.Y(_0147_),
    .A(net62),
    .B(net169));
 sg13g2_o21ai_1 _1411_ (.B1(_0147_),
    .Y(_0117_),
    .A1(_0162_),
    .A2(net169));
 sg13g2_mux2_1 _1412_ (.A0(net299),
    .A1(net58),
    .S(net167),
    .X(_0118_));
 sg13g2_mux2_1 _1413_ (.A0(net258),
    .A1(net104),
    .S(net167),
    .X(_0119_));
 sg13g2_mux2_1 _1414_ (.A0(net314),
    .A1(net66),
    .S(net169),
    .X(_0120_));
 sg13g2_mux2_1 _1415_ (.A0(net284),
    .A1(net54),
    .S(net167),
    .X(_0121_));
 sg13g2_mux2_1 _1416_ (.A0(net277),
    .A1(net98),
    .S(net167),
    .X(_0122_));
 sg13g2_mux2_1 _1417_ (.A0(net143),
    .A1(net50),
    .S(net167),
    .X(_0123_));
 sg13g2_mux2_1 _1418_ (.A0(fb_samp),
    .A1(net68),
    .S(_0186_),
    .X(_0124_));
 sg13g2_mux2_1 _1419_ (.A0(net120),
    .A1(net60),
    .S(net171),
    .X(_0125_));
 sg13g2_mux2_1 _1420_ (.A0(net297),
    .A1(net89),
    .S(net171),
    .X(_0126_));
 sg13g2_mux2_1 _1421_ (.A0(net259),
    .A1(net71),
    .S(net171),
    .X(_0127_));
 sg13g2_mux2_1 _1422_ (.A0(net308),
    .A1(\u_core.beat_cnt[3] ),
    .S(net171),
    .X(_0128_));
 sg13g2_nor2_1 _1423_ (.A(net137),
    .B(net171),
    .Y(_0148_));
 sg13g2_a21oi_1 _1424_ (.A1(_0163_),
    .A2(net171),
    .Y(_0129_),
    .B1(_0148_));
 sg13g2_mux2_1 _1425_ (.A0(net293),
    .A1(net64),
    .S(net171),
    .X(_0130_));
 sg13g2_mux2_1 _1426_ (.A0(net289),
    .A1(net75),
    .S(net171),
    .X(_0131_));
 sg13g2_nor2_1 _1427_ (.A(net162),
    .B(net170),
    .Y(_0149_));
 sg13g2_a21oi_1 _1428_ (.A1(_0164_),
    .A2(net170),
    .Y(_0132_),
    .B1(_0149_));
 sg13g2_mux2_1 _1429_ (.A0(net311),
    .A1(net48),
    .S(net170),
    .X(_0133_));
 sg13g2_nand2_1 _1430_ (.Y(_0150_),
    .A(net62),
    .B(net172));
 sg13g2_o21ai_1 _1431_ (.B1(_0150_),
    .Y(_0134_),
    .A1(_0161_),
    .A2(net170));
 sg13g2_mux2_1 _1432_ (.A0(net310),
    .A1(net58),
    .S(net170),
    .X(_0135_));
 sg13g2_mux2_1 _1433_ (.A0(net159),
    .A1(net104),
    .S(net170),
    .X(_0136_));
 sg13g2_mux2_1 _1434_ (.A0(net294),
    .A1(net66),
    .S(net172),
    .X(_0137_));
 sg13g2_mux2_1 _1435_ (.A0(net255),
    .A1(net54),
    .S(net170),
    .X(_0138_));
 sg13g2_mux2_1 _1436_ (.A0(net302),
    .A1(net98),
    .S(net172),
    .X(_0139_));
 sg13g2_mux2_1 _1437_ (.A0(net250),
    .A1(net50),
    .S(net170),
    .X(_0140_));
 sg13g2_nand2_1 _1438_ (.Y(_0151_),
    .A(net34),
    .B(_0186_));
 sg13g2_o21ai_1 _1439_ (.B1(net35),
    .Y(_0141_),
    .A1(_0154_),
    .A2(net186));
 sg13g2_o21ai_1 _1440_ (.B1(_0620_),
    .Y(_0142_),
    .A1(_0155_),
    .A2(net186));
 sg13g2_o21ai_1 _1441_ (.B1(net176),
    .Y(_0152_),
    .A1(net261),
    .A2(net169));
 sg13g2_inv_1 _1442_ (.Y(_0143_),
    .A(net262));
 sg13g2_dfrbpq_1 _1443_ (.RESET_B(net227),
    .D(net33),
    .Q(\nco_phase_acc[0] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1444_ (.RESET_B(net227),
    .D(net122),
    .Q(\nco_phase_acc[1] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net227),
    .D(net80),
    .Q(\nco_phase_acc[2] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net227),
    .D(net101),
    .Q(\nco_phase_acc[3] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net223),
    .D(net95),
    .Q(\nco_phase_acc[4] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_2 _1448_ (.RESET_B(net223),
    .D(net118),
    .Q(\nco_phase_acc[5] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1449_ (.RESET_B(net223),
    .D(net111),
    .Q(\nco_phase_acc[6] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net224),
    .D(net103),
    .Q(\nco_phase_acc[7] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1451_ (.RESET_B(net221),
    .D(net288),
    .Q(\nco_phase_acc[8] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_2 _1452_ (.RESET_B(net222),
    .D(net252),
    .Q(\nco_phase_acc[9] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1453_ (.RESET_B(net222),
    .D(net84),
    .Q(\nco_phase_acc[10] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1454_ (.RESET_B(net222),
    .D(net134),
    .Q(\nco_phase_acc[11] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_1 _1455_ (.RESET_B(net222),
    .D(net93),
    .Q(\nco_phase_acc[12] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1456_ (.RESET_B(net221),
    .D(net145),
    .Q(\nco_phase_acc[13] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1457_ (.RESET_B(net221),
    .D(net91),
    .Q(\nco_phase_acc[14] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1458_ (.RESET_B(net223),
    .D(net74),
    .Q(\nco_phase_acc[15] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _1459_ (.RESET_B(net223),
    .D(_0019_),
    .Q(\nco_phase_acc[16] ),
    .CLK(clknet_5_23__leaf_clk));
 sg13g2_dfrbpq_1 _1460_ (.RESET_B(net227),
    .D(net41),
    .Q(\nco_phase_acc[17] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1461_ (.RESET_B(net229),
    .D(net39),
    .Q(\nco_phase_acc[18] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1462_ (.RESET_B(net229),
    .D(net43),
    .Q(\nco_phase_acc[19] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1463_ (.RESET_B(net229),
    .D(net29),
    .Q(\nco_phase_acc[20] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1464_ (.RESET_B(net229),
    .D(_0024_),
    .Q(\nco_phase_acc[21] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_1 _1465_ (.RESET_B(net229),
    .D(net31),
    .Q(\nco_phase_acc[22] ),
    .CLK(clknet_5_31__leaf_clk));
 sg13g2_dfrbpq_2 _1466_ (.RESET_B(net229),
    .D(_0026_),
    .Q(clk_helper),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_2 _1467_ (.RESET_B(net232),
    .D(_0027_),
    .Q(\u_lf.kp_sel_latched[0] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1468_ (.RESET_B(net231),
    .D(_0028_),
    .Q(_0001_),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1469_ (.RESET_B(net226),
    .D(net53),
    .Q(\u_lf.i_acc[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_2 _1470_ (.RESET_B(net226),
    .D(_0030_),
    .Q(\u_lf.i_acc[1] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1471_ (.RESET_B(net226),
    .D(net154),
    .Q(\u_lf.i_acc[2] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1472_ (.RESET_B(net226),
    .D(_0032_),
    .Q(\u_lf.i_acc[3] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1473_ (.RESET_B(net231),
    .D(_0033_),
    .Q(\u_lf.i_acc[4] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1474_ (.RESET_B(net231),
    .D(_0034_),
    .Q(\u_lf.i_acc[5] ),
    .CLK(clknet_5_27__leaf_clk));
 sg13g2_dfrbpq_2 _1475_ (.RESET_B(net228),
    .D(net276),
    .Q(\u_lf.i_acc[6] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1476_ (.RESET_B(net228),
    .D(net249),
    .Q(\u_lf.i_acc[7] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _1477_ (.RESET_B(net226),
    .D(_0037_),
    .Q(\u_lf.i_acc[8] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1478_ (.RESET_B(net226),
    .D(_0038_),
    .Q(\u_lf.i_acc[9] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1479_ (.RESET_B(net226),
    .D(net265),
    .Q(\u_lf.i_acc[10] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_2 _1480_ (.RESET_B(net226),
    .D(_0040_),
    .Q(\u_lf.i_acc[11] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1481_ (.RESET_B(net220),
    .D(_0041_),
    .Q(\u_lf.i_acc[12] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1482_ (.RESET_B(net225),
    .D(net244),
    .Q(\u_lf.i_acc[13] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1483_ (.RESET_B(net225),
    .D(_0043_),
    .Q(\u_lf.i_acc[14] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1484_ (.RESET_B(net225),
    .D(net267),
    .Q(\u_lf.i_acc[15] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_2 _1485_ (.RESET_B(net220),
    .D(net126),
    .Q(\u_lf.i_acc[16] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1486_ (.RESET_B(net220),
    .D(net161),
    .Q(\u_lf.i_acc[17] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1487_ (.RESET_B(net220),
    .D(_0047_),
    .Q(\u_lf.i_acc[18] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1488_ (.RESET_B(net220),
    .D(_0048_),
    .Q(\u_lf.i_acc[19] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_2 _1489_ (.RESET_B(net220),
    .D(_0049_),
    .Q(\u_lf.i_acc[20] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net220),
    .D(net142),
    .Q(\u_lf.i_acc[21] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1491_ (.RESET_B(net211),
    .D(_0051_),
    .Q(\u_lf.i_acc[22] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net211),
    .D(net158),
    .Q(\u_lf.i_acc[23] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_2 _1493_ (.RESET_B(net211),
    .D(net274),
    .Q(\u_lf.i_acc[24] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1494_ (.RESET_B(net211),
    .D(net148),
    .Q(\u_lf.i_acc[25] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_2 _1495_ (.RESET_B(net211),
    .D(_0055_),
    .Q(\u_lf.i_acc[26] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1496_ (.RESET_B(net211),
    .D(net254),
    .Q(\u_lf.i_acc[27] ),
    .CLK(clknet_5_4__leaf_clk));
 sg13g2_dfrbpq_1 _1497_ (.RESET_B(net210),
    .D(_0057_),
    .Q(\u_lf.i_acc[28] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1498_ (.RESET_B(net211),
    .D(net107),
    .Q(\u_lf.i_acc[29] ),
    .CLK(clknet_5_5__leaf_clk));
 sg13g2_dfrbpq_1 _1499_ (.RESET_B(net228),
    .D(net88),
    .Q(\ctrl[8] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_1 _1500_ (.RESET_B(net227),
    .D(net130),
    .Q(\ctrl[9] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1501_ (.RESET_B(net227),
    .D(net124),
    .Q(\ctrl[10] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net227),
    .D(net128),
    .Q(\ctrl[11] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_1 _1503_ (.RESET_B(net223),
    .D(net78),
    .Q(\ctrl[12] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_2 _1504_ (.RESET_B(net224),
    .D(net139),
    .Q(\ctrl[13] ),
    .CLK(clknet_5_22__leaf_clk));
 sg13g2_dfrbpq_1 _1505_ (.RESET_B(net223),
    .D(net269),
    .Q(\ctrl[14] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1506_ (.RESET_B(net223),
    .D(net136),
    .Q(\ctrl[15] ),
    .CLK(clknet_5_19__leaf_clk));
 sg13g2_dfrbpq_1 _1507_ (.RESET_B(net222),
    .D(_0067_),
    .Q(\ctrl[16] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net222),
    .D(_0068_),
    .Q(\ctrl[17] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1509_ (.RESET_B(net221),
    .D(_0069_),
    .Q(\ctrl[18] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_1 _1510_ (.RESET_B(net221),
    .D(net97),
    .Q(\ctrl[19] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1511_ (.RESET_B(net221),
    .D(net116),
    .Q(\ctrl[20] ),
    .CLK(clknet_5_16__leaf_clk));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net221),
    .D(_0072_),
    .Q(\ctrl[21] ),
    .CLK(clknet_5_20__leaf_clk));
 sg13g2_dfrbpq_2 _1513_ (.RESET_B(net221),
    .D(_0073_),
    .Q(\ctrl[22] ),
    .CLK(clknet_5_17__leaf_clk));
 sg13g2_dfrbpq_2 _1514_ (.RESET_B(net220),
    .D(_0074_),
    .Q(\ctrl[23] ),
    .CLK(clknet_5_18__leaf_clk));
 sg13g2_dfrbpq_1 _1515_ (.RESET_B(net218),
    .D(_0075_),
    .Q(\u_core.have_fb ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_2 _1516_ (.RESET_B(net231),
    .D(_0076_),
    .Q(\u_lf.ki_sel_latched[0] ),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_2 _1517_ (.RESET_B(net231),
    .D(_0077_),
    .Q(_0002_),
    .CLK(clknet_5_25__leaf_clk));
 sg13g2_dfrbpq_1 _1518_ (.RESET_B(net229),
    .D(net26),
    .Q(helper_msb_d),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1519_ (.RESET_B(net216),
    .D(net114),
    .Q(\u_core.ref_samp_d ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_2 _1520_ (.RESET_B(net214),
    .D(net61),
    .Q(\u_core.beat_cnt[0] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1521_ (.RESET_B(net214),
    .D(_0080_),
    .Q(\u_core.beat_cnt[1] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _1522_ (.RESET_B(net214),
    .D(net72),
    .Q(\u_core.beat_cnt[2] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1523_ (.RESET_B(net214),
    .D(_0082_),
    .Q(\u_core.beat_cnt[3] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1524_ (.RESET_B(net214),
    .D(net47),
    .Q(\u_core.beat_cnt[4] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _1525_ (.RESET_B(net213),
    .D(net65),
    .Q(\u_core.beat_cnt[5] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_2 _1526_ (.RESET_B(net213),
    .D(_0085_),
    .Q(\u_core.beat_cnt[6] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1527_ (.RESET_B(net213),
    .D(net45),
    .Q(\u_core.beat_cnt[7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1528_ (.RESET_B(net212),
    .D(net49),
    .Q(\u_core.beat_cnt[8] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_2 _1529_ (.RESET_B(net212),
    .D(net63),
    .Q(\u_core.beat_cnt[9] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1530_ (.RESET_B(net209),
    .D(net59),
    .Q(\u_core.beat_cnt[10] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1531_ (.RESET_B(net209),
    .D(_0090_),
    .Q(\u_core.beat_cnt[11] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_2 _1532_ (.RESET_B(net209),
    .D(net67),
    .Q(\u_core.beat_cnt[12] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1533_ (.RESET_B(net208),
    .D(net55),
    .Q(\u_core.beat_cnt[13] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _1534_ (.RESET_B(net208),
    .D(_0093_),
    .Q(\u_core.beat_cnt[14] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1535_ (.RESET_B(net208),
    .D(net51),
    .Q(\u_core.beat_cnt[15] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1536_ (.RESET_B(net217),
    .D(net82),
    .Q(\phase_err_beat[3] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1537_ (.RESET_B(net217),
    .D(_0096_),
    .Q(\phase_err_beat[4] ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1538_ (.RESET_B(net217),
    .D(net286),
    .Q(\phase_err_beat[5] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1539_ (.RESET_B(net217),
    .D(_0098_),
    .Q(\phase_err_beat[6] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1540_ (.RESET_B(net217),
    .D(_0099_),
    .Q(\phase_err_beat[7] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1541_ (.RESET_B(net217),
    .D(net247),
    .Q(\phase_err_beat[8] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1542_ (.RESET_B(net219),
    .D(_0101_),
    .Q(\phase_err_beat[9] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_2 _1543_ (.RESET_B(net218),
    .D(net321),
    .Q(\phase_err_beat[10] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1544_ (.RESET_B(net218),
    .D(_0103_),
    .Q(\phase_err_beat[11] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1545_ (.RESET_B(net218),
    .D(_0104_),
    .Q(\phase_err_beat[12] ),
    .CLK(clknet_5_13__leaf_clk));
 sg13g2_dfrbpq_2 _1546_ (.RESET_B(net218),
    .D(net323),
    .Q(\phase_err_beat[13] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1547_ (.RESET_B(net218),
    .D(_0106_),
    .Q(\phase_err_beat[14] ),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_2 _1548_ (.RESET_B(net210),
    .D(_0107_),
    .Q(\phase_err_beat[15] ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_dfrbpq_1 _1549_ (.RESET_B(net214),
    .D(_0108_),
    .Q(\u_core.t_ref[0] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1550_ (.RESET_B(net214),
    .D(_0109_),
    .Q(\u_core.t_ref[1] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_1 _1551_ (.RESET_B(net215),
    .D(_0110_),
    .Q(\u_core.t_ref[2] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1552_ (.RESET_B(net216),
    .D(net291),
    .Q(\u_core.t_ref[3] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1553_ (.RESET_B(net216),
    .D(_0112_),
    .Q(\u_core.t_ref[4] ),
    .CLK(clknet_5_9__leaf_clk));
 sg13g2_dfrbpq_1 _1554_ (.RESET_B(net216),
    .D(net281),
    .Q(\u_core.t_ref[5] ),
    .CLK(clknet_5_12__leaf_clk));
 sg13g2_dfrbpq_1 _1555_ (.RESET_B(net212),
    .D(_0114_),
    .Q(\u_core.t_ref[6] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1556_ (.RESET_B(net212),
    .D(_0115_),
    .Q(\u_core.t_ref[7] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1557_ (.RESET_B(net212),
    .D(_0116_),
    .Q(\u_core.t_ref[8] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1558_ (.RESET_B(net213),
    .D(net151),
    .Q(\u_core.t_ref[9] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1559_ (.RESET_B(net208),
    .D(_0118_),
    .Q(\u_core.t_ref[10] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1560_ (.RESET_B(net208),
    .D(_0119_),
    .Q(\u_core.t_ref[11] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _1561_ (.RESET_B(net210),
    .D(net315),
    .Q(\u_core.t_ref[12] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1562_ (.RESET_B(net210),
    .D(_0121_),
    .Q(\u_core.t_ref[13] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1563_ (.RESET_B(net210),
    .D(_0122_),
    .Q(\u_core.t_ref[14] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1564_ (.RESET_B(net208),
    .D(_0123_),
    .Q(\u_core.t_ref[15] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_1 _1565_ (.RESET_B(net229),
    .D(clk_fb),
    .Q(\u_core.fb_sync[0] ),
    .CLK(clknet_5_30__leaf_clk));
 sg13g2_dfrbpq_1 _1566_ (.RESET_B(net230),
    .D(net24),
    .Q(\u_core.fb_sync[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1567_ (.RESET_B(net230),
    .D(net1),
    .Q(\u_core.ref_sync[0] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1568_ (.RESET_B(net230),
    .D(net25),
    .Q(\u_core.ref_sync[1] ),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1569_ (.RESET_B(net230),
    .D(net69),
    .Q(fb_samp),
    .CLK(clknet_5_26__leaf_clk));
 sg13g2_dfrbpq_1 _1570_ (.RESET_B(net215),
    .D(_0125_),
    .Q(\u_core.t_fb[0] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1571_ (.RESET_B(net215),
    .D(_0126_),
    .Q(\u_core.t_fb[1] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1572_ (.RESET_B(net215),
    .D(_0127_),
    .Q(\u_core.t_fb[2] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1573_ (.RESET_B(net216),
    .D(net309),
    .Q(\u_core.t_fb[3] ),
    .CLK(clknet_5_14__leaf_clk));
 sg13g2_dfrbpq_1 _1574_ (.RESET_B(net214),
    .D(_0129_),
    .Q(\u_core.t_fb[4] ),
    .CLK(clknet_5_10__leaf_clk));
 sg13g2_dfrbpq_2 _1575_ (.RESET_B(net216),
    .D(_0130_),
    .Q(\u_core.t_fb[5] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1576_ (.RESET_B(net212),
    .D(_0131_),
    .Q(\u_core.t_fb[6] ),
    .CLK(clknet_5_11__leaf_clk));
 sg13g2_dfrbpq_1 _1577_ (.RESET_B(net212),
    .D(_0132_),
    .Q(\u_core.t_fb[7] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _1578_ (.RESET_B(net212),
    .D(_0133_),
    .Q(\u_core.t_fb[8] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1579_ (.RESET_B(net213),
    .D(net156),
    .Q(\u_core.t_fb[9] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_1 _1580_ (.RESET_B(net208),
    .D(_0135_),
    .Q(\u_core.t_fb[10] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1581_ (.RESET_B(net209),
    .D(_0136_),
    .Q(\u_core.t_fb[11] ),
    .CLK(clknet_5_3__leaf_clk));
 sg13g2_dfrbpq_2 _1582_ (.RESET_B(net210),
    .D(net295),
    .Q(\u_core.t_fb[12] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1583_ (.RESET_B(net210),
    .D(_0138_),
    .Q(\u_core.t_fb[13] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1584_ (.RESET_B(net210),
    .D(net303),
    .Q(\u_core.t_fb[14] ),
    .CLK(clknet_5_6__leaf_clk));
 sg13g2_dfrbpq_1 _1585_ (.RESET_B(net208),
    .D(_0140_),
    .Q(\u_core.t_fb[15] ),
    .CLK(clknet_5_1__leaf_clk));
 sg13g2_dfrbpq_1 _1586_ (.RESET_B(net217),
    .D(net36),
    .Q(ref_samp),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1587_ (.RESET_B(net217),
    .D(net57),
    .Q(\u_core.fb_samp_d ),
    .CLK(clknet_5_15__leaf_clk));
 sg13g2_dfrbpq_1 _1588_ (.RESET_B(net218),
    .D(net173),
    .Q(phase_valid),
    .CLK(clknet_5_24__leaf_clk));
 sg13g2_dfrbpq_1 _1589_ (.RESET_B(net218),
    .D(_0143_),
    .Q(\u_core.have_ref ),
    .CLK(clknet_5_7__leaf_clk));
 sg13g2_tielo tt_um_arthfink_ddmtd_9 (.L_LO(net9));
 sg13g2_tielo tt_um_arthfink_ddmtd_10 (.L_LO(net10));
 sg13g2_tielo tt_um_arthfink_ddmtd_11 (.L_LO(net11));
 sg13g2_tielo tt_um_arthfink_ddmtd_12 (.L_LO(net12));
 sg13g2_tielo tt_um_arthfink_ddmtd_13 (.L_LO(net13));
 sg13g2_tielo tt_um_arthfink_ddmtd_14 (.L_LO(net14));
 sg13g2_tielo tt_um_arthfink_ddmtd_15 (.L_LO(net15));
 sg13g2_tielo tt_um_arthfink_ddmtd_16 (.L_LO(net16));
 sg13g2_tielo tt_um_arthfink_ddmtd_17 (.L_LO(net17));
 sg13g2_tielo tt_um_arthfink_ddmtd_18 (.L_LO(net18));
 sg13g2_tielo tt_um_arthfink_ddmtd_19 (.L_LO(net19));
 sg13g2_tielo tt_um_arthfink_ddmtd_20 (.L_LO(net20));
 sg13g2_tielo tt_um_arthfink_ddmtd_21 (.L_LO(net21));
 sg13g2_tielo tt_um_arthfink_ddmtd_22 (.L_LO(net22));
 sg13g2_tielo tt_um_arthfink_ddmtd_23 (.L_LO(net23));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 fanout163 (.A(_0577_),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(_0577_),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(_0570_),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(_0570_),
    .X(net166));
 sg13g2_buf_8 fanout167 (.A(net169),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net169),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(_0717_),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net172),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net172),
    .X(net171));
 sg13g2_buf_8 fanout172 (.A(_0621_),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_1 fanout174 (.A(net175),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(_0000_),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(_0188_),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(net180),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net180),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(net180),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(net182),
    .X(net180));
 sg13g2_buf_8 fanout181 (.A(net182),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(net184),
    .X(net182));
 sg13g2_buf_8 fanout183 (.A(uo_out[0]),
    .X(net183));
 sg13g2_buf_8 fanout184 (.A(net185),
    .X(uo_out[0]));
 sg13g2_buf_8 fanout185 (.A(net184),
    .X(net185));
 sg13g2_buf_8 fanout186 (.A(_0186_),
    .X(net186));
 sg13g2_buf_8 fanout187 (.A(net188),
    .X(net187));
 sg13g2_buf_8 fanout188 (.A(net191),
    .X(net188));
 sg13g2_buf_8 fanout189 (.A(net191),
    .X(net189));
 sg13g2_buf_1 fanout190 (.A(net191),
    .X(net190));
 sg13g2_buf_8 fanout191 (.A(_0189_),
    .X(net191));
 sg13g2_buf_8 fanout192 (.A(net193),
    .X(net192));
 sg13g2_buf_8 fanout193 (.A(net197),
    .X(net193));
 sg13g2_buf_8 fanout194 (.A(net195),
    .X(net194));
 sg13g2_buf_8 fanout195 (.A(net197),
    .X(net195));
 sg13g2_buf_8 fanout196 (.A(net197),
    .X(net196));
 sg13g2_buf_8 fanout197 (.A(\phase_err_beat[15] ),
    .X(net197));
 sg13g2_buf_8 fanout198 (.A(net200),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(net200),
    .X(net199));
 sg13g2_buf_8 fanout200 (.A(net328),
    .X(net200));
 sg13g2_buf_8 fanout201 (.A(net331),
    .X(net201));
 sg13g2_buf_8 fanout202 (.A(net332),
    .X(net202));
 sg13g2_buf_8 fanout203 (.A(net330),
    .X(net203));
 sg13g2_buf_8 fanout204 (.A(net205),
    .X(net204));
 sg13g2_buf_8 fanout205 (.A(net327),
    .X(net205));
 sg13g2_buf_8 fanout206 (.A(net333),
    .X(net206));
 sg13g2_buf_8 fanout207 (.A(\u_lf.kp_sel_latched[0] ),
    .X(net207));
 sg13g2_buf_8 fanout208 (.A(net209),
    .X(net208));
 sg13g2_buf_8 fanout209 (.A(net233),
    .X(net209));
 sg13g2_buf_8 fanout210 (.A(net211),
    .X(net210));
 sg13g2_buf_8 fanout211 (.A(net233),
    .X(net211));
 sg13g2_buf_8 fanout212 (.A(net213),
    .X(net212));
 sg13g2_buf_8 fanout213 (.A(net219),
    .X(net213));
 sg13g2_buf_8 fanout214 (.A(net216),
    .X(net214));
 sg13g2_buf_1 fanout215 (.A(net216),
    .X(net215));
 sg13g2_buf_8 fanout216 (.A(net219),
    .X(net216));
 sg13g2_buf_8 fanout217 (.A(net219),
    .X(net217));
 sg13g2_buf_8 fanout218 (.A(net219),
    .X(net218));
 sg13g2_buf_8 fanout219 (.A(net233),
    .X(net219));
 sg13g2_buf_8 fanout220 (.A(net225),
    .X(net220));
 sg13g2_buf_8 fanout221 (.A(net224),
    .X(net221));
 sg13g2_buf_8 fanout222 (.A(net224),
    .X(net222));
 sg13g2_buf_8 fanout223 (.A(net224),
    .X(net223));
 sg13g2_buf_8 fanout224 (.A(net225),
    .X(net224));
 sg13g2_buf_8 fanout225 (.A(net233),
    .X(net225));
 sg13g2_buf_8 fanout226 (.A(net232),
    .X(net226));
 sg13g2_buf_8 fanout227 (.A(net228),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(net232),
    .X(net228));
 sg13g2_buf_8 fanout229 (.A(net231),
    .X(net229));
 sg13g2_buf_1 fanout230 (.A(net231),
    .X(net230));
 sg13g2_buf_8 fanout231 (.A(net232),
    .X(net231));
 sg13g2_buf_8 fanout232 (.A(net233),
    .X(net232));
 sg13g2_buf_8 fanout233 (.A(rst_n),
    .X(net233));
 sg13g2_buf_8 fanout234 (.A(net236),
    .X(net234));
 sg13g2_buf_1 fanout235 (.A(net236),
    .X(net235));
 sg13g2_buf_8 fanout236 (.A(ena),
    .X(net236));
 sg13g2_buf_8 fanout237 (.A(net238),
    .X(net237));
 sg13g2_buf_1 fanout238 (.A(ena),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(net242),
    .X(net239));
 sg13g2_buf_8 fanout240 (.A(net242),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(net242),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(ena),
    .X(net242));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_tielo tt_um_arthfink_ddmtd_8 (.L_LO(net8));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u_core.fb_sync[0] ),
    .X(net24));
 sg13g2_dlygate4sd3_1 hold2 (.A(\u_core.ref_sync[0] ),
    .X(net25));
 sg13g2_dlygate4sd3_1 hold3 (.A(clk_helper),
    .X(net26));
 sg13g2_dlygate4sd3_1 hold4 (.A(\nco_phase_acc[20] ),
    .X(net27));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0290_),
    .X(net28));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0023_),
    .X(net29));
 sg13g2_dlygate4sd3_1 hold7 (.A(\nco_phase_acc[22] ),
    .X(net30));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0025_),
    .X(net31));
 sg13g2_dlygate4sd3_1 hold9 (.A(\nco_phase_acc[0] ),
    .X(net32));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0003_),
    .X(net33));
 sg13g2_dlygate4sd3_1 hold11 (.A(\u_core.ref_sync[1] ),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0151_),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0141_),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold14 (.A(\nco_phase_acc[18] ),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0288_),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0021_),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold17 (.A(\nco_phase_acc[17] ),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0020_),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold19 (.A(\nco_phase_acc[19] ),
    .X(net42));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0022_),
    .X(net43));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u_core.beat_cnt[7] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold22 (.A(_0086_),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u_core.beat_cnt[4] ),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0083_),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold25 (.A(\u_core.beat_cnt[8] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0087_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u_core.beat_cnt[15] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0094_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u_lf.i_acc[0] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0029_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u_core.beat_cnt[13] ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold32 (.A(_0092_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u_core.fb_samp_d ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0142_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u_core.beat_cnt[10] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0089_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u_core.beat_cnt[0] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0079_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u_core.beat_cnt[9] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0088_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u_core.beat_cnt[5] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0084_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u_core.beat_cnt[12] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0091_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u_core.fb_sync[1] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0124_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold47 (.A(\nco_phase_acc[21] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u_core.beat_cnt[2] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0081_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold50 (.A(\nco_phase_acc[15] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0018_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u_core.beat_cnt[6] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0630_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ctrl[12] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0063_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold56 (.A(\nco_phase_acc[2] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0005_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold58 (.A(\phase_err_beat[3] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0095_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold60 (.A(\nco_phase_acc[10] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0013_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold62 (.A(\nco_phase_acc[16] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0283_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold64 (.A(\ctrl[8] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0059_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold66 (.A(\u_core.beat_cnt[1] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold67 (.A(\nco_phase_acc[14] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0017_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold69 (.A(\nco_phase_acc[12] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0015_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold71 (.A(\nco_phase_acc[4] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0007_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ctrl[19] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0070_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold75 (.A(\u_core.beat_cnt[14] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0640_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold77 (.A(\nco_phase_acc[3] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0006_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold79 (.A(\nco_phase_acc[7] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0010_),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold81 (.A(\u_core.beat_cnt[11] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0637_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold83 (.A(\u_lf.i_acc[29] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0058_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold85 (.A(\u_core.t_ref[4] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0144_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold87 (.A(\nco_phase_acc[6] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0009_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold89 (.A(\u_lf.i_acc[18] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold90 (.A(ref_samp),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0078_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold92 (.A(\ctrl[20] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0071_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold94 (.A(\nco_phase_acc[5] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0008_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold96 (.A(\u_core.t_ref[0] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold97 (.A(\u_core.t_fb[0] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold98 (.A(\nco_phase_acc[1] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0004_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold100 (.A(\ctrl[10] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0061_),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold102 (.A(\u_lf.i_acc[16] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0045_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold104 (.A(\ctrl[11] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0062_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold106 (.A(\ctrl[9] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0060_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold108 (.A(\u_core.t_ref[7] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold109 (.A(_0146_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold110 (.A(\nco_phase_acc[11] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0014_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold112 (.A(\ctrl[15] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold113 (.A(_0066_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold114 (.A(\u_core.t_fb[4] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold115 (.A(\ctrl[13] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0064_),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold117 (.A(\u_lf.i_acc[19] ),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold118 (.A(\u_lf.i_acc[21] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0050_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold120 (.A(\u_core.t_ref[15] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold121 (.A(\nco_phase_acc[13] ),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0016_),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold123 (.A(\u_lf.i_acc[28] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold124 (.A(\u_lf.i_acc[25] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0054_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold126 (.A(\ctrl[23] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold127 (.A(\u_core.t_ref[9] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0117_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold129 (.A(\ctrl[22] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold130 (.A(\u_lf.i_acc[2] ),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0031_),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold132 (.A(\u_core.t_fb[9] ),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0134_),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold134 (.A(\u_lf.i_acc[23] ),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0052_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold136 (.A(\u_core.t_fb[11] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold137 (.A(\u_lf.i_acc[17] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0046_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold139 (.A(\u_core.t_fb[7] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold140 (.A(\u_lf.i_acc[13] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold141 (.A(_0042_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold142 (.A(\phase_err_beat[4] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold143 (.A(\phase_err_beat[8] ),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold144 (.A(_0100_),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold145 (.A(\u_lf.i_acc[7] ),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold146 (.A(_0036_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold147 (.A(\u_core.t_fb[15] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold148 (.A(\nco_phase_acc[9] ),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0012_),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold150 (.A(\u_lf.i_acc[27] ),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0056_),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold152 (.A(\u_core.t_fb[13] ),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold153 (.A(\u_lf.i_acc[20] ),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold154 (.A(\u_core.t_ref[2] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold155 (.A(\u_core.t_ref[11] ),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold156 (.A(\u_core.t_fb[2] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold157 (.A(\ctrl[18] ),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold158 (.A(\u_core.have_ref ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0152_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold160 (.A(\u_lf.i_acc[10] ),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0362_),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0039_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold163 (.A(\u_lf.i_acc[15] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0044_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ctrl[14] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0065_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold167 (.A(\u_lf.i_acc[26] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold168 (.A(phase_valid),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold169 (.A(\u_lf.i_acc[14] ),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold170 (.A(\u_lf.i_acc[24] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0053_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold172 (.A(\u_lf.i_acc[6] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold173 (.A(_0035_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold174 (.A(\u_core.t_ref[14] ),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold175 (.A(\u_lf.i_acc[3] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold176 (.A(\u_lf.i_acc[8] ),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold177 (.A(\u_core.t_ref[5] ),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0113_),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold179 (.A(\u_lf.i_acc[4] ),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold180 (.A(\u_core.t_ref[6] ),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold181 (.A(\u_core.t_ref[13] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold182 (.A(\phase_err_beat[5] ),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0097_),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold184 (.A(\nco_phase_acc[8] ),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold185 (.A(_0011_),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold186 (.A(\u_core.t_fb[6] ),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold187 (.A(\u_core.t_ref[3] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0111_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold189 (.A(\u_core.t_ref[8] ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold190 (.A(\u_core.t_fb[5] ),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold191 (.A(\u_core.t_fb[12] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold192 (.A(_0137_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold193 (.A(\u_lf.i_acc[22] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold194 (.A(\u_core.t_fb[1] ),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold195 (.A(\u_lf.i_acc[1] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold196 (.A(\u_core.t_ref[10] ),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold197 (.A(\u_core.have_fb ),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold198 (.A(_0622_),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold199 (.A(\u_core.t_fb[14] ),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0139_),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold201 (.A(\u_core.t_ref[1] ),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold202 (.A(\u_lf.i_acc[11] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold203 (.A(\u_lf.i_acc[5] ),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold204 (.A(\phase_err_beat[7] ),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold205 (.A(\u_core.t_fb[3] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold206 (.A(_0128_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold207 (.A(\u_core.t_fb[10] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold208 (.A(\u_core.t_fb[8] ),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold209 (.A(\u_lf.i_acc[9] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold210 (.A(\phase_err_beat[9] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold211 (.A(\u_core.t_ref[12] ),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0120_),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold213 (.A(\ctrl[21] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold214 (.A(\phase_err_beat[6] ),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold215 (.A(\ctrl[16] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0002_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold217 (.A(\phase_err_beat[10] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0102_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold219 (.A(\phase_err_beat[13] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0105_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold221 (.A(\ctrl[17] ),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold222 (.A(\u_lf.i_acc[12] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold223 (.A(\u_core.beat_cnt[3] ),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0001_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold225 (.A(\phase_err_beat[15] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold226 (.A(\u_lf.ki_sel_latched[0] ),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold227 (.A(\phase_err_beat[11] ),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold228 (.A(\phase_err_beat[14] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold229 (.A(\phase_err_beat[12] ),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold230 (.A(\u_lf.kp_sel_latched[0] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold231 (.A(\u_core.beat_cnt[11] ),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold232 (.A(\u_lf.i_acc[27] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0483_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold234 (.A(\u_lf.i_acc[16] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold235 (.A(\u_lf.i_acc[16] ),
    .X(net338));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_fill_1 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_194 ();
 sg13g2_decap_8 FILLER_0_201 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_4 FILLER_0_291 ();
 sg13g2_fill_2 FILLER_0_295 ();
 sg13g2_fill_2 FILLER_0_345 ();
 sg13g2_fill_1 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_352 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_4 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_201 ();
 sg13g2_fill_2 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_239 ();
 sg13g2_decap_8 FILLER_1_246 ();
 sg13g2_decap_8 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_decap_8 FILLER_1_267 ();
 sg13g2_decap_8 FILLER_1_274 ();
 sg13g2_decap_8 FILLER_1_281 ();
 sg13g2_fill_2 FILLER_1_288 ();
 sg13g2_fill_2 FILLER_1_329 ();
 sg13g2_fill_1 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_363 ();
 sg13g2_decap_8 FILLER_1_370 ();
 sg13g2_decap_8 FILLER_1_377 ();
 sg13g2_decap_8 FILLER_1_384 ();
 sg13g2_decap_8 FILLER_1_391 ();
 sg13g2_decap_8 FILLER_1_398 ();
 sg13g2_decap_4 FILLER_1_405 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_4 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_193 ();
 sg13g2_fill_1 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_2_239 ();
 sg13g2_decap_8 FILLER_2_246 ();
 sg13g2_decap_8 FILLER_2_253 ();
 sg13g2_decap_4 FILLER_2_260 ();
 sg13g2_fill_2 FILLER_2_268 ();
 sg13g2_fill_1 FILLER_2_297 ();
 sg13g2_fill_2 FILLER_2_334 ();
 sg13g2_fill_1 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_376 ();
 sg13g2_decap_8 FILLER_2_383 ();
 sg13g2_decap_8 FILLER_2_390 ();
 sg13g2_decap_8 FILLER_2_397 ();
 sg13g2_decap_4 FILLER_2_404 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_4 FILLER_3_154 ();
 sg13g2_fill_2 FILLER_3_204 ();
 sg13g2_fill_1 FILLER_3_206 ();
 sg13g2_decap_8 FILLER_3_246 ();
 sg13g2_decap_4 FILLER_3_253 ();
 sg13g2_fill_2 FILLER_3_261 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_decap_4 FILLER_3_380 ();
 sg13g2_decap_8 FILLER_3_393 ();
 sg13g2_decap_8 FILLER_3_400 ();
 sg13g2_fill_2 FILLER_3_407 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_4 FILLER_4_140 ();
 sg13g2_fill_2 FILLER_4_144 ();
 sg13g2_decap_4 FILLER_4_155 ();
 sg13g2_fill_2 FILLER_4_159 ();
 sg13g2_decap_8 FILLER_4_199 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_4 FILLER_4_403 ();
 sg13g2_fill_2 FILLER_4_407 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_fill_1 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_122 ();
 sg13g2_fill_2 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_131 ();
 sg13g2_decap_4 FILLER_5_159 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_fill_1 FILLER_5_203 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_fill_2 FILLER_5_237 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_fill_1 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_4 FILLER_6_91 ();
 sg13g2_fill_2 FILLER_6_108 ();
 sg13g2_fill_1 FILLER_6_110 ();
 sg13g2_decap_8 FILLER_6_124 ();
 sg13g2_fill_1 FILLER_6_131 ();
 sg13g2_fill_2 FILLER_6_168 ();
 sg13g2_fill_2 FILLER_6_181 ();
 sg13g2_fill_1 FILLER_6_183 ();
 sg13g2_fill_2 FILLER_6_194 ();
 sg13g2_fill_1 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_205 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_276 ();
 sg13g2_fill_2 FILLER_6_314 ();
 sg13g2_fill_1 FILLER_6_316 ();
 sg13g2_fill_1 FILLER_6_331 ();
 sg13g2_fill_2 FILLER_6_354 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_4 FILLER_7_84 ();
 sg13g2_fill_2 FILLER_7_88 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_fill_1 FILLER_7_136 ();
 sg13g2_fill_1 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_184 ();
 sg13g2_decap_8 FILLER_7_191 ();
 sg13g2_decap_8 FILLER_7_198 ();
 sg13g2_fill_1 FILLER_7_205 ();
 sg13g2_fill_1 FILLER_7_256 ();
 sg13g2_fill_2 FILLER_7_261 ();
 sg13g2_fill_1 FILLER_7_263 ();
 sg13g2_fill_2 FILLER_7_283 ();
 sg13g2_fill_1 FILLER_7_330 ();
 sg13g2_fill_2 FILLER_7_358 ();
 sg13g2_decap_4 FILLER_7_403 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_4 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_88 ();
 sg13g2_fill_2 FILLER_8_131 ();
 sg13g2_decap_8 FILLER_8_184 ();
 sg13g2_decap_8 FILLER_8_191 ();
 sg13g2_decap_8 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_243 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_2 FILLER_8_321 ();
 sg13g2_fill_2 FILLER_8_365 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_4 FILLER_9_77 ();
 sg13g2_fill_2 FILLER_9_81 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_fill_1 FILLER_9_162 ();
 sg13g2_fill_2 FILLER_9_181 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_fill_2 FILLER_9_203 ();
 sg13g2_fill_1 FILLER_9_247 ();
 sg13g2_decap_8 FILLER_9_253 ();
 sg13g2_decap_8 FILLER_9_260 ();
 sg13g2_decap_8 FILLER_9_271 ();
 sg13g2_decap_8 FILLER_9_278 ();
 sg13g2_decap_8 FILLER_9_285 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_fill_2 FILLER_9_312 ();
 sg13g2_fill_1 FILLER_9_314 ();
 sg13g2_fill_1 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_4 FILLER_10_84 ();
 sg13g2_fill_1 FILLER_10_88 ();
 sg13g2_fill_2 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_164 ();
 sg13g2_decap_8 FILLER_10_183 ();
 sg13g2_decap_8 FILLER_10_190 ();
 sg13g2_fill_2 FILLER_10_197 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_1 FILLER_10_228 ();
 sg13g2_fill_2 FILLER_10_242 ();
 sg13g2_fill_1 FILLER_10_244 ();
 sg13g2_fill_2 FILLER_10_252 ();
 sg13g2_fill_2 FILLER_10_267 ();
 sg13g2_fill_1 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_fill_1 FILLER_10_284 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_317 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_fill_2 FILLER_10_342 ();
 sg13g2_fill_2 FILLER_10_357 ();
 sg13g2_fill_1 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_4 FILLER_11_177 ();
 sg13g2_fill_2 FILLER_11_181 ();
 sg13g2_fill_1 FILLER_11_194 ();
 sg13g2_fill_1 FILLER_11_213 ();
 sg13g2_decap_8 FILLER_11_230 ();
 sg13g2_fill_2 FILLER_11_237 ();
 sg13g2_fill_2 FILLER_11_253 ();
 sg13g2_decap_4 FILLER_11_297 ();
 sg13g2_fill_1 FILLER_11_363 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_fill_2 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_fill_1 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_fill_2 FILLER_12_196 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_12_231 ();
 sg13g2_fill_2 FILLER_12_270 ();
 sg13g2_fill_1 FILLER_12_290 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_2 FILLER_12_346 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_91 ();
 sg13g2_fill_2 FILLER_13_128 ();
 sg13g2_fill_1 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_181 ();
 sg13g2_decap_8 FILLER_13_188 ();
 sg13g2_decap_4 FILLER_13_195 ();
 sg13g2_fill_2 FILLER_13_199 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_302 ();
 sg13g2_fill_2 FILLER_13_331 ();
 sg13g2_fill_2 FILLER_13_342 ();
 sg13g2_fill_2 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_4 FILLER_14_91 ();
 sg13g2_fill_1 FILLER_14_145 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_fill_1 FILLER_14_240 ();
 sg13g2_decap_4 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_fill_1 FILLER_14_350 ();
 sg13g2_fill_2 FILLER_14_356 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_23 ();
 sg13g2_fill_1 FILLER_15_30 ();
 sg13g2_decap_8 FILLER_15_40 ();
 sg13g2_decap_8 FILLER_15_47 ();
 sg13g2_decap_8 FILLER_15_54 ();
 sg13g2_fill_2 FILLER_15_61 ();
 sg13g2_fill_1 FILLER_15_63 ();
 sg13g2_decap_4 FILLER_15_73 ();
 sg13g2_decap_8 FILLER_15_86 ();
 sg13g2_decap_8 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_100 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_4 FILLER_15_137 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_fill_2 FILLER_15_146 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_fill_1 FILLER_15_176 ();
 sg13g2_fill_2 FILLER_15_186 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_fill_2 FILLER_15_217 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_2 FILLER_15_347 ();
 sg13g2_fill_1 FILLER_15_366 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_fill_2 FILLER_16_43 ();
 sg13g2_fill_1 FILLER_16_45 ();
 sg13g2_decap_8 FILLER_16_73 ();
 sg13g2_fill_1 FILLER_16_80 ();
 sg13g2_decap_8 FILLER_16_118 ();
 sg13g2_decap_4 FILLER_16_125 ();
 sg13g2_fill_1 FILLER_16_129 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_fill_2 FILLER_16_180 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_197 ();
 sg13g2_fill_2 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_290 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_fill_2 FILLER_16_305 ();
 sg13g2_fill_2 FILLER_16_349 ();
 sg13g2_fill_1 FILLER_16_351 ();
 sg13g2_fill_1 FILLER_16_360 ();
 sg13g2_decap_8 FILLER_16_401 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_4 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_4 ();
 sg13g2_fill_1 FILLER_17_61 ();
 sg13g2_decap_8 FILLER_17_152 ();
 sg13g2_decap_4 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_decap_4 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_213 ();
 sg13g2_fill_1 FILLER_17_217 ();
 sg13g2_fill_1 FILLER_17_222 ();
 sg13g2_decap_8 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_239 ();
 sg13g2_fill_2 FILLER_17_273 ();
 sg13g2_decap_4 FILLER_17_283 ();
 sg13g2_fill_2 FILLER_17_287 ();
 sg13g2_fill_2 FILLER_17_293 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_361 ();
 sg13g2_fill_1 FILLER_17_370 ();
 sg13g2_fill_2 FILLER_17_389 ();
 sg13g2_fill_1 FILLER_17_391 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_fill_2 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_129 ();
 sg13g2_decap_8 FILLER_18_146 ();
 sg13g2_fill_1 FILLER_18_153 ();
 sg13g2_decap_4 FILLER_18_187 ();
 sg13g2_decap_4 FILLER_18_204 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_4 FILLER_18_228 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_1 FILLER_18_292 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_4 FILLER_18_403 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_29 ();
 sg13g2_fill_2 FILLER_19_58 ();
 sg13g2_fill_2 FILLER_19_73 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_156 ();
 sg13g2_fill_2 FILLER_19_163 ();
 sg13g2_decap_4 FILLER_19_188 ();
 sg13g2_decap_8 FILLER_19_219 ();
 sg13g2_decap_4 FILLER_19_226 ();
 sg13g2_fill_1 FILLER_19_230 ();
 sg13g2_fill_2 FILLER_19_272 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_283 ();
 sg13g2_fill_2 FILLER_19_290 ();
 sg13g2_fill_1 FILLER_19_309 ();
 sg13g2_fill_1 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_22 ();
 sg13g2_fill_1 FILLER_20_36 ();
 sg13g2_fill_1 FILLER_20_51 ();
 sg13g2_decap_4 FILLER_20_79 ();
 sg13g2_decap_4 FILLER_20_96 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_decap_4 FILLER_20_162 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_fill_1 FILLER_20_223 ();
 sg13g2_decap_4 FILLER_20_233 ();
 sg13g2_fill_2 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_292 ();
 sg13g2_fill_2 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_337 ();
 sg13g2_fill_1 FILLER_20_339 ();
 sg13g2_fill_1 FILLER_20_390 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_4 ();
 sg13g2_fill_2 FILLER_21_59 ();
 sg13g2_fill_2 FILLER_21_88 ();
 sg13g2_fill_1 FILLER_21_90 ();
 sg13g2_fill_2 FILLER_21_168 ();
 sg13g2_fill_1 FILLER_21_170 ();
 sg13g2_decap_8 FILLER_21_174 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_fill_1 FILLER_21_183 ();
 sg13g2_fill_1 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_233 ();
 sg13g2_decap_8 FILLER_21_240 ();
 sg13g2_decap_4 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_282 ();
 sg13g2_fill_1 FILLER_21_307 ();
 sg13g2_fill_2 FILLER_21_340 ();
 sg13g2_fill_2 FILLER_21_357 ();
 sg13g2_fill_1 FILLER_21_404 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_4 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_191 ();
 sg13g2_fill_2 FILLER_22_205 ();
 sg13g2_fill_1 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_240 ();
 sg13g2_fill_1 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_267 ();
 sg13g2_decap_4 FILLER_22_292 ();
 sg13g2_fill_2 FILLER_22_296 ();
 sg13g2_fill_2 FILLER_22_317 ();
 sg13g2_fill_1 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_4 FILLER_22_335 ();
 sg13g2_fill_1 FILLER_22_339 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_fill_2 FILLER_23_122 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_decap_4 FILLER_23_184 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_decap_8 FILLER_23_222 ();
 sg13g2_fill_2 FILLER_23_229 ();
 sg13g2_fill_1 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_269 ();
 sg13g2_fill_2 FILLER_23_286 ();
 sg13g2_decap_4 FILLER_23_301 ();
 sg13g2_fill_2 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_328 ();
 sg13g2_decap_8 FILLER_23_335 ();
 sg13g2_fill_1 FILLER_23_342 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_24_87 ();
 sg13g2_fill_2 FILLER_24_107 ();
 sg13g2_fill_1 FILLER_24_109 ();
 sg13g2_fill_2 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_321 ();
 sg13g2_decap_4 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_49 ();
 sg13g2_fill_1 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_2 FILLER_25_190 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_fill_2 FILLER_25_246 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_313 ();
 sg13g2_decap_4 FILLER_25_320 ();
 sg13g2_fill_1 FILLER_25_324 ();
 sg13g2_fill_1 FILLER_25_330 ();
 sg13g2_fill_2 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_389 ();
 sg13g2_fill_1 FILLER_25_391 ();
 sg13g2_fill_1 FILLER_26_68 ();
 sg13g2_fill_1 FILLER_26_157 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_208 ();
 sg13g2_decap_4 FILLER_26_232 ();
 sg13g2_decap_8 FILLER_26_239 ();
 sg13g2_decap_8 FILLER_26_246 ();
 sg13g2_fill_2 FILLER_26_253 ();
 sg13g2_fill_2 FILLER_26_268 ();
 sg13g2_fill_2 FILLER_26_289 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_296 ();
 sg13g2_decap_8 FILLER_26_303 ();
 sg13g2_decap_8 FILLER_26_310 ();
 sg13g2_fill_2 FILLER_26_317 ();
 sg13g2_fill_1 FILLER_26_319 ();
 sg13g2_fill_2 FILLER_26_329 ();
 sg13g2_fill_2 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_131 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_4 FILLER_27_210 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_decap_4 FILLER_27_220 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_247 ();
 sg13g2_fill_1 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_306 ();
 sg13g2_fill_2 FILLER_27_313 ();
 sg13g2_fill_1 FILLER_27_315 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_2 FILLER_27_357 ();
 sg13g2_fill_1 FILLER_27_399 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_37 ();
 sg13g2_fill_1 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_82 ();
 sg13g2_decap_8 FILLER_28_139 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_153 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_fill_1 FILLER_28_229 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_decap_4 FILLER_28_312 ();
 sg13g2_fill_2 FILLER_28_316 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_fill_2 FILLER_28_344 ();
 sg13g2_fill_1 FILLER_28_346 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_4 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_4 ();
 sg13g2_fill_2 FILLER_29_13 ();
 sg13g2_fill_1 FILLER_29_57 ();
 sg13g2_fill_1 FILLER_29_109 ();
 sg13g2_fill_2 FILLER_29_134 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_decap_8 FILLER_29_146 ();
 sg13g2_decap_8 FILLER_29_153 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_215 ();
 sg13g2_decap_4 FILLER_29_226 ();
 sg13g2_decap_4 FILLER_29_251 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_fill_1 FILLER_29_314 ();
 sg13g2_fill_1 FILLER_29_335 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_fill_1 FILLER_29_351 ();
 sg13g2_fill_2 FILLER_29_365 ();
 sg13g2_fill_1 FILLER_29_376 ();
 sg13g2_decap_4 FILLER_30_53 ();
 sg13g2_fill_1 FILLER_30_57 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_4 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_273 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_1 FILLER_30_372 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_35 ();
 sg13g2_decap_4 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_152 ();
 sg13g2_decap_4 FILLER_31_159 ();
 sg13g2_fill_1 FILLER_31_163 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_4 FILLER_31_217 ();
 sg13g2_fill_2 FILLER_31_221 ();
 sg13g2_decap_8 FILLER_31_244 ();
 sg13g2_decap_8 FILLER_31_251 ();
 sg13g2_decap_8 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_368 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_2 FILLER_32_54 ();
 sg13g2_decap_4 FILLER_32_156 ();
 sg13g2_fill_1 FILLER_32_160 ();
 sg13g2_decap_8 FILLER_32_206 ();
 sg13g2_decap_8 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_decap_8 FILLER_32_243 ();
 sg13g2_fill_1 FILLER_32_250 ();
 sg13g2_decap_4 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_353 ();
 sg13g2_fill_1 FILLER_32_399 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_59 ();
 sg13g2_fill_2 FILLER_33_100 ();
 sg13g2_fill_1 FILLER_33_148 ();
 sg13g2_fill_2 FILLER_33_162 ();
 sg13g2_fill_1 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_241 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_fill_1 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_266 ();
 sg13g2_fill_2 FILLER_33_311 ();
 sg13g2_fill_1 FILLER_33_313 ();
 sg13g2_fill_1 FILLER_33_351 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_46 ();
 sg13g2_fill_2 FILLER_34_111 ();
 sg13g2_fill_2 FILLER_34_153 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_216 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_fill_2 FILLER_34_299 ();
 sg13g2_fill_1 FILLER_34_301 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_220 ();
 sg13g2_decap_8 FILLER_35_227 ();
 sg13g2_decap_4 FILLER_35_234 ();
 sg13g2_fill_2 FILLER_35_274 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_2 FILLER_35_332 ();
 sg13g2_fill_2 FILLER_35_347 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_4 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_159 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_decap_4 FILLER_36_235 ();
 sg13g2_fill_2 FILLER_36_239 ();
 sg13g2_fill_1 FILLER_36_268 ();
 sg13g2_decap_8 FILLER_36_309 ();
 sg13g2_decap_8 FILLER_36_316 ();
 sg13g2_decap_4 FILLER_36_323 ();
 sg13g2_fill_2 FILLER_36_362 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_97 ();
 sg13g2_fill_2 FILLER_37_143 ();
 sg13g2_fill_2 FILLER_37_167 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_decap_4 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_1 FILLER_37_266 ();
 sg13g2_fill_2 FILLER_37_280 ();
 sg13g2_fill_1 FILLER_37_373 ();
 sg13g2_decap_4 FILLER_37_383 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_397 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_7 ();
 sg13g2_fill_1 FILLER_38_47 ();
 sg13g2_fill_2 FILLER_38_108 ();
 sg13g2_fill_1 FILLER_38_110 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_fill_2 FILLER_38_184 ();
 sg13g2_fill_1 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_decap_4 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_260 ();
 sg13g2_decap_8 FILLER_38_269 ();
 sg13g2_fill_2 FILLER_38_276 ();
 sg13g2_fill_1 FILLER_38_282 ();
 sg13g2_decap_4 FILLER_38_302 ();
 sg13g2_fill_2 FILLER_38_306 ();
 sg13g2_fill_2 FILLER_38_335 ();
 sg13g2_fill_2 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_fill_1 FILLER_38_370 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
endmodule
