module tt_um_mo_module (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net1;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;

 sg13g2_inv_1 _153_ (.Y(_101_),
    .A(net51));
 sg13g2_inv_1 _154_ (.Y(_102_),
    .A(net56));
 sg13g2_inv_1 _155_ (.Y(_103_),
    .A(net68));
 sg13g2_inv_1 _156_ (.Y(_104_),
    .A(\hvsync_gen.vpos[5] ));
 sg13g2_inv_2 _157_ (.Y(_105_),
    .A(net58));
 sg13g2_inv_1 _158_ (.Y(_106_),
    .A(net78));
 sg13g2_inv_1 _159_ (.Y(_107_),
    .A(\hvsync_gen.hpos[3] ));
 sg13g2_inv_1 _160_ (.Y(_108_),
    .A(\counter[3] ));
 sg13g2_inv_1 _161_ (.Y(_002_),
    .A(\counter[0] ));
 sg13g2_nand4_1 _162_ (.B(net56),
    .C(\hvsync_gen.vpos[6] ),
    .A(net49),
    .Y(_109_),
    .D(\hvsync_gen.vpos[5] ));
 sg13g2_nand2b_1 _163_ (.Y(_110_),
    .B(net53),
    .A_N(\hvsync_gen.vpos[4] ));
 sg13g2_nand3_1 _164_ (.B(_101_),
    .C(_105_),
    .A(net66),
    .Y(_111_));
 sg13g2_nor3_1 _165_ (.A(_109_),
    .B(_110_),
    .C(_111_),
    .Y(_001_));
 sg13g2_and3_1 _166_ (.X(_112_),
    .A(\hvsync_gen.hpos[6] ),
    .B(net13),
    .C(\hvsync_gen.hpos[4] ));
 sg13g2_nand2_1 _167_ (.Y(_113_),
    .A(\hvsync_gen.hpos[7] ),
    .B(\hvsync_gen.hpos[9] ));
 sg13g2_nor3_1 _168_ (.A(\hvsync_gen.hpos[6] ),
    .B(net13),
    .C(\hvsync_gen.hpos[4] ),
    .Y(_114_));
 sg13g2_nor4_1 _169_ (.A(net45),
    .B(_112_),
    .C(_113_),
    .D(_114_),
    .Y(_000_));
 sg13g2_nor2_1 _170_ (.A(\hvsync_gen.hpos[5] ),
    .B(\counter[5] ),
    .Y(_115_));
 sg13g2_nand2_1 _171_ (.Y(_116_),
    .A(\hvsync_gen.hpos[5] ),
    .B(\counter[5] ));
 sg13g2_xnor2_1 _172_ (.Y(_117_),
    .A(net13),
    .B(\counter[5] ));
 sg13g2_nand2_1 _173_ (.Y(_118_),
    .A(\hvsync_gen.hpos[4] ),
    .B(\counter[4] ));
 sg13g2_or2_1 _174_ (.X(_119_),
    .B(\counter[4] ),
    .A(\hvsync_gen.hpos[4] ));
 sg13g2_a22oi_1 _175_ (.Y(_120_),
    .B1(\counter[0] ),
    .B2(\hvsync_gen.hpos[0] ),
    .A2(\counter[1] ),
    .A1(\hvsync_gen.hpos[1] ));
 sg13g2_nor2_1 _176_ (.A(\hvsync_gen.hpos[2] ),
    .B(\counter[2] ),
    .Y(_121_));
 sg13g2_nor2_1 _177_ (.A(\hvsync_gen.hpos[1] ),
    .B(\counter[1] ),
    .Y(_122_));
 sg13g2_or3_1 _178_ (.A(_120_),
    .B(_121_),
    .C(_122_),
    .X(_123_));
 sg13g2_a22oi_1 _179_ (.Y(_124_),
    .B1(\counter[2] ),
    .B2(\hvsync_gen.hpos[2] ),
    .A2(\counter[3] ),
    .A1(\hvsync_gen.hpos[3] ));
 sg13g2_a22oi_1 _180_ (.Y(_125_),
    .B1(_123_),
    .B2(_124_),
    .A2(_108_),
    .A1(_107_));
 sg13g2_nand2_1 _181_ (.Y(_126_),
    .A(_119_),
    .B(_125_));
 sg13g2_a21oi_1 _182_ (.A1(_118_),
    .A2(_126_),
    .Y(_127_),
    .B1(_117_));
 sg13g2_nand2_1 _183_ (.Y(_128_),
    .A(\hvsync_gen.hpos[9] ),
    .B(\hvsync_gen.hpos[8] ));
 sg13g2_nand4_1 _184_ (.B(_109_),
    .C(_113_),
    .A(_105_),
    .Y(_129_),
    .D(_128_));
 sg13g2_and3_1 _185_ (.X(_130_),
    .A(_117_),
    .B(_118_),
    .C(_126_));
 sg13g2_nor3_1 _186_ (.A(_127_),
    .B(_129_),
    .C(_130_),
    .Y(uo_out[0]));
 sg13g2_nor2_2 _187_ (.A(_101_),
    .B(_129_),
    .Y(uo_out[5]));
 sg13g2_nand3b_1 _188_ (.B(_118_),
    .C(_119_),
    .Y(_030_),
    .A_N(_117_));
 sg13g2_a221oi_1 _189_ (.B2(_124_),
    .C1(_030_),
    .B1(_123_),
    .A1(_107_),
    .Y(_031_),
    .A2(_108_));
 sg13g2_o21ai_1 _190_ (.B1(_116_),
    .Y(_032_),
    .A1(_115_),
    .A2(_118_));
 sg13g2_nand2_1 _191_ (.Y(_033_),
    .A(\hvsync_gen.hpos[6] ),
    .B(\counter[6] ));
 sg13g2_xnor2_1 _192_ (.Y(_034_),
    .A(\hvsync_gen.hpos[6] ),
    .B(\counter[6] ));
 sg13g2_inv_1 _193_ (.Y(_035_),
    .A(_034_));
 sg13g2_o21ai_1 _194_ (.B1(_035_),
    .Y(_036_),
    .A1(_031_),
    .A2(_032_));
 sg13g2_nor3_1 _195_ (.A(_031_),
    .B(_032_),
    .C(_035_),
    .Y(_037_));
 sg13g2_nor2_1 _196_ (.A(_129_),
    .B(_037_),
    .Y(_038_));
 sg13g2_and2_1 _197_ (.A(_036_),
    .B(_038_),
    .X(uo_out[1]));
 sg13g2_nor2_1 _198_ (.A(_104_),
    .B(_129_),
    .Y(uo_out[6]));
 sg13g2_xnor2_1 _199_ (.Y(_039_),
    .A(\hvsync_gen.hpos[7] ),
    .B(\counter[7] ));
 sg13g2_a21oi_1 _200_ (.A1(_033_),
    .A2(_036_),
    .Y(_040_),
    .B1(_039_));
 sg13g2_and3_1 _201_ (.X(_041_),
    .A(_033_),
    .B(_036_),
    .C(_039_));
 sg13g2_nor3_1 _202_ (.A(_129_),
    .B(_040_),
    .C(_041_),
    .Y(uo_out[2]));
 sg13g2_xor2_1 _203_ (.B(\counter[0] ),
    .A(\counter[1] ),
    .X(_003_));
 sg13g2_nand3_1 _204_ (.B(\counter[1] ),
    .C(\counter[0] ),
    .A(\counter[2] ),
    .Y(_042_));
 sg13g2_a21o_1 _205_ (.A2(\counter[0] ),
    .A1(\counter[1] ),
    .B1(\counter[2] ),
    .X(_043_));
 sg13g2_and2_1 _206_ (.A(_042_),
    .B(_043_),
    .X(_004_));
 sg13g2_nor2_2 _207_ (.A(_108_),
    .B(_042_),
    .Y(_044_));
 sg13g2_xnor2_1 _208_ (.Y(_005_),
    .A(\counter[3] ),
    .B(_042_));
 sg13g2_xor2_1 _209_ (.B(_044_),
    .A(\counter[4] ),
    .X(_006_));
 sg13g2_nand3_1 _210_ (.B(\counter[4] ),
    .C(_044_),
    .A(\counter[5] ),
    .Y(_045_));
 sg13g2_a21o_1 _211_ (.A2(_044_),
    .A1(\counter[4] ),
    .B1(\counter[5] ),
    .X(_046_));
 sg13g2_and2_1 _212_ (.A(_045_),
    .B(_046_),
    .X(_007_));
 sg13g2_nand4_1 _213_ (.B(\counter[4] ),
    .C(\counter[6] ),
    .A(\counter[5] ),
    .Y(_047_),
    .D(_044_));
 sg13g2_xnor2_1 _214_ (.Y(_008_),
    .A(\counter[6] ),
    .B(_045_));
 sg13g2_xnor2_1 _215_ (.Y(_009_),
    .A(\counter[7] ),
    .B(_047_));
 sg13g2_and2_1 _216_ (.A(net44),
    .B(net63),
    .X(_048_));
 sg13g2_nand4_1 _217_ (.B(net63),
    .C(net60),
    .A(net44),
    .Y(_049_),
    .D(net47));
 sg13g2_nor2_2 _218_ (.A(_106_),
    .B(_049_),
    .Y(_050_));
 sg13g2_nor4_1 _219_ (.A(net79),
    .B(\hvsync_gen.hpos[6] ),
    .C(net13),
    .D(_128_),
    .Y(_051_));
 sg13g2_nand2_1 _220_ (.Y(_052_),
    .A(_050_),
    .B(_051_));
 sg13g2_and2_1 _221_ (.A(net14),
    .B(_052_),
    .X(_053_));
 sg13g2_nand2_2 _222_ (.Y(_054_),
    .A(net14),
    .B(_052_));
 sg13g2_nor2_1 _223_ (.A(net44),
    .B(_054_),
    .Y(_010_));
 sg13g2_nor2_1 _224_ (.A(net44),
    .B(net63),
    .Y(_055_));
 sg13g2_nor3_1 _225_ (.A(_048_),
    .B(_054_),
    .C(_055_),
    .Y(_011_));
 sg13g2_o21ai_1 _226_ (.B1(_053_),
    .Y(_056_),
    .A1(net47),
    .A2(_048_));
 sg13g2_a21oi_1 _227_ (.A1(net47),
    .A2(_048_),
    .Y(_012_),
    .B1(_056_));
 sg13g2_a21oi_1 _228_ (.A1(net47),
    .A2(_048_),
    .Y(_057_),
    .B1(net60));
 sg13g2_nand2_1 _229_ (.Y(_058_),
    .A(net14),
    .B(_049_));
 sg13g2_nor2_1 _230_ (.A(net61),
    .B(_058_),
    .Y(_013_));
 sg13g2_o21ai_1 _231_ (.B1(net14),
    .Y(_059_),
    .A1(_106_),
    .A2(_049_));
 sg13g2_a21oi_1 _232_ (.A1(_106_),
    .A2(_049_),
    .Y(_014_),
    .B1(_059_));
 sg13g2_o21ai_1 _233_ (.B1(_053_),
    .Y(_060_),
    .A1(net13),
    .A2(_050_));
 sg13g2_a21oi_1 _234_ (.A1(net13),
    .A2(_050_),
    .Y(_015_),
    .B1(_060_));
 sg13g2_and3_2 _235_ (.X(_061_),
    .A(net73),
    .B(net13),
    .C(_050_));
 sg13g2_a21oi_1 _236_ (.A1(net13),
    .A2(_050_),
    .Y(_062_),
    .B1(net73));
 sg13g2_nor3_1 _237_ (.A(_054_),
    .B(_061_),
    .C(net74),
    .Y(_016_));
 sg13g2_xnor2_1 _238_ (.Y(_063_),
    .A(net64),
    .B(_061_));
 sg13g2_nor2_1 _239_ (.A(_054_),
    .B(_063_),
    .Y(_017_));
 sg13g2_a21oi_1 _240_ (.A1(net64),
    .A2(_061_),
    .Y(_064_),
    .B1(net45));
 sg13g2_and3_1 _241_ (.X(_065_),
    .A(net64),
    .B(net45),
    .C(_061_));
 sg13g2_nor3_1 _242_ (.A(_054_),
    .B(net65),
    .C(_065_),
    .Y(_018_));
 sg13g2_nor2_1 _243_ (.A(net76),
    .B(_065_),
    .Y(_066_));
 sg13g2_a21oi_1 _244_ (.A1(net76),
    .A2(_065_),
    .Y(_067_),
    .B1(_054_));
 sg13g2_nor2b_1 _245_ (.A(_066_),
    .B_N(_067_),
    .Y(_019_));
 sg13g2_nor3_1 _246_ (.A(\hvsync_gen.vpos[7] ),
    .B(\hvsync_gen.vpos[6] ),
    .C(\hvsync_gen.vpos[5] ),
    .Y(_068_));
 sg13g2_or2_1 _247_ (.X(_069_),
    .B(net55),
    .A(net66));
 sg13g2_nor4_1 _248_ (.A(_101_),
    .B(\hvsync_gen.vpos[8] ),
    .C(_110_),
    .D(_069_),
    .Y(_070_));
 sg13g2_nand3_1 _249_ (.B(_068_),
    .C(_070_),
    .A(net58),
    .Y(_071_));
 sg13g2_nand3_1 _250_ (.B(_050_),
    .C(net80),
    .A(net14),
    .Y(_072_));
 sg13g2_nor2b_2 _251_ (.A(_072_),
    .B_N(_071_),
    .Y(_073_));
 sg13g2_nand2b_2 _252_ (.Y(_074_),
    .B(_071_),
    .A_N(_072_));
 sg13g2_nor2_1 _253_ (.A(net55),
    .B(_073_),
    .Y(_075_));
 sg13g2_a21oi_1 _254_ (.A1(net55),
    .A2(_054_),
    .Y(_020_),
    .B1(_075_));
 sg13g2_a21oi_1 _255_ (.A1(net66),
    .A2(net55),
    .Y(_076_),
    .B1(_072_));
 sg13g2_a21o_1 _256_ (.A2(net11),
    .A1(net66),
    .B1(_076_),
    .X(_077_));
 sg13g2_and2_1 _257_ (.A(_069_),
    .B(_077_),
    .X(_021_));
 sg13g2_nand2_1 _258_ (.Y(_078_),
    .A(net51),
    .B(net11));
 sg13g2_a21oi_1 _259_ (.A1(\hvsync_gen.vpos[1] ),
    .A2(\hvsync_gen.vpos[0] ),
    .Y(_079_),
    .B1(net51));
 sg13g2_nand3_1 _260_ (.B(net51),
    .C(\hvsync_gen.vpos[0] ),
    .A(\hvsync_gen.vpos[1] ),
    .Y(_080_));
 sg13g2_nand2b_1 _261_ (.Y(_081_),
    .B(_080_),
    .A_N(_079_));
 sg13g2_o21ai_1 _262_ (.B1(_078_),
    .Y(_022_),
    .A1(_074_),
    .A2(_081_));
 sg13g2_nand2_1 _263_ (.Y(_082_),
    .A(net53),
    .B(net11));
 sg13g2_and4_1 _264_ (.A(net66),
    .B(net51),
    .C(net53),
    .D(net55),
    .X(_083_));
 sg13g2_xor2_1 _265_ (.B(_080_),
    .A(net53),
    .X(_084_));
 sg13g2_o21ai_1 _266_ (.B1(_082_),
    .Y(_023_),
    .A1(_074_),
    .A2(_084_));
 sg13g2_nand2_1 _267_ (.Y(_085_),
    .A(net72),
    .B(net11));
 sg13g2_xnor2_1 _268_ (.Y(_086_),
    .A(net72),
    .B(_083_));
 sg13g2_o21ai_1 _269_ (.B1(_085_),
    .Y(_024_),
    .A1(_074_),
    .A2(_086_));
 sg13g2_nand2_1 _270_ (.Y(_087_),
    .A(net70),
    .B(net11));
 sg13g2_a21oi_1 _271_ (.A1(\hvsync_gen.vpos[4] ),
    .A2(_083_),
    .Y(_088_),
    .B1(net70));
 sg13g2_nand3_1 _272_ (.B(net70),
    .C(_083_),
    .A(\hvsync_gen.vpos[4] ),
    .Y(_089_));
 sg13g2_nand2b_1 _273_ (.Y(_090_),
    .B(_089_),
    .A_N(_088_));
 sg13g2_o21ai_1 _274_ (.B1(_087_),
    .Y(_025_),
    .A1(_074_),
    .A2(_090_));
 sg13g2_nand2_1 _275_ (.Y(_091_),
    .A(net68),
    .B(net11));
 sg13g2_nand4_1 _276_ (.B(net68),
    .C(\hvsync_gen.vpos[5] ),
    .A(\hvsync_gen.vpos[4] ),
    .Y(_092_),
    .D(_083_));
 sg13g2_nand2_1 _277_ (.Y(_093_),
    .A(_073_),
    .B(_092_));
 sg13g2_a22oi_1 _278_ (.Y(_026_),
    .B1(_091_),
    .B2(_093_),
    .A2(_089_),
    .A1(_103_));
 sg13g2_nand2_1 _279_ (.Y(_094_),
    .A(net56),
    .B(net11));
 sg13g2_nor2_1 _280_ (.A(_102_),
    .B(_092_),
    .Y(_095_));
 sg13g2_xnor2_1 _281_ (.Y(_096_),
    .A(_102_),
    .B(_092_));
 sg13g2_o21ai_1 _282_ (.B1(_094_),
    .Y(_027_),
    .A1(_074_),
    .A2(_096_));
 sg13g2_nand2_1 _283_ (.Y(_097_),
    .A(net49),
    .B(_095_));
 sg13g2_a21oi_1 _284_ (.A1(_073_),
    .A2(_097_),
    .Y(_098_),
    .B1(net11));
 sg13g2_a21oi_1 _285_ (.A1(_073_),
    .A2(_095_),
    .Y(_099_),
    .B1(net49));
 sg13g2_nor2_1 _286_ (.A(_098_),
    .B(net50),
    .Y(_028_));
 sg13g2_nand4_1 _287_ (.B(_105_),
    .C(_073_),
    .A(net49),
    .Y(_100_),
    .D(_095_));
 sg13g2_o21ai_1 _288_ (.B1(_100_),
    .Y(_029_),
    .A1(_105_),
    .A2(_098_));
 sg13g2_dfrbpq_2 _289_ (.RESET_B(net14),
    .D(_002_),
    .Q(\counter[0] ),
    .CLK(net12));
 sg13g2_dfrbpq_2 _290_ (.RESET_B(net15),
    .D(_003_),
    .Q(\counter[1] ),
    .CLK(net12));
 sg13g2_dfrbpq_2 _291_ (.RESET_B(net15),
    .D(_004_),
    .Q(\counter[2] ),
    .CLK(net12));
 sg13g2_dfrbpq_1 _292_ (.RESET_B(net15),
    .D(_005_),
    .Q(\counter[3] ),
    .CLK(net12));
 sg13g2_dfrbpq_2 _293_ (.RESET_B(net15),
    .D(_006_),
    .Q(\counter[4] ),
    .CLK(net12));
 sg13g2_dfrbpq_2 _294_ (.RESET_B(net14),
    .D(_007_),
    .Q(\counter[5] ),
    .CLK(net12));
 sg13g2_dfrbpq_2 _295_ (.RESET_B(net15),
    .D(_008_),
    .Q(\counter[6] ),
    .CLK(\hvsync_gen.vsync ));
 sg13g2_dfrbpq_1 _296_ (.RESET_B(net14),
    .D(_009_),
    .Q(\counter[7] ),
    .CLK(net12));
 sg13g2_dfrbpq_2 _297_ (.RESET_B(net40),
    .D(_010_),
    .Q(\hvsync_gen.hpos[0] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _298_ (.RESET_B(net39),
    .D(_011_),
    .Q(\hvsync_gen.hpos[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _299_ (.RESET_B(net38),
    .D(net48),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_1 _300_ (.RESET_B(net37),
    .D(net62),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _301_ (.RESET_B(net36),
    .D(_014_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _302_ (.RESET_B(net35),
    .D(_015_),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _303_ (.RESET_B(net34),
    .D(net75),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _304_ (.RESET_B(net33),
    .D(_017_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _305_ (.RESET_B(net32),
    .D(_018_),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _306_ (.RESET_B(net43),
    .D(_019_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _307_ (.RESET_B(net31),
    .D(net46),
    .Q(hsync),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _308_ (.RESET_B(net30),
    .D(_020_),
    .Q(\hvsync_gen.vpos[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _309_ (.RESET_B(net28),
    .D(_021_),
    .Q(\hvsync_gen.vpos[1] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _310_ (.RESET_B(net26),
    .D(net52),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _311_ (.RESET_B(net24),
    .D(net54),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _312_ (.RESET_B(net22),
    .D(_024_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _313_ (.RESET_B(net41),
    .D(net71),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _314_ (.RESET_B(net27),
    .D(net69),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _315_ (.RESET_B(net23),
    .D(net57),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _316_ (.RESET_B(net29),
    .D(_028_),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_1 _317_ (.RESET_B(net25),
    .D(net59),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _318_ (.RESET_B(net42),
    .D(net67),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_tiehi _315__18 (.L_HI(net23));
 sg13g2_tiehi _311__19 (.L_HI(net24));
 sg13g2_tiehi _317__20 (.L_HI(net25));
 sg13g2_tiehi _310__21 (.L_HI(net26));
 sg13g2_tiehi _314__22 (.L_HI(net27));
 sg13g2_tiehi _309__23 (.L_HI(net28));
 sg13g2_tiehi _316__24 (.L_HI(net29));
 sg13g2_tiehi _308__25 (.L_HI(net30));
 sg13g2_tiehi _307__26 (.L_HI(net31));
 sg13g2_tiehi _305__27 (.L_HI(net32));
 sg13g2_tiehi _304__28 (.L_HI(net33));
 sg13g2_tiehi _303__29 (.L_HI(net34));
 sg13g2_tiehi _302__30 (.L_HI(net35));
 sg13g2_tiehi _301__31 (.L_HI(net36));
 sg13g2_tiehi _300__32 (.L_HI(net37));
 sg13g2_tiehi _299__33 (.L_HI(net38));
 sg13g2_tiehi _298__34 (.L_HI(net39));
 sg13g2_tiehi _297__35 (.L_HI(net40));
 sg13g2_tiehi _313__36 (.L_HI(net41));
 sg13g2_tiehi _318__37 (.L_HI(net42));
 sg13g2_tiehi _306__38 (.L_HI(net43));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_mo_module_2 (.L_LO(net2));
 sg13g2_tielo tt_um_mo_module_3 (.L_LO(net3));
 sg13g2_tielo tt_um_mo_module_4 (.L_LO(net4));
 sg13g2_tielo tt_um_mo_module_5 (.L_LO(net5));
 sg13g2_tielo tt_um_mo_module_6 (.L_LO(net6));
 sg13g2_tielo tt_um_mo_module_7 (.L_LO(net7));
 sg13g2_tielo tt_um_mo_module_8 (.L_LO(net8));
 sg13g2_tielo tt_um_mo_module_9 (.L_LO(net9));
 sg13g2_tielo tt_um_mo_module_10 (.L_LO(net10));
 sg13g2_tielo tt_um_mo_module_11 (.L_LO(net16));
 sg13g2_tielo tt_um_mo_module_12 (.L_LO(net17));
 sg13g2_tielo tt_um_mo_module_13 (.L_LO(net18));
 sg13g2_tielo tt_um_mo_module_14 (.L_LO(net19));
 sg13g2_tielo tt_um_mo_module_15 (.L_LO(net20));
 sg13g2_tielo tt_um_mo_module_16 (.L_LO(net21));
 sg13g2_tiehi _312__17 (.L_HI(net22));
 sg13g2_buf_1 _357_ (.A(net12),
    .X(uo_out[3]));
 sg13g2_buf_1 _358_ (.A(uo_out[5]),
    .X(uo_out[4]));
 sg13g2_buf_1 _359_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout11 (.A(_053_),
    .X(net11));
 sg13g2_buf_8 fanout12 (.A(\hvsync_gen.vsync ),
    .X(net12));
 sg13g2_buf_8 fanout13 (.A(net77),
    .X(net13));
 sg13g2_buf_8 fanout14 (.A(rst_n),
    .X(net14));
 sg13g2_buf_8 fanout15 (.A(rst_n),
    .X(net15));
 sg13g2_tielo tt_um_mo_module_1 (.L_LO(net1));
 sg13g2_buf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hvsync_gen.hpos[0] ),
    .X(net44));
 sg13g2_dlygate4sd3_1 hold2 (.A(\hvsync_gen.hpos[8] ),
    .X(net45));
 sg13g2_dlygate4sd3_1 hold3 (.A(_000_),
    .X(net46));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.hpos[2] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold5 (.A(_012_),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold6 (.A(\hvsync_gen.vpos[8] ),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold7 (.A(_099_),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold8 (.A(\hvsync_gen.vpos[2] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold9 (.A(_022_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold10 (.A(\hvsync_gen.vpos[3] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold11 (.A(_023_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold12 (.A(\hvsync_gen.vpos[0] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hvsync_gen.vpos[7] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold14 (.A(_027_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hvsync_gen.vpos[9] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold16 (.A(_029_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold17 (.A(\hvsync_gen.hpos[3] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold18 (.A(_057_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold19 (.A(_013_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold20 (.A(\hvsync_gen.hpos[1] ),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hvsync_gen.hpos[7] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold22 (.A(_064_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.vpos[1] ),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold24 (.A(_001_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hvsync_gen.vpos[6] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold26 (.A(_026_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hvsync_gen.vpos[5] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold28 (.A(_025_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hvsync_gen.vpos[4] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hvsync_gen.hpos[6] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold31 (.A(_062_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold32 (.A(_016_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hvsync_gen.hpos[9] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold34 (.A(\hvsync_gen.hpos[5] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold35 (.A(\hvsync_gen.hpos[4] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold36 (.A(\hvsync_gen.hpos[7] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold37 (.A(_051_),
    .X(net80));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_294 ();
 sg13g2_decap_8 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_336 ();
 sg13g2_decap_8 FILLER_22_343 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_decap_8 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_364 ();
 sg13g2_decap_8 FILLER_22_371 ();
 sg13g2_decap_8 FILLER_22_378 ();
 sg13g2_decap_8 FILLER_22_385 ();
 sg13g2_decap_8 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_399 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_8 FILLER_24_168 ();
 sg13g2_decap_8 FILLER_24_175 ();
 sg13g2_decap_8 FILLER_24_182 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_decap_8 FILLER_24_210 ();
 sg13g2_decap_8 FILLER_24_217 ();
 sg13g2_decap_8 FILLER_24_224 ();
 sg13g2_decap_8 FILLER_24_231 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_4 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_296 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_fill_2 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_205 ();
 sg13g2_decap_8 FILLER_25_215 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_decap_4 FILLER_25_229 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_fill_2 FILLER_25_270 ();
 sg13g2_fill_1 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_345 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_decap_8 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_366 ();
 sg13g2_decap_8 FILLER_25_373 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_decap_8 FILLER_25_387 ();
 sg13g2_decap_8 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_189 ();
 sg13g2_decap_4 FILLER_26_222 ();
 sg13g2_fill_2 FILLER_26_231 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_fill_2 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_337 ();
 sg13g2_decap_8 FILLER_26_344 ();
 sg13g2_decap_8 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_358 ();
 sg13g2_decap_8 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_372 ();
 sg13g2_decap_8 FILLER_26_379 ();
 sg13g2_decap_8 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_4 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_123 ();
 sg13g2_decap_4 FILLER_27_153 ();
 sg13g2_decap_8 FILLER_27_183 ();
 sg13g2_decap_8 FILLER_27_190 ();
 sg13g2_decap_4 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_216 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_238 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_fill_1 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_fill_1 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_103 ();
 sg13g2_decap_8 FILLER_28_110 ();
 sg13g2_fill_2 FILLER_28_117 ();
 sg13g2_decap_4 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_146 ();
 sg13g2_fill_2 FILLER_28_189 ();
 sg13g2_fill_1 FILLER_28_191 ();
 sg13g2_fill_1 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_285 ();
 sg13g2_decap_4 FILLER_28_290 ();
 sg13g2_fill_2 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_331 ();
 sg13g2_decap_8 FILLER_28_338 ();
 sg13g2_decap_8 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_352 ();
 sg13g2_decap_8 FILLER_28_359 ();
 sg13g2_decap_8 FILLER_28_366 ();
 sg13g2_decap_8 FILLER_28_373 ();
 sg13g2_decap_8 FILLER_28_380 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_8 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_fill_2 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_decap_4 FILLER_29_134 ();
 sg13g2_fill_1 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_156 ();
 sg13g2_fill_1 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_171 ();
 sg13g2_decap_8 FILLER_29_177 ();
 sg13g2_decap_8 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_4 FILLER_29_205 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_261 ();
 sg13g2_decap_8 FILLER_29_268 ();
 sg13g2_decap_8 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_294 ();
 sg13g2_decap_8 FILLER_29_302 ();
 sg13g2_decap_8 FILLER_29_309 ();
 sg13g2_decap_8 FILLER_29_316 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_decap_8 FILLER_29_337 ();
 sg13g2_decap_8 FILLER_29_344 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_8 FILLER_29_358 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_8 FILLER_29_379 ();
 sg13g2_decap_8 FILLER_29_386 ();
 sg13g2_decap_8 FILLER_29_393 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_97 ();
 sg13g2_decap_8 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_125 ();
 sg13g2_decap_4 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_219 ();
 sg13g2_decap_4 FILLER_30_234 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_decap_8 FILLER_30_300 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_367 ();
 sg13g2_decap_8 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_381 ();
 sg13g2_decap_8 FILLER_30_388 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_4 FILLER_31_84 ();
 sg13g2_fill_1 FILLER_31_116 ();
 sg13g2_fill_2 FILLER_31_123 ();
 sg13g2_fill_1 FILLER_31_135 ();
 sg13g2_decap_8 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_243 ();
 sg13g2_decap_4 FILLER_31_250 ();
 sg13g2_fill_1 FILLER_31_254 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_305 ();
 sg13g2_fill_1 FILLER_31_319 ();
 sg13g2_decap_8 FILLER_31_348 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_362 ();
 sg13g2_decap_8 FILLER_31_369 ();
 sg13g2_decap_8 FILLER_31_376 ();
 sg13g2_decap_8 FILLER_31_383 ();
 sg13g2_decap_8 FILLER_31_390 ();
 sg13g2_decap_8 FILLER_31_397 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_fill_2 FILLER_32_91 ();
 sg13g2_fill_1 FILLER_32_93 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_decap_8 FILLER_32_132 ();
 sg13g2_decap_4 FILLER_32_139 ();
 sg13g2_fill_2 FILLER_32_143 ();
 sg13g2_decap_8 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_183 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_1 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_32_287 ();
 sg13g2_decap_8 FILLER_32_294 ();
 sg13g2_decap_4 FILLER_32_301 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_320 ();
 sg13g2_decap_8 FILLER_32_327 ();
 sg13g2_decap_8 FILLER_32_334 ();
 sg13g2_decap_8 FILLER_32_341 ();
 sg13g2_decap_8 FILLER_32_348 ();
 sg13g2_decap_8 FILLER_32_355 ();
 sg13g2_decap_8 FILLER_32_362 ();
 sg13g2_decap_8 FILLER_32_369 ();
 sg13g2_decap_8 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_383 ();
 sg13g2_decap_8 FILLER_32_390 ();
 sg13g2_decap_8 FILLER_32_397 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_4 FILLER_33_84 ();
 sg13g2_decap_4 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_194 ();
 sg13g2_decap_8 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_208 ();
 sg13g2_fill_1 FILLER_33_230 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_decap_4 FILLER_33_297 ();
 sg13g2_fill_1 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_fill_2 FILLER_34_91 ();
 sg13g2_fill_2 FILLER_34_136 ();
 sg13g2_fill_1 FILLER_34_138 ();
 sg13g2_fill_2 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_fill_1 FILLER_34_191 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_268 ();
 sg13g2_decap_4 FILLER_34_290 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_decap_8 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_343 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_8 FILLER_34_378 ();
 sg13g2_decap_8 FILLER_34_385 ();
 sg13g2_decap_8 FILLER_34_392 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_4 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_122 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_269 ();
 sg13g2_fill_2 FILLER_35_276 ();
 sg13g2_fill_1 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_284 ();
 sg13g2_decap_8 FILLER_35_291 ();
 sg13g2_decap_8 FILLER_35_298 ();
 sg13g2_decap_8 FILLER_35_305 ();
 sg13g2_decap_8 FILLER_35_312 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_361 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_115 ();
 sg13g2_fill_1 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_162 ();
 sg13g2_decap_8 FILLER_36_169 ();
 sg13g2_decap_8 FILLER_36_176 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_decap_8 FILLER_36_190 ();
 sg13g2_fill_2 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_decap_8 FILLER_36_289 ();
 sg13g2_decap_8 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_331 ();
 sg13g2_decap_8 FILLER_36_338 ();
 sg13g2_decap_8 FILLER_36_345 ();
 sg13g2_decap_8 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_366 ();
 sg13g2_decap_8 FILLER_36_373 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_4 FILLER_37_133 ();
 sg13g2_fill_2 FILLER_37_137 ();
 sg13g2_decap_4 FILLER_37_143 ();
 sg13g2_fill_2 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_4 FILLER_37_186 ();
 sg13g2_fill_1 FILLER_37_190 ();
 sg13g2_decap_4 FILLER_37_218 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_263 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_decap_8 FILLER_37_277 ();
 sg13g2_decap_8 FILLER_37_284 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_decap_8 FILLER_37_298 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_fill_2 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_212 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_fill_1 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net1;
 assign uio_oe[1] = net2;
 assign uio_oe[2] = net3;
 assign uio_oe[3] = net4;
 assign uio_oe[4] = net5;
 assign uio_oe[5] = net6;
 assign uio_oe[6] = net7;
 assign uio_oe[7] = net8;
 assign uio_out[0] = net9;
 assign uio_out[1] = net10;
 assign uio_out[2] = net16;
 assign uio_out[3] = net17;
 assign uio_out[4] = net18;
 assign uio_out[5] = net19;
 assign uio_out[6] = net20;
 assign uio_out[7] = net21;
endmodule
