module tt_um_swenson_cqs (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire net56;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire \bp_addr_in[0] ;
 wire \bp_addr_in[10] ;
 wire \bp_addr_in[11] ;
 wire \bp_addr_in[12] ;
 wire \bp_addr_in[13] ;
 wire \bp_addr_in[14] ;
 wire \bp_addr_in[15] ;
 wire \bp_addr_in[16] ;
 wire \bp_addr_in[17] ;
 wire \bp_addr_in[18] ;
 wire \bp_addr_in[19] ;
 wire \bp_addr_in[1] ;
 wire \bp_addr_in[2] ;
 wire \bp_addr_in[3] ;
 wire \bp_addr_in[4] ;
 wire \bp_addr_in[5] ;
 wire \bp_addr_in[6] ;
 wire \bp_addr_in[7] ;
 wire \bp_addr_in[8] ;
 wire \bp_addr_in[9] ;
 wire \bp_addr_out[0] ;
 wire \bp_addr_out[10] ;
 wire \bp_addr_out[11] ;
 wire \bp_addr_out[12] ;
 wire \bp_addr_out[13] ;
 wire \bp_addr_out[14] ;
 wire \bp_addr_out[15] ;
 wire \bp_addr_out[16] ;
 wire \bp_addr_out[17] ;
 wire \bp_addr_out[18] ;
 wire \bp_addr_out[19] ;
 wire \bp_addr_out[1] ;
 wire \bp_addr_out[2] ;
 wire \bp_addr_out[3] ;
 wire \bp_addr_out[4] ;
 wire \bp_addr_out[5] ;
 wire \bp_addr_out[6] ;
 wire \bp_addr_out[7] ;
 wire \bp_addr_out[8] ;
 wire \bp_addr_out[9] ;
 wire \bp_core.addr_reg[0] ;
 wire \bp_core.addr_reg[10] ;
 wire \bp_core.addr_reg[11] ;
 wire \bp_core.addr_reg[12] ;
 wire \bp_core.addr_reg[13] ;
 wire \bp_core.addr_reg[14] ;
 wire \bp_core.addr_reg[15] ;
 wire \bp_core.addr_reg[16] ;
 wire \bp_core.addr_reg[17] ;
 wire \bp_core.addr_reg[18] ;
 wire \bp_core.addr_reg[19] ;
 wire \bp_core.addr_reg[1] ;
 wire \bp_core.addr_reg[2] ;
 wire \bp_core.addr_reg[3] ;
 wire \bp_core.addr_reg[4] ;
 wire \bp_core.addr_reg[5] ;
 wire \bp_core.addr_reg[6] ;
 wire \bp_core.addr_reg[7] ;
 wire \bp_core.addr_reg[8] ;
 wire \bp_core.addr_reg[9] ;
 wire \bp_core.bp_lambda_in[0] ;
 wire \bp_core.bp_lambda_in[1] ;
 wire \bp_core.bp_lambda_in[2] ;
 wire \bp_core.bp_lambda_in[3] ;
 wire \bp_core.bp_lambda_in[4] ;
 wire \bp_core.bp_lambda_in[5] ;
 wire \bp_core.bp_lambda_in[6] ;
 wire \bp_core.bp_lambda_in[7] ;
 wire \bp_core.bp_lambda_out[0] ;
 wire \bp_core.bp_lambda_out[1] ;
 wire \bp_core.bp_lambda_out[2] ;
 wire \bp_core.bp_lambda_out[3] ;
 wire \bp_core.bp_lambda_out[4] ;
 wire \bp_core.bp_lambda_out[5] ;
 wire \bp_core.bp_lambda_out[6] ;
 wire \bp_core.bp_lambda_out[7] ;
 wire \bp_core.bp_param_ack_out ;
 wire \bp_core.bp_param_output_data[0] ;
 wire \bp_core.bp_param_output_data[1] ;
 wire \bp_core.bp_param_output_data[2] ;
 wire \bp_core.bp_param_output_data[3] ;
 wire \bp_core.bp_param_output_data[4] ;
 wire \bp_core.bp_param_output_valid ;
 wire \bp_core.bp_param_valid_in ;
 wire \bp_core.bp_param_valid_out ;
 wire \bp_core.bp_report_addr_out[0] ;
 wire \bp_core.bp_report_addr_out[10] ;
 wire \bp_core.bp_report_addr_out[11] ;
 wire \bp_core.bp_report_addr_out[12] ;
 wire \bp_core.bp_report_addr_out[13] ;
 wire \bp_core.bp_report_addr_out[14] ;
 wire \bp_core.bp_report_addr_out[15] ;
 wire \bp_core.bp_report_addr_out[16] ;
 wire \bp_core.bp_report_addr_out[17] ;
 wire \bp_core.bp_report_addr_out[18] ;
 wire \bp_core.bp_report_addr_out[19] ;
 wire \bp_core.bp_report_addr_out[1] ;
 wire \bp_core.bp_report_addr_out[2] ;
 wire \bp_core.bp_report_addr_out[3] ;
 wire \bp_core.bp_report_addr_out[4] ;
 wire \bp_core.bp_report_addr_out[5] ;
 wire \bp_core.bp_report_addr_out[6] ;
 wire \bp_core.bp_report_addr_out[7] ;
 wire \bp_core.bp_report_addr_out[8] ;
 wire \bp_core.bp_report_addr_out[9] ;
 wire \bp_core.bp_report_valid_out ;
 wire \bp_core.bp_stride_in[0] ;
 wire \bp_core.bp_stride_in[10] ;
 wire \bp_core.bp_stride_in[11] ;
 wire \bp_core.bp_stride_in[12] ;
 wire \bp_core.bp_stride_in[13] ;
 wire \bp_core.bp_stride_in[14] ;
 wire \bp_core.bp_stride_in[15] ;
 wire \bp_core.bp_stride_in[16] ;
 wire \bp_core.bp_stride_in[17] ;
 wire \bp_core.bp_stride_in[18] ;
 wire \bp_core.bp_stride_in[19] ;
 wire \bp_core.bp_stride_in[1] ;
 wire \bp_core.bp_stride_in[2] ;
 wire \bp_core.bp_stride_in[3] ;
 wire \bp_core.bp_stride_in[4] ;
 wire \bp_core.bp_stride_in[5] ;
 wire \bp_core.bp_stride_in[6] ;
 wire \bp_core.bp_stride_in[7] ;
 wire \bp_core.bp_stride_in[8] ;
 wire \bp_core.bp_stride_in[9] ;
 wire \bp_core.bp_stride_out[0] ;
 wire \bp_core.bp_stride_out[10] ;
 wire \bp_core.bp_stride_out[11] ;
 wire \bp_core.bp_stride_out[12] ;
 wire \bp_core.bp_stride_out[13] ;
 wire \bp_core.bp_stride_out[14] ;
 wire \bp_core.bp_stride_out[15] ;
 wire \bp_core.bp_stride_out[16] ;
 wire \bp_core.bp_stride_out[17] ;
 wire \bp_core.bp_stride_out[18] ;
 wire \bp_core.bp_stride_out[19] ;
 wire \bp_core.bp_stride_out[1] ;
 wire \bp_core.bp_stride_out[2] ;
 wire \bp_core.bp_stride_out[3] ;
 wire \bp_core.bp_stride_out[4] ;
 wire \bp_core.bp_stride_out[5] ;
 wire \bp_core.bp_stride_out[6] ;
 wire \bp_core.bp_stride_out[7] ;
 wire \bp_core.bp_stride_out[8] ;
 wire \bp_core.bp_stride_out[9] ;
 wire \bp_core.busy_out ;
 wire \bp_core.data_reg[0] ;
 wire \bp_core.data_reg[1] ;
 wire \bp_core.data_reg[2] ;
 wire \bp_core.data_reg[3] ;
 wire \bp_core.data_reg[4] ;
 wire \bp_core.data_reg[5] ;
 wire \bp_core.data_reg[6] ;
 wire \bp_core.data_reg[7] ;
 wire \bp_core.init_counter[0] ;
 wire \bp_core.init_counter[10] ;
 wire \bp_core.init_counter[11] ;
 wire \bp_core.init_counter[12] ;
 wire \bp_core.init_counter[13] ;
 wire \bp_core.init_counter[14] ;
 wire \bp_core.init_counter[15] ;
 wire \bp_core.init_counter[1] ;
 wire \bp_core.init_counter[2] ;
 wire \bp_core.init_counter[3] ;
 wire \bp_core.init_counter[4] ;
 wire \bp_core.init_counter[5] ;
 wire \bp_core.init_counter[6] ;
 wire \bp_core.init_counter[7] ;
 wire \bp_core.init_counter[8] ;
 wire \bp_core.init_counter[9] ;
 wire \bp_core.initialized ;
 wire \bp_core.params_addr[0] ;
 wire \bp_core.params_addr[10] ;
 wire \bp_core.params_addr[11] ;
 wire \bp_core.params_addr[12] ;
 wire \bp_core.params_addr[13] ;
 wire \bp_core.params_addr[14] ;
 wire \bp_core.params_addr[15] ;
 wire \bp_core.params_addr[16] ;
 wire \bp_core.params_addr[17] ;
 wire \bp_core.params_addr[18] ;
 wire \bp_core.params_addr[19] ;
 wire \bp_core.params_addr[1] ;
 wire \bp_core.params_addr[2] ;
 wire \bp_core.params_addr[3] ;
 wire \bp_core.params_addr[4] ;
 wire \bp_core.params_addr[5] ;
 wire \bp_core.params_addr[6] ;
 wire \bp_core.params_addr[7] ;
 wire \bp_core.params_addr[8] ;
 wire \bp_core.params_addr[9] ;
 wire \bp_core.params_done ;
 wire \bp_core.params_forward ;
 wire \bp_core.params_module.counter[0] ;
 wire \bp_core.params_module.counter[1] ;
 wire \bp_core.params_module.counter[2] ;
 wire \bp_core.params_module.counter[3] ;
 wire \bp_core.params_module.params_ready ;
 wire \bp_core.params_module.start_load ;
 wire \bp_core.params_module.state[0] ;
 wire \bp_core.params_module.state[1] ;
 wire \bp_core.params_module.state[2] ;
 wire \bp_core.params_module.state[3] ;
 wire \bp_core.ram_addr[0] ;
 wire \bp_core.ram_addr[10] ;
 wire \bp_core.ram_addr[11] ;
 wire \bp_core.ram_addr[12] ;
 wire \bp_core.ram_addr[13] ;
 wire \bp_core.ram_addr[14] ;
 wire \bp_core.ram_addr[15] ;
 wire \bp_core.ram_addr[1] ;
 wire \bp_core.ram_addr[2] ;
 wire \bp_core.ram_addr[3] ;
 wire \bp_core.ram_addr[4] ;
 wire \bp_core.ram_addr[5] ;
 wire \bp_core.ram_addr[6] ;
 wire \bp_core.ram_addr[7] ;
 wire \bp_core.ram_addr[8] ;
 wire \bp_core.ram_addr[9] ;
 wire \bp_core.ram_rdata[0] ;
 wire \bp_core.ram_rdata[1] ;
 wire \bp_core.ram_rdata[2] ;
 wire \bp_core.ram_rdata[3] ;
 wire \bp_core.ram_rdata[4] ;
 wire \bp_core.ram_rdata[5] ;
 wire \bp_core.ram_rdata[6] ;
 wire \bp_core.ram_rdata[7] ;
 wire \bp_core.ram_start ;
 wire \bp_core.ram_wdata[0] ;
 wire \bp_core.ram_wdata[1] ;
 wire \bp_core.ram_wdata[2] ;
 wire \bp_core.ram_wdata[3] ;
 wire \bp_core.ram_wdata[4] ;
 wire \bp_core.ram_wdata[5] ;
 wire \bp_core.ram_wdata[6] ;
 wire \bp_core.ram_wdata[7] ;
 wire \bp_core.ram_we ;
 wire \bp_core.state[10] ;
 wire \bp_core.state[11] ;
 wire \bp_core.state[1] ;
 wire \bp_core.state[2] ;
 wire \bp_core.state[3] ;
 wire \bp_core.state[4] ;
 wire \bp_core.state[5] ;
 wire \bp_core.state[6] ;
 wire \bp_core.state[7] ;
 wire \bp_core.state[8] ;
 wire \bp_core.state[9] ;
 wire \bp_core.status_out[0] ;
 wire \bp_core.status_out[1] ;
 wire \bp_core.status_out[2] ;
 wire \bp_core.status_out[3] ;
 wire \bp_core.status_out[4] ;
 wire \bp_core.threshold_load_counter ;
 wire \bp_core.threshold_reg[0] ;
 wire \bp_core.threshold_reg[1] ;
 wire \bp_core.threshold_reg[2] ;
 wire \bp_core.threshold_reg[4] ;
 wire \bp_core.threshold_reg[5] ;
 wire \bp_core.valid_out ;
 wire \inter_bp.bp_report_addr_out[0] ;
 wire \inter_bp.bp_report_addr_out[10] ;
 wire \inter_bp.bp_report_addr_out[11] ;
 wire \inter_bp.bp_report_addr_out[12] ;
 wire \inter_bp.bp_report_addr_out[13] ;
 wire \inter_bp.bp_report_addr_out[14] ;
 wire \inter_bp.bp_report_addr_out[15] ;
 wire \inter_bp.bp_report_addr_out[16] ;
 wire \inter_bp.bp_report_addr_out[17] ;
 wire \inter_bp.bp_report_addr_out[18] ;
 wire \inter_bp.bp_report_addr_out[19] ;
 wire \inter_bp.bp_report_addr_out[1] ;
 wire \inter_bp.bp_report_addr_out[2] ;
 wire \inter_bp.bp_report_addr_out[3] ;
 wire \inter_bp.bp_report_addr_out[4] ;
 wire \inter_bp.bp_report_addr_out[5] ;
 wire \inter_bp.bp_report_addr_out[6] ;
 wire \inter_bp.bp_report_addr_out[7] ;
 wire \inter_bp.bp_report_addr_out[8] ;
 wire \inter_bp.bp_report_addr_out[9] ;
 wire \inter_bp.bp_report_valid_out ;
 wire \inter_bp.from_left_param_valid_prev ;
 wire \inter_bp.from_left_report_valid_prev ;
 wire \inter_bp.param_pending ;
 wire \inter_bp.param_pending_reg[0] ;
 wire \inter_bp.param_pending_reg[10] ;
 wire \inter_bp.param_pending_reg[11] ;
 wire \inter_bp.param_pending_reg[12] ;
 wire \inter_bp.param_pending_reg[13] ;
 wire \inter_bp.param_pending_reg[14] ;
 wire \inter_bp.param_pending_reg[15] ;
 wire \inter_bp.param_pending_reg[16] ;
 wire \inter_bp.param_pending_reg[17] ;
 wire \inter_bp.param_pending_reg[18] ;
 wire \inter_bp.param_pending_reg[19] ;
 wire \inter_bp.param_pending_reg[1] ;
 wire \inter_bp.param_pending_reg[20] ;
 wire \inter_bp.param_pending_reg[21] ;
 wire \inter_bp.param_pending_reg[22] ;
 wire \inter_bp.param_pending_reg[23] ;
 wire \inter_bp.param_pending_reg[24] ;
 wire \inter_bp.param_pending_reg[25] ;
 wire \inter_bp.param_pending_reg[26] ;
 wire \inter_bp.param_pending_reg[27] ;
 wire \inter_bp.param_pending_reg[28] ;
 wire \inter_bp.param_pending_reg[29] ;
 wire \inter_bp.param_pending_reg[2] ;
 wire \inter_bp.param_pending_reg[30] ;
 wire \inter_bp.param_pending_reg[31] ;
 wire \inter_bp.param_pending_reg[32] ;
 wire \inter_bp.param_pending_reg[33] ;
 wire \inter_bp.param_pending_reg[34] ;
 wire \inter_bp.param_pending_reg[35] ;
 wire \inter_bp.param_pending_reg[36] ;
 wire \inter_bp.param_pending_reg[37] ;
 wire \inter_bp.param_pending_reg[38] ;
 wire \inter_bp.param_pending_reg[39] ;
 wire \inter_bp.param_pending_reg[3] ;
 wire \inter_bp.param_pending_reg[40] ;
 wire \inter_bp.param_pending_reg[41] ;
 wire \inter_bp.param_pending_reg[42] ;
 wire \inter_bp.param_pending_reg[43] ;
 wire \inter_bp.param_pending_reg[44] ;
 wire \inter_bp.param_pending_reg[45] ;
 wire \inter_bp.param_pending_reg[46] ;
 wire \inter_bp.param_pending_reg[47] ;
 wire \inter_bp.param_pending_reg[4] ;
 wire \inter_bp.param_pending_reg[5] ;
 wire \inter_bp.param_pending_reg[6] ;
 wire \inter_bp.param_pending_reg[7] ;
 wire \inter_bp.param_pending_reg[8] ;
 wire \inter_bp.param_pending_reg[9] ;
 wire \inter_bp.param_receiving ;
 wire \inter_bp.param_rx_counter[0] ;
 wire \inter_bp.param_rx_counter[1] ;
 wire \inter_bp.param_rx_counter[2] ;
 wire \inter_bp.param_rx_counter[3] ;
 wire \inter_bp.param_rx_counter[4] ;
 wire \inter_bp.param_rx_done ;
 wire \inter_bp.param_shift_reg[0] ;
 wire \inter_bp.param_shift_reg[10] ;
 wire \inter_bp.param_shift_reg[11] ;
 wire \inter_bp.param_shift_reg[12] ;
 wire \inter_bp.param_shift_reg[13] ;
 wire \inter_bp.param_shift_reg[14] ;
 wire \inter_bp.param_shift_reg[15] ;
 wire \inter_bp.param_shift_reg[16] ;
 wire \inter_bp.param_shift_reg[17] ;
 wire \inter_bp.param_shift_reg[18] ;
 wire \inter_bp.param_shift_reg[19] ;
 wire \inter_bp.param_shift_reg[1] ;
 wire \inter_bp.param_shift_reg[20] ;
 wire \inter_bp.param_shift_reg[21] ;
 wire \inter_bp.param_shift_reg[22] ;
 wire \inter_bp.param_shift_reg[23] ;
 wire \inter_bp.param_shift_reg[24] ;
 wire \inter_bp.param_shift_reg[25] ;
 wire \inter_bp.param_shift_reg[26] ;
 wire \inter_bp.param_shift_reg[27] ;
 wire \inter_bp.param_shift_reg[28] ;
 wire \inter_bp.param_shift_reg[29] ;
 wire \inter_bp.param_shift_reg[2] ;
 wire \inter_bp.param_shift_reg[30] ;
 wire \inter_bp.param_shift_reg[31] ;
 wire \inter_bp.param_shift_reg[32] ;
 wire \inter_bp.param_shift_reg[33] ;
 wire \inter_bp.param_shift_reg[34] ;
 wire \inter_bp.param_shift_reg[35] ;
 wire \inter_bp.param_shift_reg[36] ;
 wire \inter_bp.param_shift_reg[37] ;
 wire \inter_bp.param_shift_reg[38] ;
 wire \inter_bp.param_shift_reg[39] ;
 wire \inter_bp.param_shift_reg[3] ;
 wire \inter_bp.param_shift_reg[40] ;
 wire \inter_bp.param_shift_reg[41] ;
 wire \inter_bp.param_shift_reg[42] ;
 wire \inter_bp.param_shift_reg[43] ;
 wire \inter_bp.param_shift_reg[44] ;
 wire \inter_bp.param_shift_reg[45] ;
 wire \inter_bp.param_shift_reg[46] ;
 wire \inter_bp.param_shift_reg[47] ;
 wire \inter_bp.param_shift_reg[4] ;
 wire \inter_bp.param_shift_reg[5] ;
 wire \inter_bp.param_shift_reg[6] ;
 wire \inter_bp.param_shift_reg[7] ;
 wire \inter_bp.param_shift_reg[8] ;
 wire \inter_bp.param_shift_reg[9] ;
 wire \inter_bp.param_transmitting ;
 wire \inter_bp.param_tx_counter[0] ;
 wire \inter_bp.param_tx_counter[1] ;
 wire \inter_bp.param_tx_counter[2] ;
 wire \inter_bp.param_tx_counter[3] ;
 wire \inter_bp.param_tx_counter[4] ;
 wire \inter_bp.param_tx_shift_reg[0] ;
 wire \inter_bp.param_tx_shift_reg[10] ;
 wire \inter_bp.param_tx_shift_reg[11] ;
 wire \inter_bp.param_tx_shift_reg[12] ;
 wire \inter_bp.param_tx_shift_reg[13] ;
 wire \inter_bp.param_tx_shift_reg[14] ;
 wire \inter_bp.param_tx_shift_reg[15] ;
 wire \inter_bp.param_tx_shift_reg[16] ;
 wire \inter_bp.param_tx_shift_reg[17] ;
 wire \inter_bp.param_tx_shift_reg[18] ;
 wire \inter_bp.param_tx_shift_reg[19] ;
 wire \inter_bp.param_tx_shift_reg[1] ;
 wire \inter_bp.param_tx_shift_reg[20] ;
 wire \inter_bp.param_tx_shift_reg[21] ;
 wire \inter_bp.param_tx_shift_reg[22] ;
 wire \inter_bp.param_tx_shift_reg[23] ;
 wire \inter_bp.param_tx_shift_reg[24] ;
 wire \inter_bp.param_tx_shift_reg[25] ;
 wire \inter_bp.param_tx_shift_reg[26] ;
 wire \inter_bp.param_tx_shift_reg[27] ;
 wire \inter_bp.param_tx_shift_reg[28] ;
 wire \inter_bp.param_tx_shift_reg[29] ;
 wire \inter_bp.param_tx_shift_reg[2] ;
 wire \inter_bp.param_tx_shift_reg[30] ;
 wire \inter_bp.param_tx_shift_reg[31] ;
 wire \inter_bp.param_tx_shift_reg[32] ;
 wire \inter_bp.param_tx_shift_reg[33] ;
 wire \inter_bp.param_tx_shift_reg[34] ;
 wire \inter_bp.param_tx_shift_reg[35] ;
 wire \inter_bp.param_tx_shift_reg[36] ;
 wire \inter_bp.param_tx_shift_reg[37] ;
 wire \inter_bp.param_tx_shift_reg[38] ;
 wire \inter_bp.param_tx_shift_reg[39] ;
 wire \inter_bp.param_tx_shift_reg[3] ;
 wire \inter_bp.param_tx_shift_reg[40] ;
 wire \inter_bp.param_tx_shift_reg[41] ;
 wire \inter_bp.param_tx_shift_reg[42] ;
 wire \inter_bp.param_tx_shift_reg[43] ;
 wire \inter_bp.param_tx_shift_reg[44] ;
 wire \inter_bp.param_tx_shift_reg[45] ;
 wire \inter_bp.param_tx_shift_reg[46] ;
 wire \inter_bp.param_tx_shift_reg[47] ;
 wire \inter_bp.param_tx_shift_reg[4] ;
 wire \inter_bp.param_tx_shift_reg[5] ;
 wire \inter_bp.param_tx_shift_reg[6] ;
 wire \inter_bp.param_tx_shift_reg[7] ;
 wire \inter_bp.param_tx_shift_reg[8] ;
 wire \inter_bp.param_tx_shift_reg[9] ;
 wire \inter_bp.report_receiving ;
 wire \inter_bp.report_rx_counter[0] ;
 wire \inter_bp.report_rx_counter[1] ;
 wire \inter_bp.report_rx_counter[2] ;
 wire \inter_bp.report_rx_counter[3] ;
 wire \inter_bp.report_rx_counter[4] ;
 wire \inter_bp.report_rx_done ;
 wire \inter_bp.report_shift_reg[0] ;
 wire \inter_bp.report_shift_reg[10] ;
 wire \inter_bp.report_shift_reg[11] ;
 wire \inter_bp.report_shift_reg[12] ;
 wire \inter_bp.report_shift_reg[13] ;
 wire \inter_bp.report_shift_reg[14] ;
 wire \inter_bp.report_shift_reg[15] ;
 wire \inter_bp.report_shift_reg[16] ;
 wire \inter_bp.report_shift_reg[17] ;
 wire \inter_bp.report_shift_reg[18] ;
 wire \inter_bp.report_shift_reg[19] ;
 wire \inter_bp.report_shift_reg[1] ;
 wire \inter_bp.report_shift_reg[2] ;
 wire \inter_bp.report_shift_reg[3] ;
 wire \inter_bp.report_shift_reg[4] ;
 wire \inter_bp.report_shift_reg[5] ;
 wire \inter_bp.report_shift_reg[6] ;
 wire \inter_bp.report_shift_reg[7] ;
 wire \inter_bp.report_shift_reg[8] ;
 wire \inter_bp.report_shift_reg[9] ;
 wire \inter_bp.report_transmitting ;
 wire \inter_bp.report_tx_counter[0] ;
 wire \inter_bp.report_tx_counter[1] ;
 wire \inter_bp.report_tx_counter[2] ;
 wire \inter_bp.report_tx_counter[3] ;
 wire \inter_bp.report_tx_counter[4] ;
 wire \inter_bp.report_tx_shift_reg[0] ;
 wire \inter_bp.report_tx_shift_reg[10] ;
 wire \inter_bp.report_tx_shift_reg[11] ;
 wire \inter_bp.report_tx_shift_reg[12] ;
 wire \inter_bp.report_tx_shift_reg[13] ;
 wire \inter_bp.report_tx_shift_reg[14] ;
 wire \inter_bp.report_tx_shift_reg[15] ;
 wire \inter_bp.report_tx_shift_reg[16] ;
 wire \inter_bp.report_tx_shift_reg[17] ;
 wire \inter_bp.report_tx_shift_reg[18] ;
 wire \inter_bp.report_tx_shift_reg[19] ;
 wire \inter_bp.report_tx_shift_reg[1] ;
 wire \inter_bp.report_tx_shift_reg[2] ;
 wire \inter_bp.report_tx_shift_reg[3] ;
 wire \inter_bp.report_tx_shift_reg[4] ;
 wire \inter_bp.report_tx_shift_reg[5] ;
 wire \inter_bp.report_tx_shift_reg[6] ;
 wire \inter_bp.report_tx_shift_reg[7] ;
 wire \inter_bp.report_tx_shift_reg[8] ;
 wire \inter_bp.report_tx_shift_reg[9] ;
 wire \inter_bp.serialize_param_valid_prev ;
 wire \inter_bp.serialize_report_valid_prev ;
 wire spi_cs;
 wire \spi_ctrl.addr[0] ;
 wire \spi_ctrl.addr[10] ;
 wire \spi_ctrl.addr[11] ;
 wire \spi_ctrl.addr[12] ;
 wire \spi_ctrl.addr[13] ;
 wire \spi_ctrl.addr[14] ;
 wire \spi_ctrl.addr[15] ;
 wire \spi_ctrl.addr[1] ;
 wire \spi_ctrl.addr[2] ;
 wire \spi_ctrl.addr[3] ;
 wire \spi_ctrl.addr[4] ;
 wire \spi_ctrl.addr[5] ;
 wire \spi_ctrl.addr[6] ;
 wire \spi_ctrl.addr[7] ;
 wire \spi_ctrl.addr[8] ;
 wire \spi_ctrl.addr[9] ;
 wire \spi_ctrl.bits_remaining[0] ;
 wire \spi_ctrl.bits_remaining[1] ;
 wire \spi_ctrl.bits_remaining[2] ;
 wire \spi_ctrl.bits_remaining[3] ;
 wire \spi_ctrl.fsm_state[0] ;
 wire \spi_ctrl.fsm_state[1] ;
 wire clk_regs;
 wire \spi_ctrl.spi_miso_buf ;
 wire \spi_ctrl.spi_mosi ;
 wire \spi_ctrl.writing ;
 wire net49;
 wire net50;
 wire net51;
 wire net15;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net16;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire delaynet_0_clk;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire [0:0] _1799_;
 wire [0:0] _1800_;

 sg13g2_o21ai_1 _1801_ (.B1(_1404_),
    .Y(_1405_),
    .A1(_0770_),
    .A2(_1403_));
 sg13g2_o21ai_1 _1802_ (.B1(_1405_),
    .Y(_1406_),
    .A1(_0540_),
    .A2(net723));
 sg13g2_mux2_1 _1803_ (.A0(_1406_),
    .A1(net1077),
    .S(net567),
    .X(_0321_));
 sg13g2_a21oi_1 _1804_ (.A1(_0770_),
    .A2(_1403_),
    .Y(_1407_),
    .B1(_0768_));
 sg13g2_xnor2_1 _1805_ (.Y(_1408_),
    .A(_0767_),
    .B(_1407_));
 sg13g2_nand2_1 _1806_ (.Y(_1409_),
    .A(net725),
    .B(_1408_));
 sg13g2_o21ai_1 _1807_ (.B1(_1409_),
    .Y(_1410_),
    .A1(_0541_),
    .A2(net723));
 sg13g2_mux2_1 _1808_ (.A0(_1410_),
    .A1(net1087),
    .S(net566),
    .X(_0322_));
 sg13g2_a221oi_1 _1809_ (.B2(_1403_),
    .C1(_0768_),
    .B1(_0770_),
    .A1(\bp_core.addr_reg[13] ),
    .Y(_1411_),
    .A2(\bp_core.bp_stride_out[13] ));
 sg13g2_o21ai_1 _1810_ (.B1(_0762_),
    .Y(_1412_),
    .A1(_0766_),
    .A2(_1411_));
 sg13g2_nor3_1 _1811_ (.A(_0762_),
    .B(_0766_),
    .C(_1411_),
    .Y(_1413_));
 sg13g2_nor2_1 _1812_ (.A(net719),
    .B(_1413_),
    .Y(_1414_));
 sg13g2_nor2_1 _1813_ (.A(_0542_),
    .B(net725),
    .Y(_1415_));
 sg13g2_a21o_1 _1814_ (.A2(_1414_),
    .A1(_1412_),
    .B1(_1415_),
    .X(_1416_));
 sg13g2_mux2_1 _1815_ (.A0(_1416_),
    .A1(net1104),
    .S(net566),
    .X(_0323_));
 sg13g2_o21ai_1 _1816_ (.B1(_0760_),
    .Y(_1417_),
    .A1(_0761_),
    .A2(_1413_));
 sg13g2_or3_1 _1817_ (.A(_0760_),
    .B(_0761_),
    .C(_1413_),
    .X(_1418_));
 sg13g2_nand3_1 _1818_ (.B(_1417_),
    .C(_1418_),
    .A(net725),
    .Y(_1419_));
 sg13g2_o21ai_1 _1819_ (.B1(_1419_),
    .Y(_1420_),
    .A1(_0543_),
    .A2(net725));
 sg13g2_mux2_1 _1820_ (.A0(_1420_),
    .A1(net1047),
    .S(net568),
    .X(_0324_));
 sg13g2_and2_1 _1821_ (.A(net721),
    .B(_0793_),
    .X(_1421_));
 sg13g2_nand2_1 _1822_ (.Y(_1422_),
    .A(net721),
    .B(_0793_));
 sg13g2_a21oi_1 _1823_ (.A1(\bp_core.addr_reg[16] ),
    .A2(net717),
    .Y(_1423_),
    .B1(_1421_));
 sg13g2_mux2_1 _1824_ (.A0(_1423_),
    .A1(net1019),
    .S(net568),
    .X(_0325_));
 sg13g2_nand2_1 _1825_ (.Y(_1424_),
    .A(net721),
    .B(_0796_));
 sg13g2_xor2_1 _1826_ (.B(\bp_core.addr_reg[16] ),
    .A(\bp_core.addr_reg[17] ),
    .X(_1425_));
 sg13g2_a21oi_1 _1827_ (.A1(net717),
    .A2(_1425_),
    .Y(_1426_),
    .B1(_1421_));
 sg13g2_mux2_1 _1828_ (.A0(_0793_),
    .A1(_1426_),
    .S(_1424_),
    .X(_1427_));
 sg13g2_mux2_1 _1829_ (.A0(_1427_),
    .A1(net102),
    .S(net568),
    .X(_0326_));
 sg13g2_o21ai_1 _1830_ (.B1(_0804_),
    .Y(_1428_),
    .A1(_0793_),
    .A2(_0796_));
 sg13g2_o21ai_1 _1831_ (.B1(net482),
    .Y(_1429_),
    .A1(net932),
    .A2(\bp_core.addr_reg[16] ));
 sg13g2_nor2_1 _1832_ (.A(net721),
    .B(_0726_),
    .Y(_1430_));
 sg13g2_a22oi_1 _1833_ (.Y(_1431_),
    .B1(_1429_),
    .B2(_1430_),
    .A2(_1428_),
    .A1(_0809_));
 sg13g2_mux2_1 _1834_ (.A0(_1431_),
    .A1(net1065),
    .S(net568),
    .X(_0327_));
 sg13g2_or2_1 _1835_ (.X(_1432_),
    .B(_0808_),
    .A(_0805_));
 sg13g2_xnor2_1 _1836_ (.Y(_1433_),
    .A(\bp_core.addr_reg[19] ),
    .B(_0726_));
 sg13g2_a22oi_1 _1837_ (.Y(_1434_),
    .B1(_1433_),
    .B2(net717),
    .A2(_1432_),
    .A1(_0810_));
 sg13g2_mux2_1 _1838_ (.A0(_1434_),
    .A1(net1038),
    .S(net568),
    .X(_0328_));
 sg13g2_a21oi_1 _1839_ (.A1(net198),
    .A2(\bp_core.params_forward ),
    .Y(_1435_),
    .B1(net58));
 sg13g2_a21oi_1 _1840_ (.A1(_0556_),
    .A2(\bp_core.params_module.state[0] ),
    .Y(_0329_),
    .B1(_1435_));
 sg13g2_o21ai_1 _1841_ (.B1(_1322_),
    .Y(_1436_),
    .A1(_0526_),
    .A2(_1315_));
 sg13g2_o21ai_1 _1842_ (.B1(net657),
    .Y(_1437_),
    .A1(net730),
    .A2(_0628_));
 sg13g2_mux2_1 _1843_ (.A0(_1437_),
    .A1(net1117),
    .S(_1436_),
    .X(_0330_));
 sg13g2_o21ai_1 _1844_ (.B1(net656),
    .Y(_1438_),
    .A1(net728),
    .A2(_0630_));
 sg13g2_mux2_1 _1845_ (.A0(_1438_),
    .A1(net1145),
    .S(_1436_),
    .X(_0331_));
 sg13g2_o21ai_1 _1846_ (.B1(net655),
    .Y(_1439_),
    .A1(net730),
    .A2(_0632_));
 sg13g2_nor2_1 _1847_ (.A(_1436_),
    .B(_1439_),
    .Y(_1440_));
 sg13g2_a21oi_1 _1848_ (.A1(_0544_),
    .A2(_1436_),
    .Y(_0332_),
    .B1(_1440_));
 sg13g2_o21ai_1 _1849_ (.B1(net654),
    .Y(_1441_),
    .A1(net730),
    .A2(_0634_));
 sg13g2_mux2_1 _1850_ (.A0(_1441_),
    .A1(net1150),
    .S(_1436_),
    .X(_0333_));
 sg13g2_o21ai_1 _1851_ (.B1(net653),
    .Y(_1442_),
    .A1(net728),
    .A2(_0636_));
 sg13g2_mux2_1 _1852_ (.A0(_1442_),
    .A1(net1136),
    .S(_1436_),
    .X(_0334_));
 sg13g2_nor3_1 _1853_ (.A(\bp_core.params_module.counter[3] ),
    .B(\bp_core.params_module.counter[2] ),
    .C(net738),
    .Y(_1443_));
 sg13g2_and2_1 _1854_ (.A(\bp_core.params_module.counter[0] ),
    .B(_1443_),
    .X(_1444_));
 sg13g2_inv_1 _1855_ (.Y(_1445_),
    .A(_1444_));
 sg13g2_nor3_2 _1856_ (.A(net738),
    .B(\bp_core.params_module.counter[0] ),
    .C(_1314_),
    .Y(_1446_));
 sg13g2_inv_1 _1857_ (.Y(_1447_),
    .A(_1446_));
 sg13g2_nand2_1 _1858_ (.Y(_1448_),
    .A(\bp_core.bp_stride_out[10] ),
    .B(_1342_));
 sg13g2_nor3_2 _1859_ (.A(\bp_core.params_module.counter[3] ),
    .B(\bp_core.params_module.counter[2] ),
    .C(_1309_),
    .Y(_1449_));
 sg13g2_nor3_2 _1860_ (.A(\bp_core.params_module.counter[3] ),
    .B(\bp_core.params_module.counter[2] ),
    .C(_1341_),
    .Y(_1450_));
 sg13g2_o21ai_1 _1861_ (.B1(\bp_core.params_module.counter[3] ),
    .Y(_1451_),
    .A1(\bp_core.params_module.counter[2] ),
    .A2(net738));
 sg13g2_nand2_2 _1862_ (.Y(_1452_),
    .A(_0524_),
    .B(_1443_));
 sg13g2_and2_1 _1863_ (.A(_1451_),
    .B(_1452_),
    .X(_1453_));
 sg13g2_a22oi_1 _1864_ (.Y(_1454_),
    .B1(_1449_),
    .B2(\bp_addr_out[15] ),
    .A2(_1323_),
    .A1(\bp_core.bp_stride_out[5] ));
 sg13g2_nand3_1 _1865_ (.B(_1453_),
    .C(_1454_),
    .A(_1448_),
    .Y(_1455_));
 sg13g2_a22oi_1 _1866_ (.Y(_1456_),
    .B1(_0720_),
    .B2(\bp_core.bp_lambda_out[5] ),
    .A2(_0718_),
    .A1(\bp_core.bp_lambda_out[0] ));
 sg13g2_a22oi_1 _1867_ (.Y(_1457_),
    .B1(_1446_),
    .B2(\bp_core.bp_stride_out[0] ),
    .A2(_1315_),
    .A1(\bp_core.bp_stride_out[15] ));
 sg13g2_a22oi_1 _1868_ (.Y(_1458_),
    .B1(_1450_),
    .B2(\bp_addr_out[10] ),
    .A2(_1444_),
    .A1(\bp_addr_out[5] ));
 sg13g2_nand3_1 _1869_ (.B(_1457_),
    .C(_1458_),
    .A(_1456_),
    .Y(_1459_));
 sg13g2_nor2_1 _1870_ (.A(_1455_),
    .B(_1459_),
    .Y(_1460_));
 sg13g2_and2_1 _1871_ (.A(net59),
    .B(_1451_),
    .X(_1461_));
 sg13g2_nand2_2 _1872_ (.Y(_1462_),
    .A(net59),
    .B(_1451_));
 sg13g2_o21ai_1 _1873_ (.B1(_1461_),
    .Y(_1463_),
    .A1(\bp_addr_out[0] ),
    .A2(_1452_));
 sg13g2_nand2_1 _1874_ (.Y(_1464_),
    .A(net459),
    .B(_1462_));
 sg13g2_o21ai_1 _1875_ (.B1(_1464_),
    .Y(_0335_),
    .A1(_1460_),
    .A2(_1463_));
 sg13g2_a22oi_1 _1876_ (.Y(_1465_),
    .B1(_0720_),
    .B2(\bp_core.bp_lambda_out[6] ),
    .A2(_0718_),
    .A1(\bp_core.bp_lambda_out[1] ));
 sg13g2_a22oi_1 _1877_ (.Y(_1466_),
    .B1(_1446_),
    .B2(\bp_core.bp_stride_out[1] ),
    .A2(_1323_),
    .A1(\bp_core.bp_stride_out[6] ));
 sg13g2_a22oi_1 _1878_ (.Y(_1467_),
    .B1(_1450_),
    .B2(\bp_addr_out[11] ),
    .A2(_1315_),
    .A1(\bp_core.bp_stride_out[16] ));
 sg13g2_nand2_1 _1879_ (.Y(_1468_),
    .A(\bp_core.bp_stride_out[11] ),
    .B(_1342_));
 sg13g2_a22oi_1 _1880_ (.Y(_1469_),
    .B1(_1449_),
    .B2(\bp_addr_out[16] ),
    .A2(_1444_),
    .A1(\bp_addr_out[6] ));
 sg13g2_nand3_1 _1881_ (.B(_1468_),
    .C(_1469_),
    .A(_1453_),
    .Y(_1470_));
 sg13g2_nand3_1 _1882_ (.B(_1466_),
    .C(_1467_),
    .A(_1465_),
    .Y(_1471_));
 sg13g2_nor2_1 _1883_ (.A(_1470_),
    .B(_1471_),
    .Y(_1472_));
 sg13g2_o21ai_1 _1884_ (.B1(_1461_),
    .Y(_1473_),
    .A1(\bp_addr_out[1] ),
    .A2(_1452_));
 sg13g2_nand2_1 _1885_ (.Y(_1474_),
    .A(net290),
    .B(_1462_));
 sg13g2_o21ai_1 _1886_ (.B1(_1474_),
    .Y(_0336_),
    .A1(_1472_),
    .A2(_1473_));
 sg13g2_a22oi_1 _1887_ (.Y(_1475_),
    .B1(_0720_),
    .B2(\bp_core.bp_lambda_out[7] ),
    .A2(_0718_),
    .A1(\bp_core.bp_lambda_out[2] ));
 sg13g2_nand2_1 _1888_ (.Y(_1476_),
    .A(\bp_core.bp_stride_out[7] ),
    .B(_1323_));
 sg13g2_a22oi_1 _1889_ (.Y(_1477_),
    .B1(_1449_),
    .B2(\bp_addr_out[17] ),
    .A2(_1446_),
    .A1(\bp_core.bp_stride_out[2] ));
 sg13g2_nand3_1 _1890_ (.B(_1476_),
    .C(_1477_),
    .A(_1453_),
    .Y(_1478_));
 sg13g2_a22oi_1 _1891_ (.Y(_1479_),
    .B1(_1444_),
    .B2(\bp_addr_out[7] ),
    .A2(_1342_),
    .A1(\bp_core.bp_stride_out[12] ));
 sg13g2_a22oi_1 _1892_ (.Y(_1480_),
    .B1(_1450_),
    .B2(\bp_addr_out[12] ),
    .A2(_1315_),
    .A1(\bp_core.bp_stride_out[17] ));
 sg13g2_nand3_1 _1893_ (.B(_1479_),
    .C(_1480_),
    .A(_1475_),
    .Y(_1481_));
 sg13g2_nor2_1 _1894_ (.A(_1478_),
    .B(_1481_),
    .Y(_1482_));
 sg13g2_o21ai_1 _1895_ (.B1(_1461_),
    .Y(_1483_),
    .A1(\bp_addr_out[2] ),
    .A2(_1452_));
 sg13g2_nand2_1 _1896_ (.Y(_1484_),
    .A(net952),
    .B(_1462_));
 sg13g2_o21ai_1 _1897_ (.B1(_1484_),
    .Y(_0337_),
    .A1(_1482_),
    .A2(_1483_));
 sg13g2_a22oi_1 _1898_ (.Y(_1485_),
    .B1(_1444_),
    .B2(\bp_addr_out[8] ),
    .A2(_1315_),
    .A1(\bp_core.bp_stride_out[18] ));
 sg13g2_a22oi_1 _1899_ (.Y(_1486_),
    .B1(_1446_),
    .B2(\bp_core.bp_stride_out[3] ),
    .A2(_1342_),
    .A1(\bp_core.bp_stride_out[13] ));
 sg13g2_nand2_1 _1900_ (.Y(_1487_),
    .A(_1485_),
    .B(_1486_));
 sg13g2_a22oi_1 _1901_ (.Y(_1488_),
    .B1(_1323_),
    .B2(\bp_core.bp_stride_out[8] ),
    .A2(_0718_),
    .A1(\bp_core.bp_lambda_out[3] ));
 sg13g2_a22oi_1 _1902_ (.Y(_1489_),
    .B1(_1450_),
    .B2(\bp_addr_out[13] ),
    .A2(_1449_),
    .A1(\bp_addr_out[18] ));
 sg13g2_nand3_1 _1903_ (.B(_1488_),
    .C(_1489_),
    .A(_1453_),
    .Y(_1490_));
 sg13g2_nor2_1 _1904_ (.A(_1487_),
    .B(_1490_),
    .Y(_1491_));
 sg13g2_o21ai_1 _1905_ (.B1(_1461_),
    .Y(_1492_),
    .A1(\bp_addr_out[3] ),
    .A2(_1452_));
 sg13g2_nand2_1 _1906_ (.Y(_1493_),
    .A(net296),
    .B(_1462_));
 sg13g2_o21ai_1 _1907_ (.B1(_1493_),
    .Y(_0338_),
    .A1(_1491_),
    .A2(_1492_));
 sg13g2_a22oi_1 _1908_ (.Y(_1494_),
    .B1(_1450_),
    .B2(\bp_addr_out[14] ),
    .A2(_1449_),
    .A1(\bp_addr_out[19] ));
 sg13g2_a22oi_1 _1909_ (.Y(_1495_),
    .B1(_1342_),
    .B2(\bp_core.bp_stride_out[14] ),
    .A2(_1323_),
    .A1(\bp_core.bp_stride_out[9] ));
 sg13g2_nand3_1 _1910_ (.B(_1494_),
    .C(_1495_),
    .A(_1453_),
    .Y(_1496_));
 sg13g2_a22oi_1 _1911_ (.Y(_1497_),
    .B1(_1444_),
    .B2(\bp_addr_out[9] ),
    .A2(_0718_),
    .A1(\bp_core.bp_lambda_out[4] ));
 sg13g2_a22oi_1 _1912_ (.Y(_1498_),
    .B1(_1446_),
    .B2(\bp_core.bp_stride_out[4] ),
    .A2(_1315_),
    .A1(\bp_core.bp_stride_out[19] ));
 sg13g2_nand2_1 _1913_ (.Y(_1499_),
    .A(_1497_),
    .B(_1498_));
 sg13g2_nor2_1 _1914_ (.A(_1496_),
    .B(_1499_),
    .Y(_1500_));
 sg13g2_o21ai_1 _1915_ (.B1(_1461_),
    .Y(_1501_),
    .A1(\bp_addr_out[4] ),
    .A2(_1452_));
 sg13g2_nand2_1 _1916_ (.Y(_1502_),
    .A(net959),
    .B(_1462_));
 sg13g2_o21ai_1 _1917_ (.B1(_1502_),
    .Y(_0339_),
    .A1(_1500_),
    .A2(_1501_));
 sg13g2_o21ai_1 _1918_ (.B1(_1322_),
    .Y(_1503_),
    .A1(_0526_),
    .A2(_1449_));
 sg13g2_o21ai_1 _1919_ (.B1(net657),
    .Y(_1504_),
    .A1(net729),
    .A2(_0590_));
 sg13g2_mux2_1 _1920_ (.A0(_1504_),
    .A1(net1024),
    .S(_1503_),
    .X(_0340_));
 sg13g2_o21ai_1 _1921_ (.B1(net656),
    .Y(_1505_),
    .A1(net728),
    .A2(_0592_));
 sg13g2_mux2_1 _1922_ (.A0(_1505_),
    .A1(net974),
    .S(_1503_),
    .X(_0341_));
 sg13g2_o21ai_1 _1923_ (.B1(net655),
    .Y(_1506_),
    .A1(net728),
    .A2(_0594_));
 sg13g2_mux2_1 _1924_ (.A0(_1506_),
    .A1(net985),
    .S(_1503_),
    .X(_0342_));
 sg13g2_o21ai_1 _1925_ (.B1(net654),
    .Y(_1507_),
    .A1(net728),
    .A2(_0596_));
 sg13g2_mux2_1 _1926_ (.A0(_1507_),
    .A1(net877),
    .S(_1503_),
    .X(_0343_));
 sg13g2_o21ai_1 _1927_ (.B1(net653),
    .Y(_1508_),
    .A1(net728),
    .A2(_0598_));
 sg13g2_mux2_1 _1928_ (.A0(_1508_),
    .A1(net1036),
    .S(_1503_),
    .X(_0344_));
 sg13g2_nand2_1 _1929_ (.Y(_1509_),
    .A(\bp_core.bp_lambda_out[0] ),
    .B(\bp_core.ram_rdata[0] ));
 sg13g2_or2_1 _1930_ (.X(_1510_),
    .B(\bp_core.ram_rdata[0] ),
    .A(\bp_core.bp_lambda_out[0] ));
 sg13g2_a21oi_1 _1931_ (.A1(_1509_),
    .A2(_1510_),
    .Y(_1511_),
    .B1(net609));
 sg13g2_a21oi_1 _1932_ (.A1(_0665_),
    .A2(net609),
    .Y(_0345_),
    .B1(_1511_));
 sg13g2_nand2_1 _1933_ (.Y(_1512_),
    .A(\bp_core.bp_lambda_out[1] ),
    .B(\bp_core.ram_rdata[1] ));
 sg13g2_nor2_1 _1934_ (.A(\bp_core.bp_lambda_out[1] ),
    .B(\bp_core.ram_rdata[1] ),
    .Y(_1513_));
 sg13g2_xor2_1 _1935_ (.B(\bp_core.ram_rdata[1] ),
    .A(\bp_core.bp_lambda_out[1] ),
    .X(_1514_));
 sg13g2_xnor2_1 _1936_ (.Y(_1515_),
    .A(_1509_),
    .B(_1514_));
 sg13g2_nor2_1 _1937_ (.A(net609),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_a21oi_1 _1938_ (.A1(_0664_),
    .A2(net609),
    .Y(_0346_),
    .B1(_1516_));
 sg13g2_and2_1 _1939_ (.A(\bp_core.bp_lambda_out[2] ),
    .B(\bp_core.ram_rdata[2] ),
    .X(_1517_));
 sg13g2_xnor2_1 _1940_ (.Y(_1518_),
    .A(\bp_core.bp_lambda_out[2] ),
    .B(\bp_core.ram_rdata[2] ));
 sg13g2_o21ai_1 _1941_ (.B1(_1512_),
    .Y(_1519_),
    .A1(_1509_),
    .A2(_1513_));
 sg13g2_nor2b_1 _1942_ (.A(_1518_),
    .B_N(_1519_),
    .Y(_1520_));
 sg13g2_xnor2_1 _1943_ (.Y(_1521_),
    .A(_1518_),
    .B(_1519_));
 sg13g2_nor2_1 _1944_ (.A(net609),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_a21oi_1 _1945_ (.A1(_0662_),
    .A2(net609),
    .Y(_0347_),
    .B1(_1522_));
 sg13g2_nand2_1 _1946_ (.Y(_1523_),
    .A(\bp_core.bp_lambda_out[3] ),
    .B(\bp_core.ram_rdata[3] ));
 sg13g2_xor2_1 _1947_ (.B(\bp_core.ram_rdata[3] ),
    .A(\bp_core.bp_lambda_out[3] ),
    .X(_1524_));
 sg13g2_or3_1 _1948_ (.A(_1517_),
    .B(_1520_),
    .C(_1524_),
    .X(_1525_));
 sg13g2_o21ai_1 _1949_ (.B1(_1524_),
    .Y(_1526_),
    .A1(_1517_),
    .A2(_1520_));
 sg13g2_a21oi_1 _1950_ (.A1(_1525_),
    .A2(_1526_),
    .Y(_1527_),
    .B1(net610));
 sg13g2_a21oi_1 _1951_ (.A1(_0660_),
    .A2(net609),
    .Y(_0348_),
    .B1(_1527_));
 sg13g2_xnor2_1 _1952_ (.Y(_1528_),
    .A(\bp_core.bp_lambda_out[4] ),
    .B(net363));
 sg13g2_and3_1 _1953_ (.X(_1529_),
    .A(_1523_),
    .B(_1526_),
    .C(_1528_));
 sg13g2_a21oi_1 _1954_ (.A1(_1523_),
    .A2(_1526_),
    .Y(_1530_),
    .B1(_1528_));
 sg13g2_nor2_1 _1955_ (.A(_1529_),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_nor2_1 _1956_ (.A(net610),
    .B(_1531_),
    .Y(_1532_));
 sg13g2_a21oi_1 _1957_ (.A1(_0659_),
    .A2(_0817_),
    .Y(_0349_),
    .B1(_1532_));
 sg13g2_nand2_1 _1958_ (.Y(_1533_),
    .A(\bp_core.bp_lambda_out[5] ),
    .B(\bp_core.ram_rdata[5] ));
 sg13g2_nor2_1 _1959_ (.A(\bp_core.bp_lambda_out[5] ),
    .B(\bp_core.ram_rdata[5] ),
    .Y(_1534_));
 sg13g2_xor2_1 _1960_ (.B(\bp_core.ram_rdata[5] ),
    .A(\bp_core.bp_lambda_out[5] ),
    .X(_1535_));
 sg13g2_a21oi_1 _1961_ (.A1(\bp_core.bp_lambda_out[4] ),
    .A2(\bp_core.ram_rdata[4] ),
    .Y(_1536_),
    .B1(_1530_));
 sg13g2_xnor2_1 _1962_ (.Y(_1537_),
    .A(_1535_),
    .B(_1536_));
 sg13g2_nor2_1 _1963_ (.A(net610),
    .B(_1537_),
    .Y(_1538_));
 sg13g2_a21oi_1 _1964_ (.A1(_0658_),
    .A2(net610),
    .Y(_0350_),
    .B1(_1538_));
 sg13g2_o21ai_1 _1965_ (.B1(_1533_),
    .Y(_1539_),
    .A1(_1534_),
    .A2(_1536_));
 sg13g2_and2_1 _1966_ (.A(\bp_core.bp_lambda_out[6] ),
    .B(net331),
    .X(_1540_));
 sg13g2_xor2_1 _1967_ (.B(net331),
    .A(\bp_core.bp_lambda_out[6] ),
    .X(_1541_));
 sg13g2_xor2_1 _1968_ (.B(net400),
    .A(_1539_),
    .X(_1542_));
 sg13g2_nor2_1 _1969_ (.A(net610),
    .B(_1542_),
    .Y(_1543_));
 sg13g2_a21oi_1 _1970_ (.A1(_0657_),
    .A2(net610),
    .Y(_0351_),
    .B1(_1543_));
 sg13g2_a21oi_1 _1971_ (.A1(_1539_),
    .A2(_1541_),
    .Y(_1544_),
    .B1(_1540_));
 sg13g2_xor2_1 _1972_ (.B(\bp_core.ram_rdata[7] ),
    .A(net234),
    .X(_1545_));
 sg13g2_o21ai_1 _1973_ (.B1(_0011_),
    .Y(_1546_),
    .A1(_1544_),
    .A2(_1545_));
 sg13g2_a21oi_1 _1974_ (.A1(_1544_),
    .A2(_1545_),
    .Y(_1547_),
    .B1(_1546_));
 sg13g2_a21oi_1 _1975_ (.A1(_0656_),
    .A2(net610),
    .Y(_0352_),
    .B1(_1547_));
 sg13g2_nor2_1 _1976_ (.A(\bp_core.state[2] ),
    .B(_0970_),
    .Y(_1548_));
 sg13g2_nor2_1 _1977_ (.A(_0012_),
    .B(_1548_),
    .Y(_1549_));
 sg13g2_o21ai_1 _1978_ (.B1(_1356_),
    .Y(_1550_),
    .A1(net722),
    .A2(_0667_));
 sg13g2_nor2_1 _1979_ (.A(net622),
    .B(_1550_),
    .Y(_1551_));
 sg13g2_a21oi_1 _1980_ (.A1(_0527_),
    .A2(net622),
    .Y(_0353_),
    .B1(_1551_));
 sg13g2_a21oi_1 _1981_ (.A1(net720),
    .A2(net1016),
    .Y(_1552_),
    .B1(net621));
 sg13g2_a22oi_1 _1982_ (.Y(_0354_),
    .B1(_1552_),
    .B2(_1359_),
    .A2(net617),
    .A1(_0528_));
 sg13g2_a21oi_1 _1983_ (.A1(net719),
    .A2(net955),
    .Y(_1553_),
    .B1(net621));
 sg13g2_a22oi_1 _1984_ (.Y(_0355_),
    .B1(_1553_),
    .B2(_1363_),
    .A2(net617),
    .A1(_0529_));
 sg13g2_a21oi_1 _1985_ (.A1(net719),
    .A2(net1035),
    .Y(_1554_),
    .B1(net621));
 sg13g2_a22oi_1 _1986_ (.Y(_0356_),
    .B1(_1554_),
    .B2(_1367_),
    .A2(net617),
    .A1(_0530_));
 sg13g2_a21oi_1 _1987_ (.A1(net720),
    .A2(net986),
    .Y(_1555_),
    .B1(net620));
 sg13g2_a22oi_1 _1988_ (.Y(_0357_),
    .B1(_1555_),
    .B2(net1101),
    .A2(net620),
    .A1(_0531_));
 sg13g2_a21oi_1 _1989_ (.A1(net718),
    .A2(net976),
    .Y(_1556_),
    .B1(net618));
 sg13g2_a22oi_1 _1990_ (.Y(_0358_),
    .B1(_1556_),
    .B2(_1375_),
    .A2(net620),
    .A1(_0532_));
 sg13g2_a21oi_1 _1991_ (.A1(net718),
    .A2(net989),
    .Y(_1557_),
    .B1(net619));
 sg13g2_a22oi_1 _1992_ (.Y(_0359_),
    .B1(_1557_),
    .B2(_1380_),
    .A2(net620),
    .A1(_0533_));
 sg13g2_a21oi_1 _1993_ (.A1(net720),
    .A2(net1029),
    .Y(_1558_),
    .B1(net621));
 sg13g2_a22oi_1 _1994_ (.Y(_0360_),
    .B1(_1558_),
    .B2(_1384_),
    .A2(net620),
    .A1(_0534_));
 sg13g2_a21oi_1 _1995_ (.A1(net718),
    .A2(net1010),
    .Y(_1559_),
    .B1(net619));
 sg13g2_a22oi_1 _1996_ (.Y(_0361_),
    .B1(_1559_),
    .B2(_1387_),
    .A2(net618),
    .A1(_0535_));
 sg13g2_a21oi_1 _1997_ (.A1(net718),
    .A2(net957),
    .Y(_1560_),
    .B1(net618));
 sg13g2_a22oi_1 _1998_ (.Y(_0362_),
    .B1(_1560_),
    .B2(_1392_),
    .A2(net619),
    .A1(_0536_));
 sg13g2_a21oi_1 _1999_ (.A1(net718),
    .A2(net988),
    .Y(_1561_),
    .B1(net618));
 sg13g2_a22oi_1 _2000_ (.Y(_0363_),
    .B1(_1561_),
    .B2(_1397_),
    .A2(net618),
    .A1(_0537_));
 sg13g2_a21oi_1 _2001_ (.A1(net718),
    .A2(net979),
    .Y(_1562_),
    .B1(net618));
 sg13g2_a22oi_1 _2002_ (.Y(_0364_),
    .B1(_1562_),
    .B2(_1401_),
    .A2(net618),
    .A1(_0538_));
 sg13g2_a21oi_1 _2003_ (.A1(net718),
    .A2(net1011),
    .Y(_1563_),
    .B1(net618));
 sg13g2_a22oi_1 _2004_ (.Y(_0365_),
    .B1(_1563_),
    .B2(_1405_),
    .A2(net619),
    .A1(_0540_));
 sg13g2_a21oi_1 _2005_ (.A1(net719),
    .A2(net1037),
    .Y(_1564_),
    .B1(net617));
 sg13g2_a22oi_1 _2006_ (.Y(_0366_),
    .B1(_1564_),
    .B2(_1409_),
    .A2(net620),
    .A1(_0541_));
 sg13g2_a221oi_1 _2007_ (.B2(_1414_),
    .C1(net617),
    .B1(_1412_),
    .A1(net719),
    .Y(_1565_),
    .A2(net1046));
 sg13g2_a21oi_1 _2008_ (.A1(_0542_),
    .A2(net617),
    .Y(_0367_),
    .B1(_1565_));
 sg13g2_a21oi_1 _2009_ (.A1(net719),
    .A2(net1024),
    .Y(_1566_),
    .B1(net617));
 sg13g2_a22oi_1 _2010_ (.Y(_0368_),
    .B1(_1566_),
    .B2(_1419_),
    .A2(net617),
    .A1(_0543_));
 sg13g2_a21oi_1 _2011_ (.A1(net717),
    .A2(net974),
    .Y(_1567_),
    .B1(net616));
 sg13g2_a22oi_1 _2012_ (.Y(_0369_),
    .B1(_1567_),
    .B2(_1422_),
    .A2(net616),
    .A1(_0546_));
 sg13g2_a21oi_1 _2013_ (.A1(net717),
    .A2(net985),
    .Y(_1568_),
    .B1(net616));
 sg13g2_a22oi_1 _2014_ (.Y(_0370_),
    .B1(_1568_),
    .B2(_1424_),
    .A2(net616),
    .A1(_0545_));
 sg13g2_nand2_1 _2015_ (.Y(_1569_),
    .A(net482),
    .B(net616));
 sg13g2_or2_1 _2016_ (.X(_1570_),
    .B(\bp_core.params_addr[18] ),
    .A(net721));
 sg13g2_o21ai_1 _2017_ (.B1(_1570_),
    .Y(_1571_),
    .A1(net717),
    .A2(_0804_));
 sg13g2_o21ai_1 _2018_ (.B1(_1569_),
    .Y(_0371_),
    .A1(net616),
    .A2(_1571_));
 sg13g2_nor2_1 _2019_ (.A(net721),
    .B(net1036),
    .Y(_1572_));
 sg13g2_nor3_1 _2020_ (.A(_0821_),
    .B(net616),
    .C(_1572_),
    .Y(_1573_));
 sg13g2_a21o_1 _2021_ (.A2(net616),
    .A1(net1092),
    .B1(_1573_),
    .X(_0372_));
 sg13g2_nand3_1 _2022_ (.B(_0685_),
    .C(_0687_),
    .A(\bp_core.state[9] ),
    .Y(_1574_));
 sg13g2_nand3b_1 _2023_ (.B(_0102_),
    .C(net755),
    .Y(_1575_),
    .A_N(\bp_core.state[4] ));
 sg13g2_a21o_2 _2024_ (.A2(net359),
    .A1(\bp_core.state[9] ),
    .B1(_0814_),
    .X(_1576_));
 sg13g2_nand2b_1 _2025_ (.Y(_1577_),
    .B(_0685_),
    .A_N(_1576_));
 sg13g2_nand4_1 _2026_ (.B(_1574_),
    .C(_1575_),
    .A(_0825_),
    .Y(_1578_),
    .D(_1577_));
 sg13g2_nor3_1 _2027_ (.A(net756),
    .B(\bp_core.state[4] ),
    .C(\bp_core.bp_param_valid_in ),
    .Y(_1579_));
 sg13g2_nand2b_1 _2028_ (.Y(_1580_),
    .B(net755),
    .A_N(_1579_));
 sg13g2_o21ai_1 _2029_ (.B1(_1580_),
    .Y(_1581_),
    .A1(\bp_core.state[9] ),
    .A2(_0686_));
 sg13g2_mux2_1 _2030_ (.A0(_1581_),
    .A1(net454),
    .S(_1578_),
    .X(_0373_));
 sg13g2_a21oi_1 _2031_ (.A1(net1042),
    .A2(_0687_),
    .Y(_1582_),
    .B1(_0686_));
 sg13g2_nand2_2 _2032_ (.Y(_1583_),
    .A(_1576_),
    .B(_1582_));
 sg13g2_nor2_1 _2033_ (.A(_0689_),
    .B(_0706_),
    .Y(_1584_));
 sg13g2_mux2_1 _2034_ (.A0(net585),
    .A1(net615),
    .S(net1146),
    .X(_0374_));
 sg13g2_xor2_1 _2035_ (.B(\bp_core.init_counter[0] ),
    .A(net1108),
    .X(_1585_));
 sg13g2_a22oi_1 _2036_ (.Y(_1586_),
    .B1(net585),
    .B2(_1585_),
    .A2(net614),
    .A1(net1108));
 sg13g2_inv_1 _2037_ (.Y(_0375_),
    .A(net1109));
 sg13g2_a21o_1 _2038_ (.A2(\bp_core.init_counter[0] ),
    .A1(\bp_core.init_counter[1] ),
    .B1(net1053),
    .X(_1587_));
 sg13g2_and2_1 _2039_ (.A(_0690_),
    .B(_1587_),
    .X(_1588_));
 sg13g2_a22oi_1 _2040_ (.Y(_1589_),
    .B1(net585),
    .B2(_1588_),
    .A2(net615),
    .A1(net1053));
 sg13g2_inv_1 _2041_ (.Y(_0376_),
    .A(net1054));
 sg13g2_xnor2_1 _2042_ (.Y(_1590_),
    .A(net1033),
    .B(_0690_));
 sg13g2_a22oi_1 _2043_ (.Y(_1591_),
    .B1(net585),
    .B2(_1590_),
    .A2(net615),
    .A1(net1033));
 sg13g2_inv_1 _2044_ (.Y(_0377_),
    .A(net1034));
 sg13g2_xor2_1 _2045_ (.B(_0691_),
    .A(net1044),
    .X(_1592_));
 sg13g2_a22oi_1 _2046_ (.Y(_1593_),
    .B1(net584),
    .B2(_1592_),
    .A2(net614),
    .A1(net1044));
 sg13g2_inv_1 _2047_ (.Y(_0378_),
    .A(net1045));
 sg13g2_xor2_1 _2048_ (.B(_0692_),
    .A(net1111),
    .X(_1594_));
 sg13g2_a22oi_1 _2049_ (.Y(_1595_),
    .B1(net584),
    .B2(_1594_),
    .A2(net614),
    .A1(net1111));
 sg13g2_inv_1 _2050_ (.Y(_0379_),
    .A(_1595_));
 sg13g2_a21o_1 _2051_ (.A2(_0692_),
    .A1(\bp_core.init_counter[5] ),
    .B1(net1030),
    .X(_1596_));
 sg13g2_and2_1 _2052_ (.A(_0693_),
    .B(net584),
    .X(_1597_));
 sg13g2_a22oi_1 _2053_ (.Y(_1598_),
    .B1(_1596_),
    .B2(_1597_),
    .A2(net614),
    .A1(net1030));
 sg13g2_inv_1 _2054_ (.Y(_0380_),
    .A(net1031));
 sg13g2_xnor2_1 _2055_ (.Y(_1599_),
    .A(net1021),
    .B(_0693_));
 sg13g2_a22oi_1 _2056_ (.Y(_1600_),
    .B1(net584),
    .B2(_1599_),
    .A2(net614),
    .A1(net1021));
 sg13g2_inv_1 _2057_ (.Y(_0381_),
    .A(net1022));
 sg13g2_xor2_1 _2058_ (.B(_0694_),
    .A(net1057),
    .X(_1601_));
 sg13g2_a22oi_1 _2059_ (.Y(_1602_),
    .B1(net584),
    .B2(_1601_),
    .A2(net614),
    .A1(net1057));
 sg13g2_inv_1 _2060_ (.Y(_0382_),
    .A(net1058));
 sg13g2_nand2_1 _2061_ (.Y(_1603_),
    .A(net480),
    .B(net614));
 sg13g2_a21oi_1 _2062_ (.A1(\bp_core.init_counter[8] ),
    .A2(_0694_),
    .Y(_1604_),
    .B1(net480));
 sg13g2_nand2_1 _2063_ (.Y(_1605_),
    .A(_0695_),
    .B(net584));
 sg13g2_o21ai_1 _2064_ (.B1(_1603_),
    .Y(_0383_),
    .A1(_1604_),
    .A2(_1605_));
 sg13g2_xnor2_1 _2065_ (.Y(_1606_),
    .A(net1012),
    .B(_0695_));
 sg13g2_a22oi_1 _2066_ (.Y(_1607_),
    .B1(net584),
    .B2(_1606_),
    .A2(net614),
    .A1(net1012));
 sg13g2_inv_1 _2067_ (.Y(_0384_),
    .A(net1013));
 sg13g2_xor2_1 _2068_ (.B(_0696_),
    .A(net1094),
    .X(_1608_));
 sg13g2_a22oi_1 _2069_ (.Y(_1609_),
    .B1(net584),
    .B2(_1608_),
    .A2(net615),
    .A1(net1094));
 sg13g2_inv_1 _2070_ (.Y(_0385_),
    .A(_1609_));
 sg13g2_a21o_1 _2071_ (.A2(_0696_),
    .A1(\bp_core.init_counter[11] ),
    .B1(net1075),
    .X(_1610_));
 sg13g2_and2_1 _2072_ (.A(_0697_),
    .B(net586),
    .X(_1611_));
 sg13g2_a22oi_1 _2073_ (.Y(_1612_),
    .B1(_1610_),
    .B2(_1611_),
    .A2(net615),
    .A1(net1075));
 sg13g2_inv_1 _2074_ (.Y(_0386_),
    .A(net1076));
 sg13g2_xnor2_1 _2075_ (.Y(_1613_),
    .A(net1049),
    .B(_0697_));
 sg13g2_a22oi_1 _2076_ (.Y(_1614_),
    .B1(net586),
    .B2(_1613_),
    .A2(net615),
    .A1(net1049));
 sg13g2_inv_1 _2077_ (.Y(_0387_),
    .A(net1050));
 sg13g2_xor2_1 _2078_ (.B(_0698_),
    .A(net1051),
    .X(_1615_));
 sg13g2_a22oi_1 _2079_ (.Y(_1616_),
    .B1(net586),
    .B2(_1615_),
    .A2(_1583_),
    .A1(net1051));
 sg13g2_inv_1 _2080_ (.Y(_0388_),
    .A(net1052));
 sg13g2_nand2_1 _2081_ (.Y(_1617_),
    .A(net368),
    .B(_1583_));
 sg13g2_o21ai_1 _2082_ (.B1(_1576_),
    .Y(_1618_),
    .A1(net368),
    .A2(_0699_));
 sg13g2_o21ai_1 _2083_ (.B1(net369),
    .Y(_0389_),
    .A1(_0825_),
    .A2(_1618_));
 sg13g2_nor3_1 _2084_ (.A(net292),
    .B(_0706_),
    .C(_0812_),
    .Y(_1619_));
 sg13g2_a21oi_1 _2085_ (.A1(_0549_),
    .A2(net359),
    .Y(_1620_),
    .B1(_0815_));
 sg13g2_nand2_1 _2086_ (.Y(_1621_),
    .A(_0707_),
    .B(_1620_));
 sg13g2_a21oi_1 _2087_ (.A1(net292),
    .A2(_1621_),
    .Y(_1622_),
    .B1(_1619_));
 sg13g2_inv_1 _2088_ (.Y(_0390_),
    .A(_1622_));
 sg13g2_nor3_1 _2089_ (.A(\bp_core.state[1] ),
    .B(net754),
    .C(net600),
    .Y(_1623_));
 sg13g2_a21oi_1 _2090_ (.A1(_0551_),
    .A2(net600),
    .Y(_0391_),
    .B1(_1623_));
 sg13g2_nand2_1 _2091_ (.Y(_1624_),
    .A(net357),
    .B(_0818_));
 sg13g2_a21oi_1 _2092_ (.A1(_0817_),
    .A2(_1624_),
    .Y(_0392_),
    .B1(_1511_));
 sg13g2_nand2_1 _2093_ (.Y(_1625_),
    .A(net456),
    .B(net716));
 sg13g2_a21oi_1 _2094_ (.A1(net609),
    .A2(_1625_),
    .Y(_0393_),
    .B1(_1516_));
 sg13g2_a21oi_1 _2095_ (.A1(net492),
    .A2(net716),
    .Y(_1626_),
    .B1(_0011_));
 sg13g2_nor2_1 _2096_ (.A(_1522_),
    .B(_1626_),
    .Y(_0394_));
 sg13g2_a21oi_1 _2097_ (.A1(net441),
    .A2(net716),
    .Y(_1627_),
    .B1(_0011_));
 sg13g2_nor2_1 _2098_ (.A(_1527_),
    .B(_1627_),
    .Y(_0395_));
 sg13g2_a21oi_1 _2099_ (.A1(net223),
    .A2(net716),
    .Y(_1628_),
    .B1(_0011_));
 sg13g2_nor2_1 _2100_ (.A(_1532_),
    .B(_1628_),
    .Y(_0396_));
 sg13g2_a21oi_1 _2101_ (.A1(net266),
    .A2(net716),
    .Y(_1629_),
    .B1(_0011_));
 sg13g2_nor2_1 _2102_ (.A(_1538_),
    .B(_1629_),
    .Y(_0397_));
 sg13g2_a21oi_1 _2103_ (.A1(net227),
    .A2(net716),
    .Y(_1630_),
    .B1(_0011_));
 sg13g2_nor2_1 _2104_ (.A(_1543_),
    .B(_1630_),
    .Y(_0398_));
 sg13g2_a21oi_1 _2105_ (.A1(net355),
    .A2(net716),
    .Y(_1631_),
    .B1(_0011_));
 sg13g2_nor2_1 _2106_ (.A(_1547_),
    .B(_1631_),
    .Y(_0399_));
 sg13g2_nor2_1 _2107_ (.A(_0527_),
    .B(net750),
    .Y(_1632_));
 sg13g2_a21oi_1 _2108_ (.A1(\bp_core.init_counter[0] ),
    .A2(net753),
    .Y(_1633_),
    .B1(_1632_));
 sg13g2_nand2_1 _2109_ (.Y(_1634_),
    .A(net219),
    .B(net604));
 sg13g2_o21ai_1 _2110_ (.B1(_1634_),
    .Y(_0400_),
    .A1(net601),
    .A2(_1633_));
 sg13g2_nor2_1 _2111_ (.A(_0528_),
    .B(net754),
    .Y(_1635_));
 sg13g2_a21oi_1 _2112_ (.A1(\bp_core.init_counter[1] ),
    .A2(net753),
    .Y(_1636_),
    .B1(_1635_));
 sg13g2_nand2_1 _2113_ (.Y(_1637_),
    .A(net148),
    .B(net604));
 sg13g2_o21ai_1 _2114_ (.B1(_1637_),
    .Y(_0401_),
    .A1(net605),
    .A2(_1636_));
 sg13g2_nor2_1 _2115_ (.A(_0529_),
    .B(net753),
    .Y(_1638_));
 sg13g2_a21oi_1 _2116_ (.A1(\bp_core.init_counter[2] ),
    .A2(net753),
    .Y(_1639_),
    .B1(_1638_));
 sg13g2_nand2_1 _2117_ (.Y(_1640_),
    .A(net113),
    .B(net604));
 sg13g2_o21ai_1 _2118_ (.B1(_1640_),
    .Y(_0402_),
    .A1(net605),
    .A2(_1639_));
 sg13g2_nor2_1 _2119_ (.A(_0530_),
    .B(net753),
    .Y(_1641_));
 sg13g2_a21oi_1 _2120_ (.A1(\bp_core.init_counter[3] ),
    .A2(net753),
    .Y(_1642_),
    .B1(_1641_));
 sg13g2_nand2_1 _2121_ (.Y(_1643_),
    .A(net152),
    .B(net604));
 sg13g2_o21ai_1 _2122_ (.B1(_1643_),
    .Y(_0403_),
    .A1(net604),
    .A2(_1642_));
 sg13g2_nor2_1 _2123_ (.A(_0531_),
    .B(net754),
    .Y(_1644_));
 sg13g2_a21oi_1 _2124_ (.A1(\bp_core.init_counter[4] ),
    .A2(net753),
    .Y(_1645_),
    .B1(_1644_));
 sg13g2_nand2_1 _2125_ (.Y(_1646_),
    .A(net169),
    .B(net604));
 sg13g2_o21ai_1 _2126_ (.B1(_1646_),
    .Y(_0404_),
    .A1(net603),
    .A2(_1645_));
 sg13g2_nor2_1 _2127_ (.A(_0532_),
    .B(net751),
    .Y(_1647_));
 sg13g2_a21oi_1 _2128_ (.A1(\bp_core.init_counter[5] ),
    .A2(net752),
    .Y(_1648_),
    .B1(_1647_));
 sg13g2_nand2_1 _2129_ (.Y(_1649_),
    .A(net154),
    .B(net604));
 sg13g2_o21ai_1 _2130_ (.B1(_1649_),
    .Y(_0405_),
    .A1(net603),
    .A2(_1648_));
 sg13g2_nor2_1 _2131_ (.A(_0533_),
    .B(net751),
    .Y(_1650_));
 sg13g2_a21oi_1 _2132_ (.A1(\bp_core.init_counter[6] ),
    .A2(net752),
    .Y(_1651_),
    .B1(_1650_));
 sg13g2_nand2_1 _2133_ (.Y(_1652_),
    .A(net120),
    .B(net602));
 sg13g2_o21ai_1 _2134_ (.B1(_1652_),
    .Y(_0406_),
    .A1(net602),
    .A2(_1651_));
 sg13g2_nor2_1 _2135_ (.A(_0534_),
    .B(net751),
    .Y(_1653_));
 sg13g2_a21oi_1 _2136_ (.A1(\bp_core.init_counter[7] ),
    .A2(net751),
    .Y(_1654_),
    .B1(_1653_));
 sg13g2_nand2_1 _2137_ (.Y(_1655_),
    .A(net122),
    .B(net602));
 sg13g2_o21ai_1 _2138_ (.B1(_1655_),
    .Y(_0407_),
    .A1(net602),
    .A2(_1654_));
 sg13g2_nor2_1 _2139_ (.A(_0535_),
    .B(net751),
    .Y(_1656_));
 sg13g2_a21oi_1 _2140_ (.A1(\bp_core.init_counter[8] ),
    .A2(net751),
    .Y(_1657_),
    .B1(_1656_));
 sg13g2_nand2_1 _2141_ (.Y(_1658_),
    .A(net107),
    .B(net602));
 sg13g2_o21ai_1 _2142_ (.B1(_1658_),
    .Y(_0408_),
    .A1(net602),
    .A2(_1657_));
 sg13g2_nor2_1 _2143_ (.A(_0536_),
    .B(net751),
    .Y(_1659_));
 sg13g2_a21oi_1 _2144_ (.A1(\bp_core.init_counter[9] ),
    .A2(net751),
    .Y(_1660_),
    .B1(_1659_));
 sg13g2_nand2_1 _2145_ (.Y(_1661_),
    .A(net192),
    .B(net602));
 sg13g2_o21ai_1 _2146_ (.B1(_1661_),
    .Y(_0409_),
    .A1(net602),
    .A2(_1660_));
 sg13g2_nor2_1 _2147_ (.A(_0554_),
    .B(net755),
    .Y(_1662_));
 sg13g2_a21oi_1 _2148_ (.A1(\bp_core.addr_reg[10] ),
    .A2(net755),
    .Y(_1663_),
    .B1(_1662_));
 sg13g2_nand2_1 _2149_ (.Y(_1664_),
    .A(net177),
    .B(net603));
 sg13g2_o21ai_1 _2150_ (.B1(_1664_),
    .Y(_0410_),
    .A1(net603),
    .A2(_1663_));
 sg13g2_nor2_1 _2151_ (.A(_0538_),
    .B(net754),
    .Y(_1665_));
 sg13g2_a21oi_1 _2152_ (.A1(\bp_core.init_counter[11] ),
    .A2(net752),
    .Y(_1666_),
    .B1(_1665_));
 sg13g2_nand2_1 _2153_ (.Y(_1667_),
    .A(net194),
    .B(net603));
 sg13g2_o21ai_1 _2154_ (.B1(_1667_),
    .Y(_0411_),
    .A1(net603),
    .A2(_1666_));
 sg13g2_nor2_1 _2155_ (.A(_0540_),
    .B(net752),
    .Y(_1668_));
 sg13g2_a21oi_1 _2156_ (.A1(\bp_core.init_counter[12] ),
    .A2(net752),
    .Y(_1669_),
    .B1(_1668_));
 sg13g2_nand2_1 _2157_ (.Y(_1670_),
    .A(net173),
    .B(net603));
 sg13g2_o21ai_1 _2158_ (.B1(_1670_),
    .Y(_0412_),
    .A1(net601),
    .A2(_1669_));
 sg13g2_nor2_1 _2159_ (.A(_0555_),
    .B(_0709_),
    .Y(_1671_));
 sg13g2_a21oi_1 _2160_ (.A1(\bp_core.addr_reg[13] ),
    .A2(_0709_),
    .Y(_1672_),
    .B1(_1671_));
 sg13g2_nand2_1 _2161_ (.Y(_1673_),
    .A(net131),
    .B(net600));
 sg13g2_o21ai_1 _2162_ (.B1(_1673_),
    .Y(_0413_),
    .A1(net601),
    .A2(_1672_));
 sg13g2_nor2_1 _2163_ (.A(_0542_),
    .B(net754),
    .Y(_1674_));
 sg13g2_a21oi_1 _2164_ (.A1(\bp_core.init_counter[14] ),
    .A2(net754),
    .Y(_1675_),
    .B1(_1674_));
 sg13g2_nand2_1 _2165_ (.Y(_1676_),
    .A(net141),
    .B(net600));
 sg13g2_o21ai_1 _2166_ (.B1(_1676_),
    .Y(_0414_),
    .A1(net600),
    .A2(_1675_));
 sg13g2_nor2_1 _2167_ (.A(_0543_),
    .B(net750),
    .Y(_1677_));
 sg13g2_a21oi_1 _2168_ (.A1(\bp_core.init_counter[15] ),
    .A2(net750),
    .Y(_1678_),
    .B1(_1677_));
 sg13g2_nand2_1 _2169_ (.Y(_1679_),
    .A(net171),
    .B(net600));
 sg13g2_o21ai_1 _2170_ (.B1(_1679_),
    .Y(_0415_),
    .A1(net600),
    .A2(_1678_));
 sg13g2_nand2_1 _2171_ (.Y(_1680_),
    .A(net4),
    .B(net652));
 sg13g2_o21ai_1 _2172_ (.B1(_1680_),
    .Y(_0416_),
    .A1(_0666_),
    .A2(net652));
 sg13g2_nand2_1 _2173_ (.Y(_1681_),
    .A(net5),
    .B(net652));
 sg13g2_o21ai_1 _2174_ (.B1(_1681_),
    .Y(_0417_),
    .A1(_0663_),
    .A2(net652));
 sg13g2_nand2_1 _2175_ (.Y(_1682_),
    .A(net6),
    .B(_0813_));
 sg13g2_o21ai_1 _2176_ (.B1(_1682_),
    .Y(_0418_),
    .A1(_0661_),
    .A2(net652));
 sg13g2_nor2_1 _2177_ (.A(net540),
    .B(net652),
    .Y(_1683_));
 sg13g2_a21oi_1 _2178_ (.A1(net7),
    .A2(net652),
    .Y(_0419_),
    .B1(_1683_));
 sg13g2_mux2_1 _2179_ (.A0(net1028),
    .A1(net8),
    .S(net652),
    .X(_0420_));
 sg13g2_or2_1 _2180_ (.X(_0421_),
    .B(_0700_),
    .A(net864));
 sg13g2_a21oi_2 _2181_ (.B1(_1321_),
    .Y(_1684_),
    .A2(_1447_),
    .A1(net733));
 sg13g2_o21ai_1 _2182_ (.B1(net657),
    .Y(_1685_),
    .A1(net730),
    .A2(_0600_));
 sg13g2_mux2_1 _2183_ (.A0(net1137),
    .A1(_1685_),
    .S(_1684_),
    .X(_0422_));
 sg13g2_o21ai_1 _2184_ (.B1(net656),
    .Y(_1686_),
    .A1(net729),
    .A2(_0602_));
 sg13g2_mux2_1 _2185_ (.A0(net1138),
    .A1(_1686_),
    .S(_1684_),
    .X(_0423_));
 sg13g2_o21ai_1 _2186_ (.B1(net655),
    .Y(_1687_),
    .A1(net730),
    .A2(_0604_));
 sg13g2_mux2_1 _2187_ (.A0(net1151),
    .A1(_1687_),
    .S(_1684_),
    .X(_0424_));
 sg13g2_o21ai_1 _2188_ (.B1(net654),
    .Y(_1688_),
    .A1(net729),
    .A2(_0606_));
 sg13g2_mux2_1 _2189_ (.A0(net1156),
    .A1(_1688_),
    .S(_1684_),
    .X(_0425_));
 sg13g2_o21ai_1 _2190_ (.B1(_1333_),
    .Y(_1689_),
    .A1(net736),
    .A2(_0608_));
 sg13g2_mux2_1 _2191_ (.A0(net1179),
    .A1(_1689_),
    .S(_1684_),
    .X(_0426_));
 sg13g2_and2_1 _2192_ (.A(\bp_core.ram_start ),
    .B(spi_cs),
    .X(_1690_));
 sg13g2_nand2_1 _2193_ (.Y(_1691_),
    .A(\bp_core.ram_start ),
    .B(spi_cs));
 sg13g2_nor2_1 _2194_ (.A(net673),
    .B(_1690_),
    .Y(_1692_));
 sg13g2_a22oi_1 _2195_ (.Y(_1693_),
    .B1(net583),
    .B2(net366),
    .A2(_1690_),
    .A1(net219));
 sg13g2_inv_1 _2196_ (.Y(_0427_),
    .A(net367));
 sg13g2_a22oi_1 _2197_ (.Y(_1694_),
    .B1(net581),
    .B2(net305),
    .A2(net672),
    .A1(\spi_ctrl.addr[0] ));
 sg13g2_o21ai_1 _2198_ (.B1(net306),
    .Y(_0428_),
    .A1(_0668_),
    .A2(net612));
 sg13g2_a22oi_1 _2199_ (.Y(_1695_),
    .B1(net581),
    .B2(net303),
    .A2(net671),
    .A1(\spi_ctrl.addr[1] ));
 sg13g2_o21ai_1 _2200_ (.B1(net304),
    .Y(_0429_),
    .A1(_0669_),
    .A2(net611));
 sg13g2_a22oi_1 _2201_ (.Y(_1696_),
    .B1(net581),
    .B2(net313),
    .A2(net672),
    .A1(net303));
 sg13g2_o21ai_1 _2202_ (.B1(_1696_),
    .Y(_0430_),
    .A1(_0670_),
    .A2(net612));
 sg13g2_a22oi_1 _2203_ (.Y(_1697_),
    .B1(net582),
    .B2(net264),
    .A2(net671),
    .A1(\spi_ctrl.addr[3] ));
 sg13g2_o21ai_1 _2204_ (.B1(net265),
    .Y(_0431_),
    .A1(_0671_),
    .A2(net611));
 sg13g2_a22oi_1 _2205_ (.Y(_1698_),
    .B1(net581),
    .B2(net315),
    .A2(net671),
    .A1(net264));
 sg13g2_o21ai_1 _2206_ (.B1(_1698_),
    .Y(_0432_),
    .A1(_0672_),
    .A2(net611));
 sg13g2_a22oi_1 _2207_ (.Y(_1699_),
    .B1(net581),
    .B2(net346),
    .A2(net671),
    .A1(net315));
 sg13g2_o21ai_1 _2208_ (.B1(_1699_),
    .Y(_0433_),
    .A1(_0673_),
    .A2(net611));
 sg13g2_a22oi_1 _2209_ (.Y(_1700_),
    .B1(net581),
    .B2(net316),
    .A2(net671),
    .A1(\spi_ctrl.addr[6] ));
 sg13g2_o21ai_1 _2210_ (.B1(net317),
    .Y(_0434_),
    .A1(_0674_),
    .A2(net611));
 sg13g2_a22oi_1 _2211_ (.Y(_1701_),
    .B1(net582),
    .B2(net362),
    .A2(net671),
    .A1(net316));
 sg13g2_o21ai_1 _2212_ (.B1(_1701_),
    .Y(_0435_),
    .A1(_0675_),
    .A2(net611));
 sg13g2_a22oi_1 _2213_ (.Y(_1702_),
    .B1(net582),
    .B2(net294),
    .A2(net671),
    .A1(\spi_ctrl.addr[8] ));
 sg13g2_o21ai_1 _2214_ (.B1(net295),
    .Y(_0436_),
    .A1(_0676_),
    .A2(net611));
 sg13g2_a22oi_1 _2215_ (.Y(_1703_),
    .B1(net582),
    .B2(net312),
    .A2(net671),
    .A1(net294));
 sg13g2_o21ai_1 _2216_ (.B1(_1703_),
    .Y(_0437_),
    .A1(_0677_),
    .A2(net611));
 sg13g2_a22oi_1 _2217_ (.Y(_1704_),
    .B1(net581),
    .B2(net339),
    .A2(net672),
    .A1(net312));
 sg13g2_o21ai_1 _2218_ (.B1(_1704_),
    .Y(_0438_),
    .A1(_0678_),
    .A2(net612));
 sg13g2_a22oi_1 _2219_ (.Y(_1705_),
    .B1(net581),
    .B2(net378),
    .A2(net672),
    .A1(net339));
 sg13g2_o21ai_1 _2220_ (.B1(_1705_),
    .Y(_0439_),
    .A1(_0679_),
    .A2(net612));
 sg13g2_a22oi_1 _2221_ (.Y(_1706_),
    .B1(net583),
    .B2(net238),
    .A2(net673),
    .A1(\spi_ctrl.addr[12] ));
 sg13g2_o21ai_1 _2222_ (.B1(net239),
    .Y(_0440_),
    .A1(_0680_),
    .A2(net613));
 sg13g2_a22oi_1 _2223_ (.Y(_1707_),
    .B1(net583),
    .B2(net235),
    .A2(net673),
    .A1(\spi_ctrl.addr[13] ));
 sg13g2_o21ai_1 _2224_ (.B1(net236),
    .Y(_0441_),
    .A1(_0681_),
    .A2(net613));
 sg13g2_a22oi_1 _2225_ (.Y(_1708_),
    .B1(net583),
    .B2(net252),
    .A2(net673),
    .A1(net235));
 sg13g2_o21ai_1 _2226_ (.B1(_1708_),
    .Y(_0442_),
    .A1(_0682_),
    .A2(net613));
 sg13g2_o21ai_1 _2227_ (.B1(_1322_),
    .Y(_1709_),
    .A1(_0526_),
    .A2(_1450_));
 sg13g2_o21ai_1 _2228_ (.B1(_1325_),
    .Y(_1710_),
    .A1(net735),
    .A2(_0580_));
 sg13g2_mux2_1 _2229_ (.A0(_1710_),
    .A1(net988),
    .S(_1709_),
    .X(_0443_));
 sg13g2_o21ai_1 _2230_ (.B1(net656),
    .Y(_1711_),
    .A1(net735),
    .A2(_0582_));
 sg13g2_mux2_1 _2231_ (.A0(_1711_),
    .A1(net979),
    .S(_1709_),
    .X(_0444_));
 sg13g2_o21ai_1 _2232_ (.B1(_1329_),
    .Y(_1712_),
    .A1(net735),
    .A2(_0584_));
 sg13g2_mux2_1 _2233_ (.A0(_1712_),
    .A1(net1011),
    .S(_1709_),
    .X(_0445_));
 sg13g2_o21ai_1 _2234_ (.B1(net654),
    .Y(_1713_),
    .A1(net736),
    .A2(_0586_));
 sg13g2_mux2_1 _2235_ (.A0(_1713_),
    .A1(net1037),
    .S(_1709_),
    .X(_0446_));
 sg13g2_o21ai_1 _2236_ (.B1(net653),
    .Y(_1714_),
    .A1(net736),
    .A2(_0588_));
 sg13g2_mux2_1 _2237_ (.A0(_1714_),
    .A1(net1046),
    .S(_1709_),
    .X(_0447_));
 sg13g2_a21oi_2 _2238_ (.B1(_1321_),
    .Y(_1715_),
    .A2(_1445_),
    .A1(net733));
 sg13g2_o21ai_1 _2239_ (.B1(_1325_),
    .Y(_1716_),
    .A1(net735),
    .A2(_0570_));
 sg13g2_mux2_1 _2240_ (.A0(net976),
    .A1(_1716_),
    .S(_1715_),
    .X(_0448_));
 sg13g2_o21ai_1 _2241_ (.B1(net656),
    .Y(_1717_),
    .A1(net735),
    .A2(_0572_));
 sg13g2_mux2_1 _2242_ (.A0(net989),
    .A1(_1717_),
    .S(_1715_),
    .X(_0449_));
 sg13g2_o21ai_1 _2243_ (.B1(net655),
    .Y(_1718_),
    .A1(net735),
    .A2(_0574_));
 sg13g2_mux2_1 _2244_ (.A0(net1029),
    .A1(_1718_),
    .S(_1715_),
    .X(_0450_));
 sg13g2_o21ai_1 _2245_ (.B1(net654),
    .Y(_1719_),
    .A1(net735),
    .A2(_0576_));
 sg13g2_mux2_1 _2246_ (.A0(net1010),
    .A1(_1719_),
    .S(_1715_),
    .X(_0451_));
 sg13g2_o21ai_1 _2247_ (.B1(net653),
    .Y(_1720_),
    .A1(net736),
    .A2(_0578_));
 sg13g2_mux2_1 _2248_ (.A0(net957),
    .A1(_1720_),
    .S(_1715_),
    .X(_0452_));
 sg13g2_a21o_2 _2249_ (.A2(_1452_),
    .A1(net733),
    .B1(_1321_),
    .X(_1721_));
 sg13g2_nand2_1 _2250_ (.Y(_1722_),
    .A(_0526_),
    .B(net433));
 sg13g2_nor2b_1 _2251_ (.A(_1721_),
    .B_N(net657),
    .Y(_1723_));
 sg13g2_a22oi_1 _2252_ (.Y(_0453_),
    .B1(_1722_),
    .B2(_1723_),
    .A2(_1721_),
    .A1(_0667_));
 sg13g2_o21ai_1 _2253_ (.B1(_1327_),
    .Y(_1724_),
    .A1(net737),
    .A2(_0562_));
 sg13g2_mux2_1 _2254_ (.A0(_1724_),
    .A1(net1016),
    .S(_1721_),
    .X(_0454_));
 sg13g2_o21ai_1 _2255_ (.B1(_1329_),
    .Y(_1725_),
    .A1(net736),
    .A2(_0564_));
 sg13g2_mux2_1 _2256_ (.A0(_1725_),
    .A1(net955),
    .S(_1721_),
    .X(_0455_));
 sg13g2_o21ai_1 _2257_ (.B1(net654),
    .Y(_1726_),
    .A1(net735),
    .A2(_0566_));
 sg13g2_mux2_1 _2258_ (.A0(_1726_),
    .A1(net1035),
    .S(_1721_),
    .X(_0456_));
 sg13g2_o21ai_1 _2259_ (.B1(net653),
    .Y(_1727_),
    .A1(net737),
    .A2(_0568_));
 sg13g2_mux2_1 _2260_ (.A0(_1727_),
    .A1(net986),
    .S(_1721_),
    .X(_0457_));
 sg13g2_nor3_1 _2261_ (.A(net549),
    .B(net380),
    .C(spi_cs),
    .Y(_1728_));
 sg13g2_nand2b_1 _2262_ (.Y(_1729_),
    .B(_1728_),
    .A_N(net225));
 sg13g2_nor2_1 _2263_ (.A(net1169),
    .B(_1729_),
    .Y(_1730_));
 sg13g2_nand2_1 _2264_ (.Y(_1731_),
    .A(net1173),
    .B(_1730_));
 sg13g2_inv_1 _2265_ (.Y(_1732_),
    .A(_1731_));
 sg13g2_o21ai_1 _2266_ (.B1(_0521_),
    .Y(_1733_),
    .A1(\bp_core.ram_start ),
    .A2(_0687_));
 sg13g2_a21o_1 _2267_ (.A2(_1732_),
    .A1(\spi_ctrl.fsm_state[1] ),
    .B1(_1733_),
    .X(_1734_));
 sg13g2_nand2_1 _2268_ (.Y(_1735_),
    .A(net380),
    .B(spi_cs));
 sg13g2_a21oi_1 _2269_ (.A1(_1734_),
    .A2(_1735_),
    .Y(_0458_),
    .B1(_0684_));
 sg13g2_nor2_1 _2270_ (.A(_1690_),
    .B(_1728_),
    .Y(_1736_));
 sg13g2_a21oi_1 _2271_ (.A1(\spi_ctrl.fsm_state[1] ),
    .A2(_1732_),
    .Y(_1737_),
    .B1(_1736_));
 sg13g2_a21oi_1 _2272_ (.A1(net549),
    .A2(_1734_),
    .Y(_1738_),
    .B1(_1737_));
 sg13g2_nor2_1 _2273_ (.A(_0684_),
    .B(net550),
    .Y(_0459_));
 sg13g2_o21ai_1 _2274_ (.B1(net838),
    .Y(_1739_),
    .A1(net225),
    .A2(_1737_));
 sg13g2_a21oi_1 _2275_ (.A1(net225),
    .A2(_1728_),
    .Y(_0460_),
    .B1(_1739_));
 sg13g2_nand3_1 _2276_ (.B(net613),
    .C(_1729_),
    .A(net1169),
    .Y(_1740_));
 sg13g2_o21ai_1 _2277_ (.B1(_1740_),
    .Y(_1741_),
    .A1(net1152),
    .A2(_1731_));
 sg13g2_and2_1 _2278_ (.A(net838),
    .B(net1170),
    .X(_0461_));
 sg13g2_nor3_1 _2279_ (.A(net1173),
    .B(_1690_),
    .C(_1730_),
    .Y(_1742_));
 sg13g2_nor3_1 _2280_ (.A(_0684_),
    .B(_1732_),
    .C(net1174),
    .Y(_0462_));
 sg13g2_xor2_1 _2281_ (.B(_1731_),
    .A(net1152),
    .X(_1743_));
 sg13g2_nor2_1 _2282_ (.A(_0684_),
    .B(net1153),
    .Y(_0463_));
 sg13g2_nor2_1 _2283_ (.A(_0551_),
    .B(net613),
    .Y(_1744_));
 sg13g2_nand2_2 _2284_ (.Y(_1745_),
    .A(\bp_core.ram_we ),
    .B(_1690_));
 sg13g2_a21o_1 _2285_ (.A2(net613),
    .A1(net406),
    .B1(net580),
    .X(_0464_));
 sg13g2_nor2_2 _2286_ (.A(net674),
    .B(net579),
    .Y(_1746_));
 sg13g2_nand2_1 _2287_ (.Y(_1747_),
    .A(\spi_ctrl.spi_miso_buf ),
    .B(net675));
 sg13g2_a22oi_1 _2288_ (.Y(_1748_),
    .B1(_1746_),
    .B2(net1070),
    .A2(net580),
    .A1(net357));
 sg13g2_nand2_1 _2289_ (.Y(_0465_),
    .A(_1747_),
    .B(_1748_));
 sg13g2_nand2_1 _2290_ (.Y(_1749_),
    .A(net868),
    .B(_1746_));
 sg13g2_nor2_1 _2291_ (.A(net456),
    .B(_1745_),
    .Y(_1750_));
 sg13g2_a21oi_1 _2292_ (.A1(\bp_core.ram_rdata[0] ),
    .A2(net675),
    .Y(_1751_),
    .B1(net580));
 sg13g2_o21ai_1 _2293_ (.B1(_1749_),
    .Y(_0466_),
    .A1(_1750_),
    .A2(_1751_));
 sg13g2_nand2_1 _2294_ (.Y(_1752_),
    .A(net416),
    .B(_1746_));
 sg13g2_nor2_1 _2295_ (.A(\bp_core.ram_wdata[2] ),
    .B(_1745_),
    .Y(_1753_));
 sg13g2_a21oi_1 _2296_ (.A1(\bp_core.ram_rdata[1] ),
    .A2(net674),
    .Y(_1754_),
    .B1(net579));
 sg13g2_o21ai_1 _2297_ (.B1(_1752_),
    .Y(_0467_),
    .A1(_1753_),
    .A2(_1754_));
 sg13g2_nand2_1 _2298_ (.Y(_1755_),
    .A(net388),
    .B(_1746_));
 sg13g2_nor2_1 _2299_ (.A(\bp_core.ram_wdata[3] ),
    .B(_1745_),
    .Y(_1756_));
 sg13g2_a21oi_1 _2300_ (.A1(\bp_core.ram_rdata[2] ),
    .A2(net675),
    .Y(_1757_),
    .B1(net579));
 sg13g2_o21ai_1 _2301_ (.B1(_1755_),
    .Y(_0468_),
    .A1(_1756_),
    .A2(_1757_));
 sg13g2_nand2_1 _2302_ (.Y(_1758_),
    .A(net223),
    .B(net579));
 sg13g2_nand2b_1 _2303_ (.Y(_1759_),
    .B(net674),
    .A_N(\bp_core.ram_rdata[3] ));
 sg13g2_o21ai_1 _2304_ (.B1(_1759_),
    .Y(_1760_),
    .A1(\bp_core.ram_rdata[4] ),
    .A2(net674));
 sg13g2_o21ai_1 _2305_ (.B1(_1758_),
    .Y(_0469_),
    .A1(net579),
    .A2(_1760_));
 sg13g2_a22oi_1 _2306_ (.Y(_1761_),
    .B1(_1746_),
    .B2(\bp_core.ram_rdata[5] ),
    .A2(net674),
    .A1(\bp_core.ram_rdata[4] ));
 sg13g2_o21ai_1 _2307_ (.B1(_1761_),
    .Y(_0470_),
    .A1(_0683_),
    .A2(_1745_));
 sg13g2_nand2_1 _2308_ (.Y(_1762_),
    .A(net227),
    .B(net579));
 sg13g2_nand2b_1 _2309_ (.Y(_1763_),
    .B(net674),
    .A_N(\bp_core.ram_rdata[5] ));
 sg13g2_o21ai_1 _2310_ (.B1(_1763_),
    .Y(_1764_),
    .A1(\bp_core.ram_rdata[6] ),
    .A2(net674));
 sg13g2_o21ai_1 _2311_ (.B1(_1762_),
    .Y(_0471_),
    .A1(net579),
    .A2(_1764_));
 sg13g2_nand2_1 _2312_ (.Y(_1765_),
    .A(net331),
    .B(net674));
 sg13g2_a22oi_1 _2313_ (.Y(_1766_),
    .B1(_1746_),
    .B2(\bp_core.ram_rdata[7] ),
    .A2(net579),
    .A1(\bp_core.ram_wdata[7] ));
 sg13g2_nand2_1 _2314_ (.Y(_0472_),
    .A(_1765_),
    .B(_1766_));
 sg13g2_mux2_1 _2315_ (.A0(net397),
    .A1(net495),
    .S(net680),
    .X(_0473_));
 sg13g2_mux2_1 _2316_ (.A0(net408),
    .A1(net562),
    .S(net682),
    .X(_0474_));
 sg13g2_mux2_1 _2317_ (.A0(\inter_bp.param_shift_reg[2] ),
    .A1(net490),
    .S(net683),
    .X(_0475_));
 sg13g2_mux2_1 _2318_ (.A0(\inter_bp.param_shift_reg[3] ),
    .A1(net894),
    .S(net682),
    .X(_0476_));
 sg13g2_mux2_1 _2319_ (.A0(\inter_bp.param_shift_reg[4] ),
    .A1(net510),
    .S(net681),
    .X(_0477_));
 sg13g2_mux2_1 _2320_ (.A0(\inter_bp.param_shift_reg[5] ),
    .A1(net553),
    .S(net681),
    .X(_0478_));
 sg13g2_mux2_1 _2321_ (.A0(net493),
    .A1(net514),
    .S(net681),
    .X(_0479_));
 sg13g2_mux2_1 _2322_ (.A0(\inter_bp.param_shift_reg[7] ),
    .A1(net851),
    .S(net681),
    .X(_0480_));
 sg13g2_mux2_1 _2323_ (.A0(\inter_bp.param_shift_reg[8] ),
    .A1(net531),
    .S(net681),
    .X(_0481_));
 sg13g2_mux2_1 _2324_ (.A0(\inter_bp.param_shift_reg[9] ),
    .A1(net860),
    .S(net682),
    .X(_0482_));
 sg13g2_mux2_1 _2325_ (.A0(\inter_bp.param_shift_reg[10] ),
    .A1(net842),
    .S(net681),
    .X(_0483_));
 sg13g2_mux2_1 _2326_ (.A0(\inter_bp.param_shift_reg[11] ),
    .A1(net523),
    .S(net681),
    .X(_0484_));
 sg13g2_mux2_1 _2327_ (.A0(\inter_bp.param_shift_reg[12] ),
    .A1(net470),
    .S(net681),
    .X(_0485_));
 sg13g2_mux2_1 _2328_ (.A0(net484),
    .A1(net565),
    .S(net683),
    .X(_0486_));
 sg13g2_mux2_1 _2329_ (.A0(\inter_bp.param_shift_reg[14] ),
    .A1(net900),
    .S(net683),
    .X(_0487_));
 sg13g2_mux2_1 _2330_ (.A0(\inter_bp.param_shift_reg[15] ),
    .A1(net875),
    .S(net680),
    .X(_0488_));
 sg13g2_mux2_1 _2331_ (.A0(\inter_bp.param_shift_reg[16] ),
    .A1(net845),
    .S(net680),
    .X(_0489_));
 sg13g2_mux2_1 _2332_ (.A0(\inter_bp.param_shift_reg[17] ),
    .A1(net476),
    .S(net676),
    .X(_0490_));
 sg13g2_mux2_1 _2333_ (.A0(net888),
    .A1(net896),
    .S(net680),
    .X(_0491_));
 sg13g2_mux2_1 _2334_ (.A0(\inter_bp.param_shift_reg[19] ),
    .A1(net560),
    .S(net679),
    .X(_0492_));
 sg13g2_mux2_1 _2335_ (.A0(\inter_bp.param_shift_reg[20] ),
    .A1(net478),
    .S(_0944_),
    .X(_0493_));
 sg13g2_mux2_1 _2336_ (.A0(\inter_bp.param_shift_reg[21] ),
    .A1(net488),
    .S(net679),
    .X(_0494_));
 sg13g2_mux2_1 _2337_ (.A0(net444),
    .A1(net509),
    .S(net683),
    .X(_0495_));
 sg13g2_mux2_1 _2338_ (.A0(\inter_bp.param_shift_reg[23] ),
    .A1(net474),
    .S(net676),
    .X(_0496_));
 sg13g2_mux2_1 _2339_ (.A0(\inter_bp.param_shift_reg[24] ),
    .A1(net551),
    .S(net683),
    .X(_0497_));
 sg13g2_mux2_1 _2340_ (.A0(net429),
    .A1(net473),
    .S(net676),
    .X(_0498_));
 sg13g2_mux2_1 _2341_ (.A0(net498),
    .A1(net870),
    .S(net683),
    .X(_0499_));
 sg13g2_mux2_1 _2342_ (.A0(net451),
    .A1(net472),
    .S(net676),
    .X(_0500_));
 sg13g2_mux2_1 _2343_ (.A0(\inter_bp.param_shift_reg[28] ),
    .A1(net518),
    .S(net683),
    .X(_0501_));
 sg13g2_mux2_1 _2344_ (.A0(\inter_bp.param_shift_reg[29] ),
    .A1(net527),
    .S(net676),
    .X(_0502_));
 sg13g2_mux2_1 _2345_ (.A0(net849),
    .A1(net859),
    .S(net680),
    .X(_0503_));
 sg13g2_mux2_1 _2346_ (.A0(net427),
    .A1(net536),
    .S(net676),
    .X(_0504_));
 sg13g2_mux2_1 _2347_ (.A0(\inter_bp.param_shift_reg[32] ),
    .A1(net464),
    .S(net680),
    .X(_0505_));
 sg13g2_mux2_1 _2348_ (.A0(\inter_bp.param_shift_reg[33] ),
    .A1(net468),
    .S(net676),
    .X(_0506_));
 sg13g2_mux2_1 _2349_ (.A0(\inter_bp.param_shift_reg[34] ),
    .A1(net500),
    .S(net680),
    .X(_0507_));
 sg13g2_mux2_1 _2350_ (.A0(\inter_bp.param_shift_reg[35] ),
    .A1(net507),
    .S(net676),
    .X(_0508_));
 sg13g2_mux2_1 _2351_ (.A0(\inter_bp.param_shift_reg[36] ),
    .A1(net466),
    .S(net679),
    .X(_0509_));
 sg13g2_mux2_1 _2352_ (.A0(\inter_bp.param_shift_reg[37] ),
    .A1(net546),
    .S(net677),
    .X(_0510_));
 sg13g2_mux2_1 _2353_ (.A0(net462),
    .A1(net545),
    .S(net678),
    .X(_0511_));
 sg13g2_mux2_1 _2354_ (.A0(\inter_bp.param_shift_reg[39] ),
    .A1(net543),
    .S(net677),
    .X(_0512_));
 sg13g2_mux2_1 _2355_ (.A0(\inter_bp.param_shift_reg[40] ),
    .A1(net883),
    .S(net678),
    .X(_0513_));
 sg13g2_mux2_1 _2356_ (.A0(net349),
    .A1(net885),
    .S(net677),
    .X(_0514_));
 sg13g2_mux2_1 _2357_ (.A0(\inter_bp.param_shift_reg[42] ),
    .A1(net873),
    .S(net678),
    .X(_0515_));
 sg13g2_mux2_1 _2358_ (.A0(\inter_bp.param_shift_reg[43] ),
    .A1(net537),
    .S(net677),
    .X(_0516_));
 sg13g2_mux2_1 _2359_ (.A0(\inter_bp.param_shift_reg[44] ),
    .A1(net496),
    .S(net678),
    .X(_0517_));
 sg13g2_mux2_1 _2360_ (.A0(\inter_bp.param_shift_reg[45] ),
    .A1(net558),
    .S(net677),
    .X(_0518_));
 sg13g2_mux2_1 _2361_ (.A0(\inter_bp.param_shift_reg[46] ),
    .A1(net502),
    .S(net677),
    .X(_0519_));
 sg13g2_mux2_1 _2362_ (.A0(\inter_bp.param_shift_reg[47] ),
    .A1(net541),
    .S(net677),
    .X(_0520_));
 sg13g2_inv_1 _2403__2 (.Y(net56),
    .A(clknet_1_0__leaf_clk));
 sg13g2_inv_1 _2364_ (.Y(_0521_),
    .A(net380));
 sg13g2_inv_1 _2365_ (.Y(_0522_),
    .A(_0100_));
 sg13g2_inv_1 _2366_ (.Y(_0523_),
    .A(_0099_));
 sg13g2_inv_4 _2367_ (.A(net1149),
    .Y(_0524_));
 sg13g2_inv_1 _2368_ (.Y(_0525_),
    .A(net756));
 sg13g2_inv_4 _2369_ (.A(net733),
    .Y(_0526_));
 sg13g2_inv_1 _2370_ (.Y(_0527_),
    .A(net1134));
 sg13g2_inv_1 _2371_ (.Y(_0528_),
    .A(net446));
 sg13g2_inv_1 _2372_ (.Y(_0529_),
    .A(net333));
 sg13g2_inv_4 _2373_ (.A(net1106),
    .Y(_0530_));
 sg13g2_inv_2 _2374_ (.Y(_0531_),
    .A(net371));
 sg13g2_inv_1 _2375_ (.Y(_0532_),
    .A(net1157));
 sg13g2_inv_1 _2376_ (.Y(_0533_),
    .A(net1119));
 sg13g2_inv_2 _2377_ (.Y(_0534_),
    .A(net1130));
 sg13g2_inv_2 _2378_ (.Y(_0535_),
    .A(net1118));
 sg13g2_inv_2 _2379_ (.Y(_0536_),
    .A(net1055));
 sg13g2_inv_1 _2380_ (.Y(_0537_),
    .A(net1061));
 sg13g2_inv_2 _2381_ (.Y(_0538_),
    .A(net1115));
 sg13g2_inv_2 _2382_ (.Y(_0539_),
    .A(\bp_core.bp_stride_out[11] ));
 sg13g2_inv_2 _2383_ (.Y(_0540_),
    .A(net1127));
 sg13g2_inv_1 _2384_ (.Y(_0541_),
    .A(net1126));
 sg13g2_inv_2 _2385_ (.Y(_0542_),
    .A(net1133));
 sg13g2_inv_2 _2386_ (.Y(_0543_),
    .A(net1129));
 sg13g2_inv_1 _2387_ (.Y(_0544_),
    .A(net1093));
 sg13g2_inv_1 _2388_ (.Y(_0545_),
    .A(net932));
 sg13g2_inv_1 _2389_ (.Y(_0546_),
    .A(net1120));
 sg13g2_inv_1 _2390_ (.Y(_0547_),
    .A(net722));
 sg13g2_inv_1 _2391_ (.Y(_0548_),
    .A(net1132));
 sg13g2_inv_1 _2392_ (.Y(_0549_),
    .A(net1110));
 sg13g2_inv_1 _2393_ (.Y(_0550_),
    .A(net292));
 sg13g2_inv_1 _2394_ (.Y(_0551_),
    .A(net879));
 sg13g2_inv_1 _2395_ (.Y(_0552_),
    .A(net10));
 sg13g2_inv_1 _2396_ (.Y(_0553_),
    .A(net968));
 sg13g2_inv_1 _2397_ (.Y(_0554_),
    .A(net1012));
 sg13g2_inv_1 _2398_ (.Y(_0555_),
    .A(net1049));
 sg13g2_inv_1 _2399_ (.Y(_0556_),
    .A(net198));
 sg13g2_inv_1 _2400_ (.Y(_0557_),
    .A(net1063));
 sg13g2_inv_1 _2401_ (.Y(_0558_),
    .A(net996));
 sg13g2_inv_1 _2402_ (.Y(_0559_),
    .A(net229));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_inv_1 _2404_ (.Y(_0560_),
    .A(net353));
 sg13g2_inv_1 _2405_ (.Y(_0561_),
    .A(net394));
 sg13g2_inv_2 _2406_ (.Y(_0562_),
    .A(net902));
 sg13g2_inv_1 _2407_ (.Y(_0563_),
    .A(net408));
 sg13g2_inv_1 _2408_ (.Y(_0564_),
    .A(net991));
 sg13g2_inv_1 _2409_ (.Y(_0565_),
    .A(net926));
 sg13g2_inv_2 _2410_ (.Y(_0566_),
    .A(net994));
 sg13g2_inv_1 _2411_ (.Y(_0567_),
    .A(net904));
 sg13g2_inv_1 _2412_ (.Y(_0568_),
    .A(net931));
 sg13g2_inv_1 _2413_ (.Y(_0569_),
    .A(net534));
 sg13g2_inv_1 _2414_ (.Y(_0570_),
    .A(net950));
 sg13g2_inv_1 _2415_ (.Y(_0571_),
    .A(net927));
 sg13g2_inv_1 _2416_ (.Y(_0572_),
    .A(net909));
 sg13g2_inv_1 _2417_ (.Y(_0573_),
    .A(net493));
 sg13g2_inv_1 _2418_ (.Y(_0574_),
    .A(net999));
 sg13g2_inv_1 _2419_ (.Y(_0575_),
    .A(net907));
 sg13g2_inv_1 _2420_ (.Y(_0576_),
    .A(net995));
 sg13g2_inv_1 _2421_ (.Y(_0577_),
    .A(net934));
 sg13g2_inv_2 _2422_ (.Y(_0578_),
    .A(net983));
 sg13g2_inv_1 _2423_ (.Y(_0579_),
    .A(net920));
 sg13g2_inv_1 _2424_ (.Y(_0580_),
    .A(net966));
 sg13g2_inv_1 _2425_ (.Y(_0581_),
    .A(net891));
 sg13g2_inv_1 _2426_ (.Y(_0582_),
    .A(net936));
 sg13g2_inv_1 _2427_ (.Y(_0583_),
    .A(net533));
 sg13g2_inv_1 _2428_ (.Y(_0584_),
    .A(net937));
 sg13g2_inv_1 _2429_ (.Y(_0585_),
    .A(net853));
 sg13g2_inv_1 _2430_ (.Y(_0586_),
    .A(net970));
 sg13g2_inv_1 _2431_ (.Y(_0587_),
    .A(net484));
 sg13g2_inv_1 _2432_ (.Y(_0588_),
    .A(net1018));
 sg13g2_inv_1 _2433_ (.Y(_0589_),
    .A(net1004));
 sg13g2_inv_1 _2434_ (.Y(_0590_),
    .A(net1043));
 sg13g2_inv_1 _2435_ (.Y(_0591_),
    .A(net1005));
 sg13g2_inv_1 _2436_ (.Y(_0592_),
    .A(\bp_addr_in[16] ));
 sg13g2_inv_1 _2437_ (.Y(_0593_),
    .A(net940));
 sg13g2_inv_1 _2438_ (.Y(_0594_),
    .A(net911));
 sg13g2_inv_1 _2439_ (.Y(_0595_),
    .A(net529));
 sg13g2_inv_1 _2440_ (.Y(_0596_),
    .A(\bp_addr_in[18] ));
 sg13g2_inv_1 _2441_ (.Y(_0597_),
    .A(net888));
 sg13g2_inv_1 _2442_ (.Y(_0598_),
    .A(net984));
 sg13g2_inv_1 _2443_ (.Y(_0599_),
    .A(net882));
 sg13g2_inv_1 _2444_ (.Y(_0600_),
    .A(net1014));
 sg13g2_inv_1 _2445_ (.Y(_0601_),
    .A(net942));
 sg13g2_inv_2 _2446_ (.Y(_0602_),
    .A(\bp_core.bp_stride_in[1] ));
 sg13g2_inv_1 _2447_ (.Y(_0603_),
    .A(net856));
 sg13g2_inv_1 _2448_ (.Y(_0604_),
    .A(net563));
 sg13g2_inv_1 _2449_ (.Y(_0605_),
    .A(net444));
 sg13g2_inv_2 _2450_ (.Y(_0606_),
    .A(net982));
 sg13g2_inv_1 _2451_ (.Y(_0607_),
    .A(net935));
 sg13g2_inv_1 _2452_ (.Y(_0608_),
    .A(net903));
 sg13g2_inv_1 _2453_ (.Y(_0609_),
    .A(net881));
 sg13g2_inv_2 _2454_ (.Y(_0610_),
    .A(net548));
 sg13g2_inv_1 _2455_ (.Y(_0611_),
    .A(net429));
 sg13g2_inv_1 _2456_ (.Y(_0612_),
    .A(\bp_core.bp_stride_in[6] ));
 sg13g2_inv_1 _2457_ (.Y(_0613_),
    .A(net498));
 sg13g2_inv_2 _2458_ (.Y(_0614_),
    .A(net951));
 sg13g2_inv_1 _2459_ (.Y(_0615_),
    .A(net451));
 sg13g2_inv_1 _2460_ (.Y(_0616_),
    .A(net947));
 sg13g2_inv_1 _2461_ (.Y(_0617_),
    .A(net525));
 sg13g2_inv_2 _2462_ (.Y(_0618_),
    .A(net1165));
 sg13g2_inv_1 _2463_ (.Y(_0619_),
    .A(net961));
 sg13g2_inv_1 _2464_ (.Y(_0620_),
    .A(net906));
 sg13g2_inv_1 _2465_ (.Y(_0621_),
    .A(net849));
 sg13g2_inv_1 _2466_ (.Y(_0622_),
    .A(net925));
 sg13g2_inv_1 _2467_ (.Y(_0623_),
    .A(net866));
 sg13g2_inv_2 _2468_ (.Y(_0624_),
    .A(net954));
 sg13g2_inv_1 _2469_ (.Y(_0625_),
    .A(net898));
 sg13g2_inv_1 _2470_ (.Y(_0626_),
    .A(net949));
 sg13g2_inv_1 _2471_ (.Y(_0627_),
    .A(net921));
 sg13g2_inv_2 _2472_ (.Y(_0628_),
    .A(net977));
 sg13g2_inv_1 _2473_ (.Y(_0629_),
    .A(net912));
 sg13g2_inv_1 _2474_ (.Y(_0630_),
    .A(net844));
 sg13g2_inv_1 _2475_ (.Y(_0631_),
    .A(net515));
 sg13g2_inv_1 _2476_ (.Y(_0632_),
    .A(net1006));
 sg13g2_inv_1 _2477_ (.Y(_0633_),
    .A(net948));
 sg13g2_inv_1 _2478_ (.Y(_0634_),
    .A(net928));
 sg13g2_inv_1 _2479_ (.Y(_0635_),
    .A(net462));
 sg13g2_inv_2 _2480_ (.Y(_0636_),
    .A(net967));
 sg13g2_inv_1 _2481_ (.Y(_0637_),
    .A(net939));
 sg13g2_inv_1 _2482_ (.Y(_0638_),
    .A(\bp_core.bp_lambda_in[0] ));
 sg13g2_inv_1 _2483_ (.Y(_0639_),
    .A(net945));
 sg13g2_inv_1 _2484_ (.Y(_0640_),
    .A(net978));
 sg13g2_inv_1 _2485_ (.Y(_0641_),
    .A(net971));
 sg13g2_inv_1 _2486_ (.Y(_0642_),
    .A(\bp_core.bp_lambda_in[3] ));
 sg13g2_inv_1 _2487_ (.Y(_0643_),
    .A(net862));
 sg13g2_inv_1 _2488_ (.Y(_0644_),
    .A(net938));
 sg13g2_inv_1 _2489_ (.Y(_0645_),
    .A(net917));
 sg13g2_inv_2 _2490_ (.Y(_0646_),
    .A(\bp_core.bp_lambda_in[5] ));
 sg13g2_inv_1 _2491_ (.Y(_0647_),
    .A(net886));
 sg13g2_inv_2 _2492_ (.Y(_0648_),
    .A(net1143));
 sg13g2_inv_1 _2493_ (.Y(_0649_),
    .A(net992));
 sg13g2_inv_2 _2494_ (.Y(_0650_),
    .A(net919));
 sg13g2_inv_1 _2495_ (.Y(_0651_),
    .A(net910));
 sg13g2_inv_1 _2496_ (.Y(_0652_),
    .A(\bp_core.bp_lambda_out[1] ));
 sg13g2_inv_1 _2497_ (.Y(_0653_),
    .A(net344));
 sg13g2_inv_1 _2498_ (.Y(_0654_),
    .A(net164));
 sg13g2_inv_1 _2499_ (.Y(_0655_),
    .A(net342));
 sg13g2_inv_1 _2500_ (.Y(_0656_),
    .A(net384));
 sg13g2_inv_1 _2501_ (.Y(_0657_),
    .A(net341));
 sg13g2_inv_1 _2502_ (.Y(_0658_),
    .A(net360));
 sg13g2_inv_1 _2503_ (.Y(_0659_),
    .A(net347));
 sg13g2_inv_1 _2504_ (.Y(_0660_),
    .A(net373));
 sg13g2_inv_1 _2505_ (.Y(_0661_),
    .A(net516));
 sg13g2_inv_1 _2506_ (.Y(_0662_),
    .A(net364));
 sg13g2_inv_1 _2507_ (.Y(_0663_),
    .A(net453));
 sg13g2_inv_1 _2508_ (.Y(_0664_),
    .A(net412));
 sg13g2_inv_1 _2509_ (.Y(_0665_),
    .A(net250));
 sg13g2_inv_1 _2510_ (.Y(_0666_),
    .A(net335));
 sg13g2_inv_2 _2511_ (.Y(_0667_),
    .A(\bp_core.params_addr[0] ));
 sg13g2_inv_1 _2512_ (.Y(_0668_),
    .A(net148));
 sg13g2_inv_1 _2513_ (.Y(_0669_),
    .A(net113));
 sg13g2_inv_1 _2514_ (.Y(_0670_),
    .A(net152));
 sg13g2_inv_1 _2515_ (.Y(_0671_),
    .A(net169));
 sg13g2_inv_1 _2516_ (.Y(_0672_),
    .A(net154));
 sg13g2_inv_1 _2517_ (.Y(_0673_),
    .A(net120));
 sg13g2_inv_1 _2518_ (.Y(_0674_),
    .A(net122));
 sg13g2_inv_1 _2519_ (.Y(_0675_),
    .A(net107));
 sg13g2_inv_1 _2520_ (.Y(_0676_),
    .A(net192));
 sg13g2_inv_1 _2521_ (.Y(_0677_),
    .A(net177));
 sg13g2_inv_1 _2522_ (.Y(_0678_),
    .A(net194));
 sg13g2_inv_1 _2523_ (.Y(_0679_),
    .A(net173));
 sg13g2_inv_1 _2524_ (.Y(_0680_),
    .A(net131));
 sg13g2_inv_1 _2525_ (.Y(_0681_),
    .A(net141));
 sg13g2_inv_1 _2526_ (.Y(_0682_),
    .A(net171));
 sg13g2_inv_1 _2527_ (.Y(_0683_),
    .A(net266));
 sg13g2_inv_2 _2528_ (.Y(\bp_core.params_module.state[0] ),
    .A(net77));
 sg13g2_inv_2 _2529_ (.Y(_0684_),
    .A(net838));
 sg13g2_nor2b_2 _2530_ (.A(net2),
    .B_N(net1),
    .Y(_0685_));
 sg13g2_nand2b_2 _2531_ (.Y(_0686_),
    .B(net1),
    .A_N(net2));
 sg13g2_or2_1 _2532_ (.X(_0687_),
    .B(\spi_ctrl.fsm_state[0] ),
    .A(\spi_ctrl.fsm_state[1] ));
 sg13g2_inv_4 _2533_ (.A(_0687_),
    .Y(spi_cs));
 sg13g2_nor2_1 _2534_ (.A(_0686_),
    .B(_0687_),
    .Y(_0688_));
 sg13g2_nand2_1 _2535_ (.Y(_0689_),
    .A(net1042),
    .B(_0688_));
 sg13g2_nand3_1 _2536_ (.B(\bp_core.init_counter[0] ),
    .C(net1053),
    .A(\bp_core.init_counter[1] ),
    .Y(_0690_));
 sg13g2_and4_1 _2537_ (.A(\bp_core.init_counter[1] ),
    .B(\bp_core.init_counter[0] ),
    .C(net1033),
    .D(\bp_core.init_counter[2] ),
    .X(_0691_));
 sg13g2_and2_1 _2538_ (.A(net1044),
    .B(_0691_),
    .X(_0692_));
 sg13g2_nand3_1 _2539_ (.B(net1030),
    .C(_0692_),
    .A(\bp_core.init_counter[5] ),
    .Y(_0693_));
 sg13g2_and4_1 _2540_ (.A(\bp_core.init_counter[5] ),
    .B(net1021),
    .C(net1030),
    .D(_0692_),
    .X(_0694_));
 sg13g2_nand3_1 _2541_ (.B(\bp_core.init_counter[8] ),
    .C(_0694_),
    .A(net480),
    .Y(_0695_));
 sg13g2_nor2_1 _2542_ (.A(_0554_),
    .B(_0695_),
    .Y(_0696_));
 sg13g2_nand3_1 _2543_ (.B(net1075),
    .C(_0696_),
    .A(\bp_core.init_counter[11] ),
    .Y(_0697_));
 sg13g2_nor2_1 _2544_ (.A(_0555_),
    .B(_0697_),
    .Y(_0698_));
 sg13g2_and2_1 _2545_ (.A(net1051),
    .B(_0698_),
    .X(_0699_));
 sg13g2_and4_1 _2546_ (.A(net1042),
    .B(net368),
    .C(_0688_),
    .D(_0699_),
    .X(_0700_));
 sg13g2_nand2_1 _2547_ (.Y(_0701_),
    .A(\bp_core.state[4] ),
    .B(net241));
 sg13g2_nor3_1 _2548_ (.A(net943),
    .B(net1166),
    .C(net963),
    .Y(_0702_));
 sg13g2_nor2_1 _2549_ (.A(net505),
    .B(net929),
    .Y(_0703_));
 sg13g2_nor4_1 _2550_ (.A(net722),
    .B(net1132),
    .C(net505),
    .D(net929),
    .Y(_0704_));
 sg13g2_a22oi_1 _2551_ (.Y(_0705_),
    .B1(_0702_),
    .B2(_0704_),
    .A2(net242),
    .A1(_0686_));
 sg13g2_nor2b_2 _2552_ (.A(net359),
    .B_N(net864),
    .Y(_0706_));
 sg13g2_nor2_1 _2553_ (.A(_0686_),
    .B(_0706_),
    .Y(_0707_));
 sg13g2_nor2_1 _2554_ (.A(net215),
    .B(net1042),
    .Y(_0708_));
 sg13g2_nor2b_2 _2555_ (.A(net1),
    .B_N(net2),
    .Y(_0709_));
 sg13g2_nand2b_2 _2556_ (.Y(_0710_),
    .B(net2),
    .A_N(net1));
 sg13g2_nor3_1 _2557_ (.A(net1110),
    .B(net310),
    .C(net749),
    .Y(_0711_));
 sg13g2_a21oi_1 _2558_ (.A1(_0708_),
    .A2(_0711_),
    .Y(_0712_),
    .B1(_0707_));
 sg13g2_nor2_1 _2559_ (.A(net359),
    .B(net749),
    .Y(_0713_));
 sg13g2_nor4_1 _2560_ (.A(net756),
    .B(net1140),
    .C(net359),
    .D(net750),
    .Y(_0714_));
 sg13g2_nor4_1 _2561_ (.A(_0700_),
    .B(_0705_),
    .C(_0712_),
    .D(_0714_),
    .Y(_0104_));
 sg13g2_nor3_1 _2562_ (.A(net1125),
    .B(net922),
    .C(net77),
    .Y(_0715_));
 sg13g2_nor2_1 _2563_ (.A(\bp_core.params_module.counter[2] ),
    .B(net738),
    .Y(_0716_));
 sg13g2_nand2_2 _2564_ (.Y(_0717_),
    .A(\bp_core.params_module.counter[3] ),
    .B(_0716_));
 sg13g2_nor2_2 _2565_ (.A(\bp_core.params_module.counter[0] ),
    .B(_0717_),
    .Y(_0718_));
 sg13g2_o21ai_1 _2566_ (.B1(net1097),
    .Y(_0719_),
    .A1(\bp_core.params_module.counter[0] ),
    .A2(_0717_));
 sg13g2_nor2_2 _2567_ (.A(_0524_),
    .B(_0717_),
    .Y(_0720_));
 sg13g2_nand2_1 _2568_ (.Y(_0721_),
    .A(net756),
    .B(net733));
 sg13g2_nor2_1 _2569_ (.A(_0720_),
    .B(_0721_),
    .Y(_0722_));
 sg13g2_nor2_1 _2570_ (.A(net59),
    .B(_0722_),
    .Y(_0723_));
 sg13g2_nor2_1 _2571_ (.A(net1098),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_nor2_1 _2572_ (.A(_0715_),
    .B(_0724_),
    .Y(_0103_));
 sg13g2_nand2b_1 _2573_ (.Y(_0725_),
    .B(net943),
    .A_N(net241));
 sg13g2_nor3_1 _2574_ (.A(\bp_core.addr_reg[17] ),
    .B(\bp_core.addr_reg[16] ),
    .C(\bp_core.addr_reg[18] ),
    .Y(_0726_));
 sg13g2_nor2b_1 _2575_ (.A(net1092),
    .B_N(_0726_),
    .Y(_0727_));
 sg13g2_inv_1 _2576_ (.Y(_0728_),
    .A(_0727_));
 sg13g2_nand2_1 _2577_ (.Y(_0729_),
    .A(\bp_core.addr_reg[1] ),
    .B(\bp_core.bp_stride_out[1] ));
 sg13g2_nand2_2 _2578_ (.Y(_0730_),
    .A(net1134),
    .B(net1137));
 sg13g2_xnor2_1 _2579_ (.Y(_0731_),
    .A(net1163),
    .B(net1138));
 sg13g2_o21ai_1 _2580_ (.B1(_0729_),
    .Y(_0732_),
    .A1(_0730_),
    .A2(_0731_));
 sg13g2_nand2_1 _2581_ (.Y(_0733_),
    .A(\bp_core.addr_reg[3] ),
    .B(\bp_core.bp_stride_out[3] ));
 sg13g2_nor2_1 _2582_ (.A(\bp_core.addr_reg[3] ),
    .B(\bp_core.bp_stride_out[3] ),
    .Y(_0734_));
 sg13g2_xnor2_1 _2583_ (.Y(_0735_),
    .A(\bp_core.addr_reg[3] ),
    .B(\bp_core.bp_stride_out[3] ));
 sg13g2_nand2_1 _2584_ (.Y(_0736_),
    .A(net333),
    .B(\bp_core.bp_stride_out[2] ));
 sg13g2_xnor2_1 _2585_ (.Y(_0737_),
    .A(net1141),
    .B(\bp_core.bp_stride_out[2] ));
 sg13g2_nor2_1 _2586_ (.A(_0735_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_o21ai_1 _2587_ (.B1(_0733_),
    .Y(_0739_),
    .A1(_0734_),
    .A2(_0736_));
 sg13g2_a21o_2 _2588_ (.A2(_0738_),
    .A1(_0732_),
    .B1(_0739_),
    .X(_0740_));
 sg13g2_nor2_1 _2589_ (.A(\bp_core.addr_reg[7] ),
    .B(\bp_core.bp_stride_out[7] ),
    .Y(_0741_));
 sg13g2_xnor2_1 _2590_ (.Y(_0742_),
    .A(\bp_core.addr_reg[7] ),
    .B(\bp_core.bp_stride_out[7] ));
 sg13g2_nand2_1 _2591_ (.Y(_0743_),
    .A(net1119),
    .B(\bp_core.bp_stride_out[6] ));
 sg13g2_xor2_1 _2592_ (.B(\bp_core.bp_stride_out[6] ),
    .A(\bp_core.addr_reg[6] ),
    .X(_0744_));
 sg13g2_nand2b_1 _2593_ (.Y(_0745_),
    .B(_0744_),
    .A_N(_0742_));
 sg13g2_nor2_1 _2594_ (.A(\bp_core.addr_reg[5] ),
    .B(\bp_core.bp_stride_out[5] ),
    .Y(_0746_));
 sg13g2_xnor2_1 _2595_ (.Y(_0747_),
    .A(\bp_core.addr_reg[5] ),
    .B(\bp_core.bp_stride_out[5] ));
 sg13g2_nand2_1 _2596_ (.Y(_0748_),
    .A(net371),
    .B(net1183));
 sg13g2_xnor2_1 _2597_ (.Y(_0749_),
    .A(\bp_core.addr_reg[4] ),
    .B(\bp_core.bp_stride_out[4] ));
 sg13g2_nor3_1 _2598_ (.A(_0745_),
    .B(_0747_),
    .C(_0749_),
    .Y(_0750_));
 sg13g2_a22oi_1 _2599_ (.Y(_0751_),
    .B1(\bp_core.addr_reg[5] ),
    .B2(\bp_core.bp_stride_out[5] ),
    .A2(\bp_core.bp_stride_out[4] ),
    .A1(\bp_core.addr_reg[4] ));
 sg13g2_or2_1 _2600_ (.X(_0752_),
    .B(_0751_),
    .A(_0746_));
 sg13g2_a22oi_1 _2601_ (.Y(_0753_),
    .B1(\bp_core.addr_reg[7] ),
    .B2(\bp_core.bp_stride_out[7] ),
    .A2(\bp_core.bp_stride_out[6] ),
    .A1(\bp_core.addr_reg[6] ));
 sg13g2_or2_1 _2602_ (.X(_0754_),
    .B(_0753_),
    .A(_0741_));
 sg13g2_o21ai_1 _2603_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0745_),
    .A2(_0752_));
 sg13g2_a21oi_1 _2604_ (.A1(_0740_),
    .A2(_0750_),
    .Y(_0756_),
    .B1(_0755_));
 sg13g2_a21o_2 _2605_ (.A2(_0750_),
    .A1(_0740_),
    .B1(_0755_),
    .X(_0757_));
 sg13g2_and2_1 _2606_ (.A(\bp_core.addr_reg[15] ),
    .B(\bp_core.bp_stride_out[15] ),
    .X(_0758_));
 sg13g2_or2_1 _2607_ (.X(_0759_),
    .B(\bp_core.bp_stride_out[15] ),
    .A(\bp_core.addr_reg[15] ));
 sg13g2_nor2b_2 _2608_ (.A(_0758_),
    .B_N(_0759_),
    .Y(_0760_));
 sg13g2_and2_1 _2609_ (.A(\bp_core.addr_reg[14] ),
    .B(\bp_core.bp_stride_out[14] ),
    .X(_0761_));
 sg13g2_xnor2_1 _2610_ (.Y(_0762_),
    .A(\bp_core.addr_reg[14] ),
    .B(\bp_core.bp_stride_out[14] ));
 sg13g2_inv_1 _2611_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_and2_1 _2612_ (.A(_0760_),
    .B(_0763_),
    .X(_0764_));
 sg13g2_nand2_1 _2613_ (.Y(_0765_),
    .A(\bp_core.addr_reg[13] ),
    .B(\bp_core.bp_stride_out[13] ));
 sg13g2_nor2_1 _2614_ (.A(\bp_core.addr_reg[13] ),
    .B(\bp_core.bp_stride_out[13] ),
    .Y(_0766_));
 sg13g2_xor2_1 _2615_ (.B(net1184),
    .A(\bp_core.addr_reg[13] ),
    .X(_0767_));
 sg13g2_and2_1 _2616_ (.A(\bp_core.addr_reg[12] ),
    .B(\bp_core.bp_stride_out[12] ),
    .X(_0768_));
 sg13g2_nand2_1 _2617_ (.Y(_0769_),
    .A(\bp_core.addr_reg[12] ),
    .B(\bp_core.bp_stride_out[12] ));
 sg13g2_xor2_1 _2618_ (.B(\bp_core.bp_stride_out[12] ),
    .A(\bp_core.addr_reg[12] ),
    .X(_0770_));
 sg13g2_nand4_1 _2619_ (.B(_0763_),
    .C(_0767_),
    .A(_0760_),
    .Y(_0771_),
    .D(_0770_));
 sg13g2_xnor2_1 _2620_ (.Y(_0772_),
    .A(\bp_core.addr_reg[11] ),
    .B(\bp_core.bp_stride_out[11] ));
 sg13g2_nand2_1 _2621_ (.Y(_0773_),
    .A(\bp_core.addr_reg[10] ),
    .B(\bp_core.bp_stride_out[10] ));
 sg13g2_xnor2_1 _2622_ (.Y(_0774_),
    .A(\bp_core.addr_reg[10] ),
    .B(\bp_core.bp_stride_out[10] ));
 sg13g2_nor2_1 _2623_ (.A(_0772_),
    .B(_0774_),
    .Y(_0775_));
 sg13g2_and2_1 _2624_ (.A(\bp_core.addr_reg[8] ),
    .B(\bp_core.bp_stride_out[8] ),
    .X(_0776_));
 sg13g2_nand2_1 _2625_ (.Y(_0777_),
    .A(\bp_core.addr_reg[8] ),
    .B(\bp_core.bp_stride_out[8] ));
 sg13g2_xor2_1 _2626_ (.B(\bp_core.bp_stride_out[8] ),
    .A(\bp_core.addr_reg[8] ),
    .X(_0778_));
 sg13g2_nand2_1 _2627_ (.Y(_0779_),
    .A(\bp_core.addr_reg[9] ),
    .B(\bp_core.bp_stride_out[9] ));
 sg13g2_nor2_1 _2628_ (.A(\bp_core.addr_reg[9] ),
    .B(\bp_core.bp_stride_out[9] ),
    .Y(_0780_));
 sg13g2_xor2_1 _2629_ (.B(\bp_core.bp_stride_out[9] ),
    .A(\bp_core.addr_reg[9] ),
    .X(_0781_));
 sg13g2_nand3_1 _2630_ (.B(_0778_),
    .C(_0781_),
    .A(_0775_),
    .Y(_0782_));
 sg13g2_nor2_1 _2631_ (.A(_0771_),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_a21oi_1 _2632_ (.A1(_0777_),
    .A2(_0779_),
    .Y(_0784_),
    .B1(_0780_));
 sg13g2_a21oi_1 _2633_ (.A1(_0538_),
    .A2(_0539_),
    .Y(_0785_),
    .B1(_0773_));
 sg13g2_a221oi_1 _2634_ (.B2(_0784_),
    .C1(_0785_),
    .B1(_0775_),
    .A1(\bp_core.addr_reg[11] ),
    .Y(_0786_),
    .A2(\bp_core.bp_stride_out[11] ));
 sg13g2_o21ai_1 _2635_ (.B1(_0765_),
    .Y(_0787_),
    .A1(_0766_),
    .A2(_0769_));
 sg13g2_a21oi_1 _2636_ (.A1(_0759_),
    .A2(_0761_),
    .Y(_0788_),
    .B1(_0758_));
 sg13g2_o21ai_1 _2637_ (.B1(_0788_),
    .Y(_0789_),
    .A1(_0771_),
    .A2(_0786_));
 sg13g2_a221oi_1 _2638_ (.B2(_0764_),
    .C1(_0789_),
    .B1(_0787_),
    .A1(_0757_),
    .Y(_0790_),
    .A2(_0783_));
 sg13g2_nand2_1 _2639_ (.Y(_0791_),
    .A(\bp_core.bp_stride_out[16] ),
    .B(\bp_core.addr_reg[16] ));
 sg13g2_xnor2_1 _2640_ (.Y(_0792_),
    .A(\bp_core.bp_stride_out[16] ),
    .B(\bp_core.addr_reg[16] ));
 sg13g2_xor2_1 _2641_ (.B(_0792_),
    .A(_0790_),
    .X(_0793_));
 sg13g2_xor2_1 _2642_ (.B(\bp_core.addr_reg[17] ),
    .A(\bp_core.bp_stride_out[17] ),
    .X(_0794_));
 sg13g2_o21ai_1 _2643_ (.B1(_0791_),
    .Y(_0795_),
    .A1(_0790_),
    .A2(_0792_));
 sg13g2_xor2_1 _2644_ (.B(_0795_),
    .A(_0794_),
    .X(_0796_));
 sg13g2_nand2b_1 _2645_ (.Y(_0797_),
    .B(_0794_),
    .A_N(_0792_));
 sg13g2_a21oi_1 _2646_ (.A1(_0544_),
    .A2(_0545_),
    .Y(_0798_),
    .B1(_0791_));
 sg13g2_a21oi_1 _2647_ (.A1(\bp_core.bp_stride_out[17] ),
    .A2(\bp_core.addr_reg[17] ),
    .Y(_0799_),
    .B1(_0798_));
 sg13g2_o21ai_1 _2648_ (.B1(_0799_),
    .Y(_0800_),
    .A1(_0790_),
    .A2(_0797_));
 sg13g2_and2_1 _2649_ (.A(\bp_core.bp_stride_out[18] ),
    .B(\bp_core.addr_reg[18] ),
    .X(_0801_));
 sg13g2_or2_1 _2650_ (.X(_0802_),
    .B(\bp_core.addr_reg[18] ),
    .A(\bp_core.bp_stride_out[18] ));
 sg13g2_nand2b_1 _2651_ (.Y(_0803_),
    .B(_0802_),
    .A_N(_0801_));
 sg13g2_xnor2_1 _2652_ (.Y(_0804_),
    .A(_0800_),
    .B(_0803_));
 sg13g2_nor3_1 _2653_ (.A(_0793_),
    .B(_0796_),
    .C(_0804_),
    .Y(_0805_));
 sg13g2_a21oi_1 _2654_ (.A1(_0800_),
    .A2(_0802_),
    .Y(_0806_),
    .B1(_0801_));
 sg13g2_xnor2_1 _2655_ (.Y(_0807_),
    .A(\bp_core.bp_stride_out[19] ),
    .B(\bp_core.addr_reg[19] ));
 sg13g2_xnor2_1 _2656_ (.Y(_0808_),
    .A(_0806_),
    .B(_0807_));
 sg13g2_nor2_1 _2657_ (.A(net717),
    .B(_0805_),
    .Y(_0809_));
 sg13g2_a21oi_1 _2658_ (.A1(_0805_),
    .A2(_0808_),
    .Y(_0810_),
    .B1(net717));
 sg13g2_a21oi_1 _2659_ (.A1(net1132),
    .A2(_0728_),
    .Y(_0811_),
    .B1(_0810_));
 sg13g2_a21oi_1 _2660_ (.A1(_0725_),
    .A2(_0811_),
    .Y(_0008_),
    .B1(net749));
 sg13g2_nand3_1 _2661_ (.B(net1110),
    .C(_0685_),
    .A(net756),
    .Y(_0812_));
 sg13g2_nor2_2 _2662_ (.A(net292),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_nor2_1 _2663_ (.A(\bp_core.initialized ),
    .B(net359),
    .Y(_0814_));
 sg13g2_nor2_1 _2664_ (.A(net756),
    .B(_0549_),
    .Y(_0815_));
 sg13g2_o21ai_1 _2665_ (.B1(_0685_),
    .Y(_0816_),
    .A1(_0814_),
    .A2(_0815_));
 sg13g2_o21ai_1 _2666_ (.B1(_0816_),
    .Y(_0010_),
    .A1(net292),
    .A2(_0812_));
 sg13g2_nand3_1 _2667_ (.B(spi_cs),
    .C(net755),
    .A(net1166),
    .Y(_0817_));
 sg13g2_inv_4 _2668_ (.A(net610),
    .Y(_0011_));
 sg13g2_and3_1 _2669_ (.X(_0012_),
    .A(net167),
    .B(\bp_core.state[2] ),
    .C(net755));
 sg13g2_nor3_1 _2670_ (.A(_0686_),
    .B(spi_cs),
    .C(_0708_),
    .Y(_0013_));
 sg13g2_nand2_2 _2671_ (.Y(_0818_),
    .A(net310),
    .B(_0685_));
 sg13g2_nand2_1 _2672_ (.Y(_0819_),
    .A(net215),
    .B(_0688_));
 sg13g2_nand2_1 _2673_ (.Y(_0003_),
    .A(net716),
    .B(_0819_));
 sg13g2_nor3_1 _2674_ (.A(_0687_),
    .B(_0703_),
    .C(net749),
    .Y(_0004_));
 sg13g2_nand2_1 _2675_ (.Y(_0820_),
    .A(net1132),
    .B(_0727_));
 sg13g2_and2_1 _2676_ (.A(net721),
    .B(_0808_),
    .X(_0821_));
 sg13g2_nand3_1 _2677_ (.B(_0805_),
    .C(_0808_),
    .A(net721),
    .Y(_0822_));
 sg13g2_nand2_1 _2678_ (.Y(_0823_),
    .A(net929),
    .B(_0687_));
 sg13g2_nand3_1 _2679_ (.B(_0822_),
    .C(_0823_),
    .A(_0820_),
    .Y(_0824_));
 sg13g2_and2_1 _2680_ (.A(net755),
    .B(_0824_),
    .X(_0009_));
 sg13g2_a21o_2 _2681_ (.A2(_0699_),
    .A1(net368),
    .B1(_0689_),
    .X(_0825_));
 sg13g2_nor2_2 _2682_ (.A(_0550_),
    .B(_0812_),
    .Y(_0826_));
 sg13g2_o21ai_1 _2683_ (.B1(_0825_),
    .Y(_0007_),
    .A1(_0550_),
    .A2(_0812_));
 sg13g2_o21ai_1 _2684_ (.B1(_0713_),
    .Y(_0827_),
    .A1(net756),
    .A2(\bp_core.bp_param_valid_in ));
 sg13g2_nand2b_1 _2685_ (.Y(_0828_),
    .B(net963),
    .A_N(net167));
 sg13g2_o21ai_1 _2686_ (.B1(_0827_),
    .Y(_0006_),
    .A1(net749),
    .A2(_0828_));
 sg13g2_nand3_1 _2687_ (.B(net733),
    .C(_0720_),
    .A(net756),
    .Y(_0829_));
 sg13g2_nand2b_1 _2688_ (.Y(_0830_),
    .B(\bp_core.bp_param_ack_out ),
    .A_N(net922));
 sg13g2_o21ai_1 _2689_ (.B1(_0829_),
    .Y(_1800_[0]),
    .A1(net77),
    .A2(net923));
 sg13g2_nand2b_1 _2690_ (.Y(_0831_),
    .B(net198),
    .A_N(net1026));
 sg13g2_nand2b_1 _2691_ (.Y(_0000_),
    .B(_0831_),
    .A_N(_1800_[0]));
 sg13g2_nor2_1 _2692_ (.A(\bp_core.state[1] ),
    .B(net505),
    .Y(_0832_));
 sg13g2_nor3_1 _2693_ (.A(spi_cs),
    .B(net749),
    .C(net506),
    .Y(_0005_));
 sg13g2_a22oi_1 _2694_ (.Y(_0833_),
    .B1(_0719_),
    .B2(net59),
    .A2(net1026),
    .A1(net198));
 sg13g2_inv_1 _2695_ (.Y(_0002_),
    .A(net1099));
 sg13g2_nand2_1 _2696_ (.Y(_0834_),
    .A(_0525_),
    .B(net731));
 sg13g2_nand2_1 _2697_ (.Y(_0835_),
    .A(net922),
    .B(\bp_core.params_module.state[0] ));
 sg13g2_and2_1 _2698_ (.A(_0834_),
    .B(_0835_),
    .X(_0836_));
 sg13g2_nand2_1 _2699_ (.Y(_0837_),
    .A(net733),
    .B(net1098));
 sg13g2_nand2_1 _2700_ (.Y(_0001_),
    .A(_0836_),
    .B(_0837_));
 sg13g2_nand2_1 _2701_ (.Y(_0838_),
    .A(\bp_core.bp_param_output_data[0] ),
    .B(\bp_core.bp_param_output_valid ));
 sg13g2_o21ai_1 _2702_ (.B1(_0838_),
    .Y(uo_out[3]),
    .A1(_0560_),
    .A2(\bp_core.bp_param_output_valid ));
 sg13g2_mux2_1 _2703_ (.A0(\bp_core.status_out[1] ),
    .A1(\bp_core.bp_param_output_data[1] ),
    .S(\bp_core.bp_param_output_valid ),
    .X(uo_out[4]));
 sg13g2_nand2_1 _2704_ (.Y(_0839_),
    .A(\bp_core.bp_param_output_valid ),
    .B(\bp_core.bp_param_output_data[2] ));
 sg13g2_o21ai_1 _2705_ (.B1(_0839_),
    .Y(uo_out[5]),
    .A1(\bp_core.bp_param_output_valid ),
    .A2(_0561_));
 sg13g2_mux2_1 _2706_ (.A0(\bp_core.status_out[3] ),
    .A1(\bp_core.bp_param_output_data[3] ),
    .S(\bp_core.bp_param_output_valid ),
    .X(uo_out[6]));
 sg13g2_mux2_1 _2707_ (.A0(\bp_core.status_out[4] ),
    .A1(\bp_core.bp_param_output_data[4] ),
    .S(\bp_core.bp_param_output_valid ),
    .X(uo_out[7]));
 sg13g2_and2_1 _2708_ (.A(\bp_core.bp_param_ack_out ),
    .B(\inter_bp.param_pending ),
    .X(_0840_));
 sg13g2_nand2_1 _2709_ (.Y(_0841_),
    .A(\bp_core.bp_param_ack_out ),
    .B(\inter_bp.param_pending ));
 sg13g2_nor2b_2 _2710_ (.A(\bp_core.bp_param_valid_in ),
    .B_N(\inter_bp.param_rx_done ),
    .Y(_0842_));
 sg13g2_nand2b_2 _2711_ (.Y(_0843_),
    .B(net890),
    .A_N(\bp_core.bp_param_valid_in ));
 sg13g2_nand2b_1 _2712_ (.Y(_0844_),
    .B(net1140),
    .A_N(net1125));
 sg13g2_nand3_1 _2713_ (.B(net685),
    .C(_0844_),
    .A(net704),
    .Y(_0072_));
 sg13g2_nand2_1 _2714_ (.Y(_0845_),
    .A(net397),
    .B(net695));
 sg13g2_nor2_1 _2715_ (.A(\inter_bp.param_pending_reg[0] ),
    .B(net708),
    .Y(_0846_));
 sg13g2_o21ai_1 _2716_ (.B1(net688),
    .Y(_0847_),
    .A1(\bp_addr_in[0] ),
    .A2(_0840_));
 sg13g2_o21ai_1 _2717_ (.B1(_0845_),
    .Y(_0044_),
    .A1(_0846_),
    .A2(_0847_));
 sg13g2_a21oi_1 _2718_ (.A1(_0562_),
    .A2(net714),
    .Y(_0848_),
    .B1(net697));
 sg13g2_o21ai_1 _2719_ (.B1(_0848_),
    .Y(_0849_),
    .A1(net562),
    .A2(net714));
 sg13g2_o21ai_1 _2720_ (.B1(_0849_),
    .Y(_0055_),
    .A1(_0563_),
    .A2(net690));
 sg13g2_a21oi_1 _2721_ (.A1(_0564_),
    .A2(net710),
    .Y(_0850_),
    .B1(net698));
 sg13g2_o21ai_1 _2722_ (.B1(_0850_),
    .Y(_0851_),
    .A1(net490),
    .A2(net709));
 sg13g2_o21ai_1 _2723_ (.B1(_0851_),
    .Y(_0056_),
    .A1(_0565_),
    .A2(net691));
 sg13g2_a21oi_1 _2724_ (.A1(_0566_),
    .A2(net714),
    .Y(_0852_),
    .B1(net696));
 sg13g2_o21ai_1 _2725_ (.B1(_0852_),
    .Y(_0853_),
    .A1(net894),
    .A2(net711));
 sg13g2_o21ai_1 _2726_ (.B1(_0853_),
    .Y(_0057_),
    .A1(_0567_),
    .A2(net690));
 sg13g2_a21oi_1 _2727_ (.A1(_0568_),
    .A2(net713),
    .Y(_0854_),
    .B1(net696));
 sg13g2_o21ai_1 _2728_ (.B1(_0854_),
    .Y(_0855_),
    .A1(net510),
    .A2(net713));
 sg13g2_o21ai_1 _2729_ (.B1(_0855_),
    .Y(_0058_),
    .A1(_0569_),
    .A2(net689));
 sg13g2_a21oi_1 _2730_ (.A1(_0570_),
    .A2(net712),
    .Y(_0856_),
    .B1(net696));
 sg13g2_o21ai_1 _2731_ (.B1(_0856_),
    .Y(_0857_),
    .A1(net553),
    .A2(net712));
 sg13g2_o21ai_1 _2732_ (.B1(_0857_),
    .Y(_0059_),
    .A1(_0571_),
    .A2(net689));
 sg13g2_a21oi_1 _2733_ (.A1(_0572_),
    .A2(net712),
    .Y(_0858_),
    .B1(net696));
 sg13g2_o21ai_1 _2734_ (.B1(_0858_),
    .Y(_0859_),
    .A1(net514),
    .A2(net713));
 sg13g2_o21ai_1 _2735_ (.B1(_0859_),
    .Y(_0060_),
    .A1(_0573_),
    .A2(net689));
 sg13g2_a21oi_1 _2736_ (.A1(_0574_),
    .A2(net711),
    .Y(_0860_),
    .B1(net696));
 sg13g2_o21ai_1 _2737_ (.B1(_0860_),
    .Y(_0861_),
    .A1(net851),
    .A2(net711));
 sg13g2_o21ai_1 _2738_ (.B1(_0861_),
    .Y(_0061_),
    .A1(_0575_),
    .A2(net689));
 sg13g2_a21oi_1 _2739_ (.A1(_0576_),
    .A2(net712),
    .Y(_0862_),
    .B1(net696));
 sg13g2_o21ai_1 _2740_ (.B1(_0862_),
    .Y(_0863_),
    .A1(net531),
    .A2(net712));
 sg13g2_o21ai_1 _2741_ (.B1(_0863_),
    .Y(_0062_),
    .A1(_0577_),
    .A2(net689));
 sg13g2_a21oi_1 _2742_ (.A1(_0578_),
    .A2(net711),
    .Y(_0864_),
    .B1(net696));
 sg13g2_o21ai_1 _2743_ (.B1(_0864_),
    .Y(_0865_),
    .A1(net860),
    .A2(net711));
 sg13g2_o21ai_1 _2744_ (.B1(_0865_),
    .Y(_0063_),
    .A1(_0579_),
    .A2(net690));
 sg13g2_a21oi_1 _2745_ (.A1(_0580_),
    .A2(net711),
    .Y(_0866_),
    .B1(net697));
 sg13g2_o21ai_1 _2746_ (.B1(_0866_),
    .Y(_0867_),
    .A1(net842),
    .A2(net711));
 sg13g2_o21ai_1 _2747_ (.B1(_0867_),
    .Y(_0045_),
    .A1(_0581_),
    .A2(net689));
 sg13g2_a21oi_1 _2748_ (.A1(_0582_),
    .A2(net711),
    .Y(_0868_),
    .B1(net697));
 sg13g2_o21ai_1 _2749_ (.B1(_0868_),
    .Y(_0869_),
    .A1(net523),
    .A2(net713));
 sg13g2_o21ai_1 _2750_ (.B1(_0869_),
    .Y(_0046_),
    .A1(_0583_),
    .A2(net689));
 sg13g2_a21oi_1 _2751_ (.A1(_0584_),
    .A2(net713),
    .Y(_0870_),
    .B1(net696));
 sg13g2_o21ai_1 _2752_ (.B1(_0870_),
    .Y(_0871_),
    .A1(net470),
    .A2(net713));
 sg13g2_o21ai_1 _2753_ (.B1(_0871_),
    .Y(_0047_),
    .A1(_0585_),
    .A2(net689));
 sg13g2_a21oi_1 _2754_ (.A1(_0586_),
    .A2(net709),
    .Y(_0872_),
    .B1(net698));
 sg13g2_o21ai_1 _2755_ (.B1(_0872_),
    .Y(_0873_),
    .A1(net565),
    .A2(net710));
 sg13g2_o21ai_1 _2756_ (.B1(_0873_),
    .Y(_0048_),
    .A1(_0587_),
    .A2(net691));
 sg13g2_a21oi_1 _2757_ (.A1(_0588_),
    .A2(net710),
    .Y(_0874_),
    .B1(net698));
 sg13g2_o21ai_1 _2758_ (.B1(_0874_),
    .Y(_0875_),
    .A1(net900),
    .A2(net710));
 sg13g2_o21ai_1 _2759_ (.B1(_0875_),
    .Y(_0049_),
    .A1(_0589_),
    .A2(net691));
 sg13g2_a21oi_1 _2760_ (.A1(_0590_),
    .A2(net707),
    .Y(_0876_),
    .B1(net695));
 sg13g2_o21ai_1 _2761_ (.B1(_0876_),
    .Y(_0877_),
    .A1(net875),
    .A2(net707));
 sg13g2_o21ai_1 _2762_ (.B1(_0877_),
    .Y(_0050_),
    .A1(_0591_),
    .A2(net688));
 sg13g2_a21oi_1 _2763_ (.A1(_0592_),
    .A2(net706),
    .Y(_0878_),
    .B1(net695));
 sg13g2_o21ai_1 _2764_ (.B1(_0878_),
    .Y(_0879_),
    .A1(net845),
    .A2(net706));
 sg13g2_o21ai_1 _2765_ (.B1(_0879_),
    .Y(_0051_),
    .A1(_0593_),
    .A2(net688));
 sg13g2_a21oi_1 _2766_ (.A1(_0594_),
    .A2(net700),
    .Y(_0880_),
    .B1(net694));
 sg13g2_o21ai_1 _2767_ (.B1(_0880_),
    .Y(_0881_),
    .A1(net476),
    .A2(net700));
 sg13g2_o21ai_1 _2768_ (.B1(_0881_),
    .Y(_0052_),
    .A1(_0595_),
    .A2(net684));
 sg13g2_a21oi_1 _2769_ (.A1(_0596_),
    .A2(net706),
    .Y(_0882_),
    .B1(net695));
 sg13g2_o21ai_1 _2770_ (.B1(_0882_),
    .Y(_0883_),
    .A1(net896),
    .A2(net706));
 sg13g2_o21ai_1 _2771_ (.B1(net897),
    .Y(_0053_),
    .A1(_0597_),
    .A2(net688));
 sg13g2_a21oi_1 _2772_ (.A1(_0598_),
    .A2(net700),
    .Y(_0884_),
    .B1(net694));
 sg13g2_o21ai_1 _2773_ (.B1(_0884_),
    .Y(_0885_),
    .A1(net560),
    .A2(net700));
 sg13g2_o21ai_1 _2774_ (.B1(_0885_),
    .Y(_0054_),
    .A1(_0599_),
    .A2(net687));
 sg13g2_a21oi_1 _2775_ (.A1(_0600_),
    .A2(net707),
    .Y(_0886_),
    .B1(_0842_));
 sg13g2_o21ai_1 _2776_ (.B1(_0886_),
    .Y(_0887_),
    .A1(net478),
    .A2(net707));
 sg13g2_o21ai_1 _2777_ (.B1(_0887_),
    .Y(_0073_),
    .A1(_0601_),
    .A2(_0843_));
 sg13g2_a21oi_1 _2778_ (.A1(_0602_),
    .A2(net700),
    .Y(_0888_),
    .B1(net692));
 sg13g2_o21ai_1 _2779_ (.B1(_0888_),
    .Y(_0889_),
    .A1(net488),
    .A2(net700));
 sg13g2_o21ai_1 _2780_ (.B1(_0889_),
    .Y(_0084_),
    .A1(_0603_),
    .A2(net687));
 sg13g2_a21oi_1 _2781_ (.A1(_0604_),
    .A2(net709),
    .Y(_0890_),
    .B1(net698));
 sg13g2_o21ai_1 _2782_ (.B1(_0890_),
    .Y(_0891_),
    .A1(net509),
    .A2(net709));
 sg13g2_o21ai_1 _2783_ (.B1(_0891_),
    .Y(_0085_),
    .A1(_0605_),
    .A2(net691));
 sg13g2_a21oi_1 _2784_ (.A1(_0606_),
    .A2(net700),
    .Y(_0892_),
    .B1(net692));
 sg13g2_o21ai_1 _2785_ (.B1(_0892_),
    .Y(_0893_),
    .A1(net474),
    .A2(net699));
 sg13g2_o21ai_1 _2786_ (.B1(_0893_),
    .Y(_0086_),
    .A1(_0607_),
    .A2(net684));
 sg13g2_a21oi_1 _2787_ (.A1(_0608_),
    .A2(net710),
    .Y(_0894_),
    .B1(net698));
 sg13g2_o21ai_1 _2788_ (.B1(_0894_),
    .Y(_0895_),
    .A1(net551),
    .A2(net709));
 sg13g2_o21ai_1 _2789_ (.B1(_0895_),
    .Y(_0087_),
    .A1(_0609_),
    .A2(net691));
 sg13g2_a21oi_1 _2790_ (.A1(_0610_),
    .A2(net699),
    .Y(_0896_),
    .B1(net692));
 sg13g2_o21ai_1 _2791_ (.B1(_0896_),
    .Y(_0897_),
    .A1(net473),
    .A2(net699));
 sg13g2_o21ai_1 _2792_ (.B1(_0897_),
    .Y(_0088_),
    .A1(_0611_),
    .A2(net684));
 sg13g2_a21oi_1 _2793_ (.A1(_0612_),
    .A2(net710),
    .Y(_0898_),
    .B1(net698));
 sg13g2_o21ai_1 _2794_ (.B1(_0898_),
    .Y(_0899_),
    .A1(net870),
    .A2(net709));
 sg13g2_o21ai_1 _2795_ (.B1(net871),
    .Y(_0089_),
    .A1(_0613_),
    .A2(net691));
 sg13g2_a21oi_1 _2796_ (.A1(_0614_),
    .A2(net699),
    .Y(_0900_),
    .B1(net692));
 sg13g2_o21ai_1 _2797_ (.B1(_0900_),
    .Y(_0901_),
    .A1(net472),
    .A2(net699));
 sg13g2_o21ai_1 _2798_ (.B1(_0901_),
    .Y(_0090_),
    .A1(_0615_),
    .A2(net684));
 sg13g2_a21oi_1 _2799_ (.A1(_0616_),
    .A2(net709),
    .Y(_0902_),
    .B1(net698));
 sg13g2_o21ai_1 _2800_ (.B1(_0902_),
    .Y(_0903_),
    .A1(net518),
    .A2(net709));
 sg13g2_o21ai_1 _2801_ (.B1(_0903_),
    .Y(_0091_),
    .A1(_0617_),
    .A2(net691));
 sg13g2_a21oi_1 _2802_ (.A1(_0618_),
    .A2(net699),
    .Y(_0904_),
    .B1(net692));
 sg13g2_o21ai_1 _2803_ (.B1(_0904_),
    .Y(_0905_),
    .A1(net527),
    .A2(net701));
 sg13g2_o21ai_1 _2804_ (.B1(_0905_),
    .Y(_0092_),
    .A1(_0619_),
    .A2(net684));
 sg13g2_a21oi_1 _2805_ (.A1(_0620_),
    .A2(net707),
    .Y(_0906_),
    .B1(net695));
 sg13g2_o21ai_1 _2806_ (.B1(_0906_),
    .Y(_0907_),
    .A1(net859),
    .A2(net707));
 sg13g2_o21ai_1 _2807_ (.B1(_0907_),
    .Y(_0074_),
    .A1(_0621_),
    .A2(net688));
 sg13g2_nand2_1 _2808_ (.Y(_0908_),
    .A(net427),
    .B(net692));
 sg13g2_nor2_1 _2809_ (.A(\inter_bp.param_pending_reg[31] ),
    .B(net699),
    .Y(_0909_));
 sg13g2_o21ai_1 _2810_ (.B1(net685),
    .Y(_0910_),
    .A1(\bp_core.bp_stride_in[11] ),
    .A2(_0840_));
 sg13g2_o21ai_1 _2811_ (.B1(_0908_),
    .Y(_0075_),
    .A1(_0909_),
    .A2(_0910_));
 sg13g2_a21oi_1 _2812_ (.A1(_0622_),
    .A2(net706),
    .Y(_0911_),
    .B1(net695));
 sg13g2_o21ai_1 _2813_ (.B1(_0911_),
    .Y(_0912_),
    .A1(net464),
    .A2(net707));
 sg13g2_o21ai_1 _2814_ (.B1(_0912_),
    .Y(_0076_),
    .A1(_0623_),
    .A2(net688));
 sg13g2_a21oi_1 _2815_ (.A1(_0624_),
    .A2(net699),
    .Y(_0913_),
    .B1(net692));
 sg13g2_o21ai_1 _2816_ (.B1(_0913_),
    .Y(_0914_),
    .A1(net468),
    .A2(net701));
 sg13g2_o21ai_1 _2817_ (.B1(_0914_),
    .Y(_0077_),
    .A1(_0625_),
    .A2(net684));
 sg13g2_a21oi_1 _2818_ (.A1(_0626_),
    .A2(net706),
    .Y(_0915_),
    .B1(net695));
 sg13g2_o21ai_1 _2819_ (.B1(_0915_),
    .Y(_0916_),
    .A1(net500),
    .A2(net706));
 sg13g2_o21ai_1 _2820_ (.B1(_0916_),
    .Y(_0078_),
    .A1(_0627_),
    .A2(net688));
 sg13g2_a21oi_1 _2821_ (.A1(_0628_),
    .A2(net702),
    .Y(_0917_),
    .B1(net692));
 sg13g2_o21ai_1 _2822_ (.B1(_0917_),
    .Y(_0918_),
    .A1(net507),
    .A2(net701));
 sg13g2_o21ai_1 _2823_ (.B1(_0918_),
    .Y(_0079_),
    .A1(_0629_),
    .A2(net684));
 sg13g2_a21oi_1 _2824_ (.A1(_0630_),
    .A2(net706),
    .Y(_0919_),
    .B1(net694));
 sg13g2_o21ai_1 _2825_ (.B1(_0919_),
    .Y(_0920_),
    .A1(net466),
    .A2(net700));
 sg13g2_o21ai_1 _2826_ (.B1(_0920_),
    .Y(_0080_),
    .A1(_0631_),
    .A2(net684));
 sg13g2_a21oi_1 _2827_ (.A1(_0632_),
    .A2(net702),
    .Y(_0921_),
    .B1(net693));
 sg13g2_o21ai_1 _2828_ (.B1(_0921_),
    .Y(_0922_),
    .A1(net546),
    .A2(net702));
 sg13g2_o21ai_1 _2829_ (.B1(_0922_),
    .Y(_0081_),
    .A1(_0633_),
    .A2(net685));
 sg13g2_a21oi_1 _2830_ (.A1(_0634_),
    .A2(net705),
    .Y(_0923_),
    .B1(net694));
 sg13g2_o21ai_1 _2831_ (.B1(_0923_),
    .Y(_0924_),
    .A1(net545),
    .A2(net701));
 sg13g2_o21ai_1 _2832_ (.B1(_0924_),
    .Y(_0082_),
    .A1(_0635_),
    .A2(net686));
 sg13g2_a21oi_1 _2833_ (.A1(_0636_),
    .A2(net702),
    .Y(_0925_),
    .B1(net693));
 sg13g2_o21ai_1 _2834_ (.B1(_0925_),
    .Y(_0926_),
    .A1(net543),
    .A2(net702));
 sg13g2_o21ai_1 _2835_ (.B1(_0926_),
    .Y(_0083_),
    .A1(_0637_),
    .A2(net685));
 sg13g2_a21oi_1 _2836_ (.A1(_0638_),
    .A2(net704),
    .Y(_0927_),
    .B1(net694));
 sg13g2_o21ai_1 _2837_ (.B1(_0927_),
    .Y(_0928_),
    .A1(net883),
    .A2(net704));
 sg13g2_o21ai_1 _2838_ (.B1(_0928_),
    .Y(_0064_),
    .A1(_0639_),
    .A2(net686));
 sg13g2_nand2_1 _2839_ (.Y(_0929_),
    .A(net349),
    .B(net693));
 sg13g2_nor2_1 _2840_ (.A(\inter_bp.param_pending_reg[41] ),
    .B(net702),
    .Y(_0930_));
 sg13g2_o21ai_1 _2841_ (.B1(net686),
    .Y(_0931_),
    .A1(\bp_core.bp_lambda_in[1] ),
    .A2(_0840_));
 sg13g2_o21ai_1 _2842_ (.B1(_0929_),
    .Y(_0065_),
    .A1(_0930_),
    .A2(_0931_));
 sg13g2_a21oi_1 _2843_ (.A1(_0640_),
    .A2(net704),
    .Y(_0932_),
    .B1(net694));
 sg13g2_o21ai_1 _2844_ (.B1(_0932_),
    .Y(_0933_),
    .A1(net873),
    .A2(net704));
 sg13g2_o21ai_1 _2845_ (.B1(_0933_),
    .Y(_0066_),
    .A1(_0641_),
    .A2(net686));
 sg13g2_a21oi_1 _2846_ (.A1(_0642_),
    .A2(net702),
    .Y(_0934_),
    .B1(net693));
 sg13g2_o21ai_1 _2847_ (.B1(_0934_),
    .Y(_0935_),
    .A1(net537),
    .A2(net703));
 sg13g2_o21ai_1 _2848_ (.B1(_0935_),
    .Y(_0067_),
    .A1(_0643_),
    .A2(net685));
 sg13g2_a21oi_1 _2849_ (.A1(_0644_),
    .A2(net704),
    .Y(_0936_),
    .B1(net693));
 sg13g2_o21ai_1 _2850_ (.B1(_0936_),
    .Y(_0937_),
    .A1(net496),
    .A2(net705));
 sg13g2_o21ai_1 _2851_ (.B1(_0937_),
    .Y(_0068_),
    .A1(_0645_),
    .A2(net686));
 sg13g2_a21oi_1 _2852_ (.A1(_0646_),
    .A2(net703),
    .Y(_0938_),
    .B1(net693));
 sg13g2_o21ai_1 _2853_ (.B1(_0938_),
    .Y(_0939_),
    .A1(net558),
    .A2(net703));
 sg13g2_o21ai_1 _2854_ (.B1(_0939_),
    .Y(_0069_),
    .A1(_0647_),
    .A2(net685));
 sg13g2_a21oi_1 _2855_ (.A1(_0648_),
    .A2(net702),
    .Y(_0940_),
    .B1(net693));
 sg13g2_o21ai_1 _2856_ (.B1(_0940_),
    .Y(_0941_),
    .A1(net502),
    .A2(net703));
 sg13g2_o21ai_1 _2857_ (.B1(_0941_),
    .Y(_0070_),
    .A1(_0649_),
    .A2(net685));
 sg13g2_a21oi_1 _2858_ (.A1(_0650_),
    .A2(net703),
    .Y(_0942_),
    .B1(net693));
 sg13g2_o21ai_1 _2859_ (.B1(_0942_),
    .Y(_0943_),
    .A1(net541),
    .A2(net703));
 sg13g2_o21ai_1 _2860_ (.B1(_0943_),
    .Y(_0071_),
    .A1(_0651_),
    .A2(net685));
 sg13g2_nand2_2 _2861_ (.Y(_0944_),
    .A(\inter_bp.param_rx_done ),
    .B(\bp_core.bp_param_valid_in ));
 sg13g2_o21ai_1 _2862_ (.B1(net677),
    .Y(_0093_),
    .A1(\bp_core.bp_param_ack_out ),
    .A2(_0553_));
 sg13g2_nor3_1 _2863_ (.A(\inter_bp.from_left_param_valid_prev ),
    .B(_0552_),
    .C(net968),
    .Y(_0945_));
 sg13g2_nor2_1 _2864_ (.A(net890),
    .B(_0945_),
    .Y(_0946_));
 sg13g2_nor4_2 _2865_ (.A(_0552_),
    .B(\inter_bp.param_rx_done ),
    .C(_0558_),
    .Y(_0947_),
    .D(_0945_));
 sg13g2_nand3_1 _2866_ (.B(\inter_bp.param_receiving ),
    .C(_0946_),
    .A(net10),
    .Y(_0948_));
 sg13g2_and3_2 _2867_ (.X(_0949_),
    .A(net1181),
    .B(net288),
    .C(net395));
 sg13g2_nand3b_1 _2868_ (.B(net229),
    .C(_0949_),
    .Y(_0950_),
    .A_N(\inter_bp.param_rx_counter[3] ));
 sg13g2_nor2_1 _2869_ (.A(_0948_),
    .B(net230),
    .Y(_0094_));
 sg13g2_nand2_1 _2870_ (.Y(_0951_),
    .A(net855),
    .B(net11));
 sg13g2_nor2_1 _2871_ (.A(net746),
    .B(_0951_),
    .Y(_0952_));
 sg13g2_and2_1 _2872_ (.A(net461),
    .B(_0952_),
    .X(_0953_));
 sg13g2_and2_1 _2873_ (.A(net308),
    .B(net448),
    .X(_0954_));
 sg13g2_nor3_1 _2874_ (.A(net322),
    .B(\inter_bp.report_rx_counter[1] ),
    .C(net1063),
    .Y(_0955_));
 sg13g2_and3_1 _2875_ (.X(_0096_),
    .A(net608),
    .B(_0954_),
    .C(net1064));
 sg13g2_nor2b_1 _2876_ (.A(\inter_bp.param_transmitting ),
    .B_N(\inter_bp.report_transmitting ),
    .Y(_0956_));
 sg13g2_a22oi_1 _2877_ (.Y(_0957_),
    .B1(_0956_),
    .B2(\inter_bp.report_tx_shift_reg[0] ),
    .A2(\inter_bp.param_tx_shift_reg[0] ),
    .A1(\inter_bp.param_transmitting ));
 sg13g2_inv_1 _2878_ (.Y(uio_out[6]),
    .A(_0957_));
 sg13g2_a22oi_1 _2879_ (.Y(_0958_),
    .B1(_0956_),
    .B2(\inter_bp.report_tx_shift_reg[1] ),
    .A2(\inter_bp.param_tx_shift_reg[1] ),
    .A1(\inter_bp.param_transmitting ));
 sg13g2_inv_1 _2880_ (.Y(uio_out[7]),
    .A(_0958_));
 sg13g2_a22oi_1 _2881_ (.Y(_0959_),
    .B1(\bp_core.threshold_reg[5] ),
    .B2(_0658_),
    .A2(_0657_),
    .A1(_0523_));
 sg13g2_nand2b_1 _2882_ (.Y(_0960_),
    .B(\bp_core.data_reg[5] ),
    .A_N(\bp_core.threshold_reg[5] ));
 sg13g2_nor2_1 _2883_ (.A(_0659_),
    .B(\bp_core.threshold_reg[4] ),
    .Y(_0961_));
 sg13g2_nand2_1 _2884_ (.Y(_0962_),
    .A(_0659_),
    .B(\bp_core.threshold_reg[4] ));
 sg13g2_o21ai_1 _2885_ (.B1(_0962_),
    .Y(_0963_),
    .A1(_0101_),
    .A2(\bp_core.data_reg[3] ));
 sg13g2_a22oi_1 _2886_ (.Y(_0964_),
    .B1(\bp_core.data_reg[0] ),
    .B2(_0666_),
    .A2(\bp_core.data_reg[1] ),
    .A1(_0663_));
 sg13g2_a221oi_1 _2887_ (.B2(_0664_),
    .C1(_0964_),
    .B1(\bp_core.threshold_reg[1] ),
    .A1(\bp_core.threshold_reg[2] ),
    .Y(_0965_),
    .A2(_0662_));
 sg13g2_a221oi_1 _2888_ (.B2(\bp_core.data_reg[2] ),
    .C1(_0965_),
    .B1(_0661_),
    .A1(_0101_),
    .Y(_0966_),
    .A2(\bp_core.data_reg[3] ));
 sg13g2_o21ai_1 _2889_ (.B1(_0960_),
    .Y(_0967_),
    .A1(_0963_),
    .A2(_0966_));
 sg13g2_o21ai_1 _2890_ (.B1(_0959_),
    .Y(_0968_),
    .A1(_0961_),
    .A2(_0967_));
 sg13g2_a22oi_1 _2891_ (.Y(_0969_),
    .B1(\bp_core.data_reg[6] ),
    .B2(_0099_),
    .A2(\bp_core.data_reg[7] ),
    .A1(_0100_));
 sg13g2_nand2_1 _2892_ (.Y(_0970_),
    .A(net722),
    .B(net755));
 sg13g2_a221oi_1 _2893_ (.B2(_0969_),
    .C1(_0970_),
    .B1(_0968_),
    .A1(_0522_),
    .Y(_0971_),
    .A2(_0656_));
 sg13g2_nand3_1 _2894_ (.B(net2),
    .C(net1),
    .A(net3),
    .Y(_0972_));
 sg13g2_nor2b_2 _2895_ (.A(net741),
    .B_N(_0972_),
    .Y(_0973_));
 sg13g2_nor2b_1 _2896_ (.A(net574),
    .B_N(_0973_),
    .Y(_0974_));
 sg13g2_inv_2 _2897_ (.Y(_0034_),
    .A(net570));
 sg13g2_nor2b_1 _2898_ (.A(net741),
    .B_N(net4),
    .Y(_0975_));
 sg13g2_a21oi_1 _2899_ (.A1(net741),
    .A2(\inter_bp.bp_report_addr_out[0] ),
    .Y(_0976_),
    .B1(_0975_));
 sg13g2_nor3_1 _2900_ (.A(net576),
    .B(_0973_),
    .C(_0976_),
    .Y(_0977_));
 sg13g2_a21oi_1 _2901_ (.A1(\bp_core.addr_reg[0] ),
    .A2(net577),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_o21ai_1 _2902_ (.B1(_0978_),
    .Y(_0014_),
    .A1(_0653_),
    .A2(_0034_));
 sg13g2_nand2b_1 _2903_ (.Y(_0979_),
    .B(net742),
    .A_N(\inter_bp.bp_report_addr_out[1] ));
 sg13g2_o21ai_1 _2904_ (.B1(_0979_),
    .Y(_0980_),
    .A1(net5),
    .A2(net741));
 sg13g2_nor3_1 _2905_ (.A(net576),
    .B(_0973_),
    .C(_0980_),
    .Y(_0981_));
 sg13g2_a21o_1 _2906_ (.A2(net576),
    .A1(net446),
    .B1(_0981_),
    .X(_0982_));
 sg13g2_a21o_1 _2907_ (.A2(net570),
    .A1(net247),
    .B1(_0982_),
    .X(_0025_));
 sg13g2_nor2b_1 _2908_ (.A(net741),
    .B_N(net6),
    .Y(_0983_));
 sg13g2_a21oi_1 _2909_ (.A1(net741),
    .A2(\inter_bp.bp_report_addr_out[2] ),
    .Y(_0984_),
    .B1(_0983_));
 sg13g2_nor3_1 _2910_ (.A(net577),
    .B(_0973_),
    .C(_0984_),
    .Y(_0985_));
 sg13g2_a21oi_1 _2911_ (.A1(net333),
    .A2(net576),
    .Y(_0986_),
    .B1(_0985_));
 sg13g2_o21ai_1 _2912_ (.B1(net334),
    .Y(_0026_),
    .A1(_0654_),
    .A2(_0034_));
 sg13g2_nand2b_1 _2913_ (.Y(_0987_),
    .B(net742),
    .A_N(\inter_bp.bp_report_addr_out[3] ));
 sg13g2_o21ai_1 _2914_ (.B1(_0987_),
    .Y(_0988_),
    .A1(net7),
    .A2(net741));
 sg13g2_nor2_1 _2915_ (.A(_0973_),
    .B(_0988_),
    .Y(_0989_));
 sg13g2_nor2_1 _2916_ (.A(net576),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_a21oi_1 _2917_ (.A1(_0530_),
    .A2(net576),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_a21o_1 _2918_ (.A2(net570),
    .A1(net847),
    .B1(_0991_),
    .X(_0027_));
 sg13g2_nor2b_1 _2919_ (.A(net741),
    .B_N(net8),
    .Y(_0992_));
 sg13g2_a21oi_1 _2920_ (.A1(net743),
    .A2(\inter_bp.bp_report_addr_out[4] ),
    .Y(_0993_),
    .B1(_0992_));
 sg13g2_nor3_1 _2921_ (.A(net576),
    .B(_0973_),
    .C(_0993_),
    .Y(_0994_));
 sg13g2_a21o_1 _2922_ (.A2(net576),
    .A1(net371),
    .B1(_0994_),
    .X(_0995_));
 sg13g2_a21o_1 _2923_ (.A2(net571),
    .A1(net115),
    .B1(net372),
    .X(_0028_));
 sg13g2_nand2_1 _2924_ (.Y(_0996_),
    .A(net742),
    .B(net281));
 sg13g2_a22oi_1 _2925_ (.Y(_0997_),
    .B1(net570),
    .B2(\bp_core.bp_report_addr_out[5] ),
    .A2(net575),
    .A1(\bp_core.addr_reg[5] ));
 sg13g2_o21ai_1 _2926_ (.B1(_0997_),
    .Y(_0029_),
    .A1(net575),
    .A2(net282));
 sg13g2_nand2_1 _2927_ (.Y(_0998_),
    .A(net742),
    .B(net328));
 sg13g2_a22oi_1 _2928_ (.Y(_0999_),
    .B1(net571),
    .B2(net208),
    .A2(net575),
    .A1(\bp_core.addr_reg[6] ));
 sg13g2_o21ai_1 _2929_ (.B1(_0999_),
    .Y(_0030_),
    .A1(net578),
    .A2(net329));
 sg13g2_nand2_1 _2930_ (.Y(_1000_),
    .A(net742),
    .B(net261));
 sg13g2_a22oi_1 _2931_ (.Y(_1001_),
    .B1(net569),
    .B2(net124),
    .A2(net575),
    .A1(\bp_core.addr_reg[7] ));
 sg13g2_o21ai_1 _2932_ (.B1(_1001_),
    .Y(_0031_),
    .A1(net575),
    .A2(net262));
 sg13g2_nand2_1 _2933_ (.Y(_1002_),
    .A(net742),
    .B(net298));
 sg13g2_a22oi_1 _2934_ (.Y(_1003_),
    .B1(net570),
    .B2(net74),
    .A2(net575),
    .A1(\bp_core.addr_reg[8] ));
 sg13g2_o21ai_1 _2935_ (.B1(_1003_),
    .Y(_0032_),
    .A1(net575),
    .A2(net299));
 sg13g2_nand2_1 _2936_ (.Y(_1004_),
    .A(net740),
    .B(net278));
 sg13g2_a22oi_1 _2937_ (.Y(_1005_),
    .B1(net571),
    .B2(net145),
    .A2(net573),
    .A1(\bp_core.addr_reg[9] ));
 sg13g2_o21ai_1 _2938_ (.B1(_1005_),
    .Y(_0033_),
    .A1(net573),
    .A2(net279));
 sg13g2_nand2_1 _2939_ (.Y(_1006_),
    .A(net742),
    .B(net336));
 sg13g2_a22oi_1 _2940_ (.Y(_1007_),
    .B1(net570),
    .B2(net64),
    .A2(net577),
    .A1(\bp_core.addr_reg[10] ));
 sg13g2_o21ai_1 _2941_ (.B1(_1007_),
    .Y(_0015_),
    .A1(net575),
    .A2(net337));
 sg13g2_nand2_1 _2942_ (.Y(_1008_),
    .A(net739),
    .B(net442));
 sg13g2_a22oi_1 _2943_ (.Y(_1009_),
    .B1(net569),
    .B2(\bp_core.bp_report_addr_out[11] ),
    .A2(net572),
    .A1(\bp_core.addr_reg[11] ));
 sg13g2_o21ai_1 _2944_ (.B1(_1009_),
    .Y(_0016_),
    .A1(net572),
    .A2(_1008_));
 sg13g2_nand2_1 _2945_ (.Y(_1010_),
    .A(net739),
    .B(net392));
 sg13g2_a22oi_1 _2946_ (.Y(_1011_),
    .B1(net569),
    .B2(net203),
    .A2(net572),
    .A1(\bp_core.addr_reg[12] ));
 sg13g2_o21ai_1 _2947_ (.B1(_1011_),
    .Y(_0017_),
    .A1(net572),
    .A2(_1010_));
 sg13g2_nand2_1 _2948_ (.Y(_1012_),
    .A(net740),
    .B(net254));
 sg13g2_a22oi_1 _2949_ (.Y(_1013_),
    .B1(net571),
    .B2(\bp_core.bp_report_addr_out[13] ),
    .A2(net573),
    .A1(\bp_core.addr_reg[13] ));
 sg13g2_o21ai_1 _2950_ (.B1(_1013_),
    .Y(_0018_),
    .A1(net573),
    .A2(net255));
 sg13g2_nand2_1 _2951_ (.Y(_1014_),
    .A(net739),
    .B(net414));
 sg13g2_a22oi_1 _2952_ (.Y(_1015_),
    .B1(net569),
    .B2(net275),
    .A2(net574),
    .A1(\bp_core.addr_reg[14] ));
 sg13g2_o21ai_1 _2953_ (.B1(_1015_),
    .Y(_0019_),
    .A1(net572),
    .A2(_1014_));
 sg13g2_nand2_1 _2954_ (.Y(_1016_),
    .A(net739),
    .B(net286));
 sg13g2_a22oi_1 _2955_ (.Y(_1017_),
    .B1(net569),
    .B2(\bp_core.bp_report_addr_out[15] ),
    .A2(net572),
    .A1(\bp_core.addr_reg[15] ));
 sg13g2_o21ai_1 _2956_ (.B1(_1017_),
    .Y(_0020_),
    .A1(net572),
    .A2(_1016_));
 sg13g2_nand2_1 _2957_ (.Y(_1018_),
    .A(net740),
    .B(\inter_bp.bp_report_addr_out[16] ));
 sg13g2_nor2_1 _2958_ (.A(net573),
    .B(_1018_),
    .Y(_1019_));
 sg13g2_a221oi_1 _2959_ (.B2(_0655_),
    .C1(_1019_),
    .B1(net569),
    .A1(_0546_),
    .Y(_0021_),
    .A2(net574));
 sg13g2_nand3_1 _2960_ (.B(\inter_bp.bp_report_addr_out[16] ),
    .C(\inter_bp.bp_report_addr_out[17] ),
    .A(net739),
    .Y(_1020_));
 sg13g2_o21ai_1 _2961_ (.B1(net739),
    .Y(_1021_),
    .A1(\inter_bp.bp_report_addr_out[16] ),
    .A2(\inter_bp.bp_report_addr_out[17] ));
 sg13g2_nand2b_1 _2962_ (.Y(_1022_),
    .B(_1020_),
    .A_N(_1021_));
 sg13g2_a22oi_1 _2963_ (.Y(_1023_),
    .B1(net569),
    .B2(net156),
    .A2(net572),
    .A1(net932));
 sg13g2_o21ai_1 _2964_ (.B1(_1023_),
    .Y(_0022_),
    .A1(net573),
    .A2(_1022_));
 sg13g2_nand4_1 _2965_ (.B(\inter_bp.bp_report_addr_out[16] ),
    .C(\inter_bp.bp_report_addr_out[17] ),
    .A(net739),
    .Y(_1024_),
    .D(\inter_bp.bp_report_addr_out[18] ));
 sg13g2_nand2_1 _2966_ (.Y(_1025_),
    .A(net739),
    .B(\inter_bp.bp_report_addr_out[18] ));
 sg13g2_nand2_1 _2967_ (.Y(_1026_),
    .A(_1020_),
    .B(_1025_));
 sg13g2_nand2_1 _2968_ (.Y(_1027_),
    .A(_1024_),
    .B(_1026_));
 sg13g2_a22oi_1 _2969_ (.Y(_1028_),
    .B1(net569),
    .B2(net972),
    .A2(net574),
    .A1(net482));
 sg13g2_o21ai_1 _2970_ (.B1(_1028_),
    .Y(_0023_),
    .A1(net574),
    .A2(_1027_));
 sg13g2_nand3_1 _2971_ (.B(net980),
    .C(_1024_),
    .A(net743),
    .Y(_1029_));
 sg13g2_a21oi_1 _2972_ (.A1(net743),
    .A2(net980),
    .Y(_1030_),
    .B1(_1024_));
 sg13g2_a21oi_1 _2973_ (.A1(net1121),
    .A2(_0973_),
    .Y(_1031_),
    .B1(_1030_));
 sg13g2_nand2_1 _2974_ (.Y(_1032_),
    .A(_1029_),
    .B(_1031_));
 sg13g2_mux2_1 _2975_ (.A0(net1122),
    .A1(net1092),
    .S(net574),
    .X(_0024_));
 sg13g2_o21ai_1 _2976_ (.B1(_0978_),
    .Y(_0038_),
    .A1(_0560_),
    .A2(_0034_));
 sg13g2_a21o_1 _2977_ (.A2(net571),
    .A1(net382),
    .B1(_0982_),
    .X(_0039_));
 sg13g2_o21ai_1 _2978_ (.B1(net334),
    .Y(_0040_),
    .A1(_0561_),
    .A2(_0034_));
 sg13g2_a21o_1 _2979_ (.A2(net570),
    .A1(net351),
    .B1(_0991_),
    .X(_0041_));
 sg13g2_a21o_1 _2980_ (.A2(net570),
    .A1(net405),
    .B1(net372),
    .X(_0042_));
 sg13g2_nor3_1 _2981_ (.A(\spi_ctrl.fsm_state[1] ),
    .B(\spi_ctrl.bits_remaining[3] ),
    .C(\spi_ctrl.bits_remaining[2] ),
    .Y(_1033_));
 sg13g2_a21oi_1 _2982_ (.A1(_0521_),
    .A2(\spi_ctrl.writing ),
    .Y(_1034_),
    .B1(\spi_ctrl.bits_remaining[1] ));
 sg13g2_nand3_1 _2983_ (.B(_1033_),
    .C(_1034_),
    .A(\spi_ctrl.fsm_state[0] ),
    .Y(_1035_));
 sg13g2_and2_1 _2984_ (.A(\spi_ctrl.fsm_state[1] ),
    .B(\spi_ctrl.fsm_state[0] ),
    .X(_1036_));
 sg13g2_nor2b_1 _2985_ (.A(\spi_ctrl.fsm_state[0] ),
    .B_N(\spi_ctrl.fsm_state[1] ),
    .Y(_1037_));
 sg13g2_a22oi_1 _2986_ (.Y(_1038_),
    .B1(net673),
    .B2(\spi_ctrl.addr[15] ),
    .A2(_1036_),
    .A1(\bp_core.ram_rdata[7] ));
 sg13g2_nand2_1 _2987_ (.Y(\spi_ctrl.spi_mosi ),
    .A(_1035_),
    .B(_1038_));
 sg13g2_nor2_1 _2988_ (.A(\bp_core.state[1] ),
    .B(\bp_core.state[5] ),
    .Y(_1039_));
 sg13g2_nor3_1 _2989_ (.A(_0687_),
    .B(net750),
    .C(_1039_),
    .Y(_1040_));
 sg13g2_a21oi_1 _2990_ (.A1(\bp_core.state[3] ),
    .A2(_0685_),
    .Y(_1041_),
    .B1(_1040_));
 sg13g2_inv_1 _2991_ (.Y(_1799_[0]),
    .A(net600));
 sg13g2_or2_1 _2992_ (.X(uo_out[1]),
    .B(\bp_core.valid_out ),
    .A(\bp_core.bp_param_output_valid ));
 sg13g2_nor2b_2 _2993_ (.A(net1083),
    .B_N(\bp_core.bp_param_valid_out ),
    .Y(_1042_));
 sg13g2_nor2_1 _2994_ (.A(\inter_bp.param_transmitting ),
    .B(net670),
    .Y(_1043_));
 sg13g2_nand2_1 _2995_ (.Y(_1044_),
    .A(net520),
    .B(\inter_bp.param_tx_counter[1] ));
 sg13g2_nand2_1 _2996_ (.Y(_1045_),
    .A(net270),
    .B(net1067));
 sg13g2_nor4_1 _2997_ (.A(net914),
    .B(net670),
    .C(_1044_),
    .D(_1045_),
    .Y(_1046_));
 sg13g2_nor2_1 _2998_ (.A(net642),
    .B(net1068),
    .Y(_0095_));
 sg13g2_nor2b_2 _2999_ (.A(\inter_bp.serialize_report_valid_prev ),
    .B_N(net57),
    .Y(_1047_));
 sg13g2_nor2_1 _3000_ (.A(net1114),
    .B(net660),
    .Y(_1048_));
 sg13g2_nand2b_1 _3001_ (.Y(_1049_),
    .B(net1007),
    .A_N(net1040));
 sg13g2_nand2b_1 _3002_ (.Y(_1050_),
    .B(net555),
    .A_N(net1079));
 sg13g2_nor4_1 _3003_ (.A(net325),
    .B(net660),
    .C(_1049_),
    .D(_1050_),
    .Y(_1051_));
 sg13g2_nor2_1 _3004_ (.A(net634),
    .B(_1051_),
    .Y(_0097_));
 sg13g2_a21oi_1 _3005_ (.A1(net720),
    .A2(_0548_),
    .Y(_1052_),
    .B1(net749));
 sg13g2_nor2b_1 _3006_ (.A(_0811_),
    .B_N(_1052_),
    .Y(_0035_));
 sg13g2_nor2_1 _3007_ (.A(net242),
    .B(net750),
    .Y(_0043_));
 sg13g2_nor3_1 _3008_ (.A(_0525_),
    .B(net359),
    .C(net749),
    .Y(_0037_));
 sg13g2_and3_1 _3009_ (.X(_0036_),
    .A(_0525_),
    .B(net1140),
    .C(_0713_));
 sg13g2_a21oi_1 _3010_ (.A1(net10),
    .A2(\inter_bp.param_receiving ),
    .Y(_1053_),
    .B1(_0945_));
 sg13g2_or2_1 _3011_ (.X(_1054_),
    .B(_1053_),
    .A(\inter_bp.param_rx_done ));
 sg13g2_a22oi_1 _3012_ (.Y(_1055_),
    .B1(net599),
    .B2(net397),
    .A2(net651),
    .A1(net926));
 sg13g2_inv_1 _3013_ (.Y(_0106_),
    .A(_1055_));
 sg13g2_a22oi_1 _3014_ (.Y(_1056_),
    .B1(net598),
    .B2(net408),
    .A2(net651),
    .A1(\inter_bp.param_shift_reg[3] ));
 sg13g2_inv_1 _3015_ (.Y(_0107_),
    .A(net409));
 sg13g2_a22oi_1 _3016_ (.Y(_1057_),
    .B1(net597),
    .B2(net926),
    .A2(net649),
    .A1(net534));
 sg13g2_inv_1 _3017_ (.Y(_0108_),
    .A(_1057_));
 sg13g2_a22oi_1 _3018_ (.Y(_1058_),
    .B1(net598),
    .B2(net904),
    .A2(net650),
    .A1(\inter_bp.param_shift_reg[5] ));
 sg13g2_inv_1 _3019_ (.Y(_0109_),
    .A(net905));
 sg13g2_a22oi_1 _3020_ (.Y(_1059_),
    .B1(net597),
    .B2(net534),
    .A2(net649),
    .A1(net493));
 sg13g2_inv_1 _3021_ (.Y(_0110_),
    .A(_1059_));
 sg13g2_a22oi_1 _3022_ (.Y(_1060_),
    .B1(net598),
    .B2(net927),
    .A2(net650),
    .A1(net907));
 sg13g2_inv_1 _3023_ (.Y(_0111_),
    .A(_1060_));
 sg13g2_a22oi_1 _3024_ (.Y(_1061_),
    .B1(net597),
    .B2(net493),
    .A2(net649),
    .A1(\inter_bp.param_shift_reg[8] ));
 sg13g2_inv_1 _3025_ (.Y(_0112_),
    .A(net494));
 sg13g2_a22oi_1 _3026_ (.Y(_1062_),
    .B1(net598),
    .B2(net907),
    .A2(net650),
    .A1(\inter_bp.param_shift_reg[9] ));
 sg13g2_inv_1 _3027_ (.Y(_0113_),
    .A(net908));
 sg13g2_a22oi_1 _3028_ (.Y(_1063_),
    .B1(net597),
    .B2(net934),
    .A2(net649),
    .A1(net891));
 sg13g2_inv_1 _3029_ (.Y(_0114_),
    .A(_1063_));
 sg13g2_a22oi_1 _3030_ (.Y(_1064_),
    .B1(net598),
    .B2(net920),
    .A2(net650),
    .A1(net533));
 sg13g2_inv_1 _3031_ (.Y(_0115_),
    .A(_1064_));
 sg13g2_a22oi_1 _3032_ (.Y(_1065_),
    .B1(net597),
    .B2(net891),
    .A2(net649),
    .A1(net853));
 sg13g2_inv_1 _3033_ (.Y(_0116_),
    .A(_1065_));
 sg13g2_a22oi_1 _3034_ (.Y(_1066_),
    .B1(net597),
    .B2(net533),
    .A2(net649),
    .A1(net484));
 sg13g2_inv_1 _3035_ (.Y(_0117_),
    .A(_1066_));
 sg13g2_a22oi_1 _3036_ (.Y(_1067_),
    .B1(net597),
    .B2(net853),
    .A2(net649),
    .A1(\inter_bp.param_shift_reg[14] ));
 sg13g2_inv_1 _3037_ (.Y(_0118_),
    .A(net854));
 sg13g2_a22oi_1 _3038_ (.Y(_1068_),
    .B1(net597),
    .B2(net484),
    .A2(net649),
    .A1(\inter_bp.param_shift_reg[15] ));
 sg13g2_inv_1 _3039_ (.Y(_0119_),
    .A(net485));
 sg13g2_a22oi_1 _3040_ (.Y(_1069_),
    .B1(net595),
    .B2(net1004),
    .A2(net647),
    .A1(net940));
 sg13g2_inv_1 _3041_ (.Y(_0120_),
    .A(_1069_));
 sg13g2_a22oi_1 _3042_ (.Y(_1070_),
    .B1(net595),
    .B2(net1005),
    .A2(net647),
    .A1(net529));
 sg13g2_inv_1 _3043_ (.Y(_0121_),
    .A(_1070_));
 sg13g2_a22oi_1 _3044_ (.Y(_1071_),
    .B1(net596),
    .B2(net940),
    .A2(net648),
    .A1(net888));
 sg13g2_inv_1 _3045_ (.Y(_0122_),
    .A(_1071_));
 sg13g2_a22oi_1 _3046_ (.Y(_1072_),
    .B1(net595),
    .B2(net529),
    .A2(net647),
    .A1(\inter_bp.param_shift_reg[19] ));
 sg13g2_inv_1 _3047_ (.Y(_0123_),
    .A(net530));
 sg13g2_a22oi_1 _3048_ (.Y(_1073_),
    .B1(net595),
    .B2(net888),
    .A2(net647),
    .A1(\inter_bp.param_shift_reg[20] ));
 sg13g2_inv_1 _3049_ (.Y(_0124_),
    .A(net889));
 sg13g2_a22oi_1 _3050_ (.Y(_1074_),
    .B1(net592),
    .B2(net882),
    .A2(net646),
    .A1(net856));
 sg13g2_inv_1 _3051_ (.Y(_0125_),
    .A(_1074_));
 sg13g2_a22oi_1 _3052_ (.Y(_1075_),
    .B1(net599),
    .B2(net942),
    .A2(net651),
    .A1(net444));
 sg13g2_inv_1 _3053_ (.Y(_0126_),
    .A(_1075_));
 sg13g2_a22oi_1 _3054_ (.Y(_1076_),
    .B1(net592),
    .B2(net856),
    .A2(net646),
    .A1(net935));
 sg13g2_inv_1 _3055_ (.Y(_0127_),
    .A(_1076_));
 sg13g2_a22oi_1 _3056_ (.Y(_1077_),
    .B1(net599),
    .B2(net444),
    .A2(net651),
    .A1(\inter_bp.param_shift_reg[24] ));
 sg13g2_inv_1 _3057_ (.Y(_0128_),
    .A(net445));
 sg13g2_a22oi_1 _3058_ (.Y(_1078_),
    .B1(net592),
    .B2(net935),
    .A2(net643),
    .A1(net429));
 sg13g2_inv_1 _3059_ (.Y(_0129_),
    .A(_1078_));
 sg13g2_a22oi_1 _3060_ (.Y(_1079_),
    .B1(net599),
    .B2(net881),
    .A2(net651),
    .A1(net498));
 sg13g2_inv_1 _3061_ (.Y(_0130_),
    .A(_1079_));
 sg13g2_a22oi_1 _3062_ (.Y(_1080_),
    .B1(net591),
    .B2(net429),
    .A2(net643),
    .A1(\inter_bp.param_shift_reg[27] ));
 sg13g2_inv_1 _3063_ (.Y(_0131_),
    .A(net430));
 sg13g2_a22oi_1 _3064_ (.Y(_1081_),
    .B1(net599),
    .B2(net498),
    .A2(net651),
    .A1(\inter_bp.param_shift_reg[28] ));
 sg13g2_inv_1 _3065_ (.Y(_0132_),
    .A(net499));
 sg13g2_a22oi_1 _3066_ (.Y(_1082_),
    .B1(net591),
    .B2(net451),
    .A2(net643),
    .A1(\inter_bp.param_shift_reg[29] ));
 sg13g2_inv_1 _3067_ (.Y(_0133_),
    .A(net452));
 sg13g2_a22oi_1 _3068_ (.Y(_1083_),
    .B1(net599),
    .B2(net525),
    .A2(net651),
    .A1(\inter_bp.param_shift_reg[30] ));
 sg13g2_inv_1 _3069_ (.Y(_0134_),
    .A(net526));
 sg13g2_a22oi_1 _3070_ (.Y(_1084_),
    .B1(net591),
    .B2(net961),
    .A2(net643),
    .A1(net427));
 sg13g2_inv_1 _3071_ (.Y(_0135_),
    .A(_1084_));
 sg13g2_a22oi_1 _3072_ (.Y(_1085_),
    .B1(net595),
    .B2(net849),
    .A2(net647),
    .A1(\inter_bp.param_shift_reg[32] ));
 sg13g2_inv_1 _3073_ (.Y(_0136_),
    .A(net850));
 sg13g2_a22oi_1 _3074_ (.Y(_1086_),
    .B1(net591),
    .B2(net427),
    .A2(net643),
    .A1(net898));
 sg13g2_inv_1 _3075_ (.Y(_0137_),
    .A(_1086_));
 sg13g2_a22oi_1 _3076_ (.Y(_1087_),
    .B1(net595),
    .B2(net866),
    .A2(net647),
    .A1(\inter_bp.param_shift_reg[34] ));
 sg13g2_inv_1 _3077_ (.Y(_0138_),
    .A(net867));
 sg13g2_a22oi_1 _3078_ (.Y(_1088_),
    .B1(net592),
    .B2(net898),
    .A2(net643),
    .A1(\inter_bp.param_shift_reg[35] ));
 sg13g2_inv_1 _3079_ (.Y(_0139_),
    .A(net899));
 sg13g2_a22oi_1 _3080_ (.Y(_1089_),
    .B1(net595),
    .B2(net921),
    .A2(net647),
    .A1(net515));
 sg13g2_inv_1 _3081_ (.Y(_0140_),
    .A(_1089_));
 sg13g2_a22oi_1 _3082_ (.Y(_1090_),
    .B1(net593),
    .B2(net912),
    .A2(net644),
    .A1(\inter_bp.param_shift_reg[37] ));
 sg13g2_inv_1 _3083_ (.Y(_0141_),
    .A(net913));
 sg13g2_a22oi_1 _3084_ (.Y(_1091_),
    .B1(net595),
    .B2(net515),
    .A2(net647),
    .A1(net462));
 sg13g2_inv_1 _3085_ (.Y(_0142_),
    .A(_1091_));
 sg13g2_a22oi_1 _3086_ (.Y(_1092_),
    .B1(net593),
    .B2(net948),
    .A2(net644),
    .A1(net939));
 sg13g2_inv_1 _3087_ (.Y(_0143_),
    .A(_1092_));
 sg13g2_a22oi_1 _3088_ (.Y(_1093_),
    .B1(net596),
    .B2(net462),
    .A2(net648),
    .A1(\inter_bp.param_shift_reg[40] ));
 sg13g2_inv_1 _3089_ (.Y(_0144_),
    .A(net463));
 sg13g2_a22oi_1 _3090_ (.Y(_1094_),
    .B1(net593),
    .B2(net939),
    .A2(net644),
    .A1(net349));
 sg13g2_inv_1 _3091_ (.Y(_0145_),
    .A(_1094_));
 sg13g2_a22oi_1 _3092_ (.Y(_1095_),
    .B1(net594),
    .B2(net945),
    .A2(net645),
    .A1(net971));
 sg13g2_inv_1 _3093_ (.Y(_0146_),
    .A(_1095_));
 sg13g2_a22oi_1 _3094_ (.Y(_1096_),
    .B1(net594),
    .B2(net349),
    .A2(net644),
    .A1(net862));
 sg13g2_inv_1 _3095_ (.Y(_0147_),
    .A(_1096_));
 sg13g2_a22oi_1 _3096_ (.Y(_1097_),
    .B1(net594),
    .B2(net971),
    .A2(net645),
    .A1(net917));
 sg13g2_inv_1 _3097_ (.Y(_0148_),
    .A(_1097_));
 sg13g2_a22oi_1 _3098_ (.Y(_1098_),
    .B1(net593),
    .B2(net862),
    .A2(net645),
    .A1(net886));
 sg13g2_inv_1 _3099_ (.Y(_0149_),
    .A(_1098_));
 sg13g2_a22oi_1 _3100_ (.Y(_1099_),
    .B1(net593),
    .B2(net917),
    .A2(net645),
    .A1(\inter_bp.param_shift_reg[46] ));
 sg13g2_inv_1 _3101_ (.Y(_0150_),
    .A(net918));
 sg13g2_a22oi_1 _3102_ (.Y(_1100_),
    .B1(net593),
    .B2(net886),
    .A2(net644),
    .A1(net910));
 sg13g2_inv_1 _3103_ (.Y(_0151_),
    .A(_1100_));
 sg13g2_mux2_1 _3104_ (.A0(net12),
    .A1(net992),
    .S(net593),
    .X(_0152_));
 sg13g2_mux2_1 _3105_ (.A0(net13),
    .A1(net910),
    .S(net593),
    .X(_0153_));
 sg13g2_nand2b_1 _3106_ (.Y(_1101_),
    .B(net11),
    .A_N(net461));
 sg13g2_nor2_2 _3107_ (.A(net746),
    .B(_1101_),
    .Y(_1102_));
 sg13g2_nor2_1 _3108_ (.A(_0952_),
    .B(_1102_),
    .Y(_1103_));
 sg13g2_nor3_1 _3109_ (.A(net308),
    .B(_0952_),
    .C(_1102_),
    .Y(_1104_));
 sg13g2_a21oi_1 _3110_ (.A1(net308),
    .A2(net608),
    .Y(_0154_),
    .B1(_1104_));
 sg13g2_xor2_1 _3111_ (.B(net308),
    .A(net1086),
    .X(_1105_));
 sg13g2_a22oi_1 _3112_ (.Y(_1106_),
    .B1(_1105_),
    .B2(net608),
    .A2(net589),
    .A1(net1086));
 sg13g2_inv_1 _3113_ (.Y(_0155_),
    .A(_1106_));
 sg13g2_nand3b_1 _3114_ (.B(net308),
    .C(net1086),
    .Y(_1107_),
    .A_N(net590));
 sg13g2_nor2_1 _3115_ (.A(_0557_),
    .B(_1107_),
    .Y(_1108_));
 sg13g2_a21oi_1 _3116_ (.A1(_0557_),
    .A2(_1107_),
    .Y(_1109_),
    .B1(_1102_));
 sg13g2_nor2b_1 _3117_ (.A(_1108_),
    .B_N(_1109_),
    .Y(_0156_));
 sg13g2_nand4_1 _3118_ (.B(net308),
    .C(\inter_bp.report_rx_counter[2] ),
    .A(\inter_bp.report_rx_counter[1] ),
    .Y(_1110_),
    .D(net448));
 sg13g2_a21oi_1 _3119_ (.A1(_1101_),
    .A2(_1110_),
    .Y(_1111_),
    .B1(net590));
 sg13g2_nor2_1 _3120_ (.A(net448),
    .B(_1108_),
    .Y(_1112_));
 sg13g2_nor2_1 _3121_ (.A(_1111_),
    .B(net449),
    .Y(_0157_));
 sg13g2_nand2b_1 _3122_ (.Y(_1113_),
    .B(net322),
    .A_N(_1111_));
 sg13g2_nand2b_1 _3123_ (.Y(_1114_),
    .B(net607),
    .A_N(net322));
 sg13g2_o21ai_1 _3124_ (.B1(net323),
    .Y(_0158_),
    .A1(_1110_),
    .A2(_1114_));
 sg13g2_a22oi_1 _3125_ (.Y(_1115_),
    .B1(net589),
    .B2(net257),
    .A2(net607),
    .A1(\inter_bp.report_shift_reg[2] ));
 sg13g2_inv_1 _3126_ (.Y(_0159_),
    .A(net258));
 sg13g2_a22oi_1 _3127_ (.Y(_1116_),
    .B1(net589),
    .B2(net273),
    .A2(net607),
    .A1(\inter_bp.report_shift_reg[3] ));
 sg13g2_inv_1 _3128_ (.Y(_0160_),
    .A(net274));
 sg13g2_a22oi_1 _3129_ (.Y(_1117_),
    .B1(net589),
    .B2(net410),
    .A2(net607),
    .A1(\inter_bp.report_shift_reg[4] ));
 sg13g2_inv_1 _3130_ (.Y(_0161_),
    .A(net411));
 sg13g2_a22oi_1 _3131_ (.Y(_1118_),
    .B1(net589),
    .B2(net486),
    .A2(net607),
    .A1(\inter_bp.report_shift_reg[5] ));
 sg13g2_inv_1 _3132_ (.Y(_0162_),
    .A(net487));
 sg13g2_a22oi_1 _3133_ (.Y(_1119_),
    .B1(net589),
    .B2(net858),
    .A2(net607),
    .A1(net426));
 sg13g2_inv_1 _3134_ (.Y(_0163_),
    .A(_1119_));
 sg13g2_a22oi_1 _3135_ (.Y(_1120_),
    .B1(net588),
    .B2(net504),
    .A2(net606),
    .A1(net539));
 sg13g2_inv_1 _3136_ (.Y(_0164_),
    .A(_1120_));
 sg13g2_a22oi_1 _3137_ (.Y(_1121_),
    .B1(net589),
    .B2(net426),
    .A2(net607),
    .A1(net386));
 sg13g2_inv_1 _3138_ (.Y(_0165_),
    .A(_1121_));
 sg13g2_a22oi_1 _3139_ (.Y(_1122_),
    .B1(net588),
    .B2(net539),
    .A2(net608),
    .A1(net418));
 sg13g2_inv_1 _3140_ (.Y(_0166_),
    .A(_1122_));
 sg13g2_a22oi_1 _3141_ (.Y(_1123_),
    .B1(net589),
    .B2(net386),
    .A2(net607),
    .A1(\inter_bp.report_shift_reg[10] ));
 sg13g2_inv_1 _3142_ (.Y(_0167_),
    .A(net387));
 sg13g2_a22oi_1 _3143_ (.Y(_1124_),
    .B1(net588),
    .B2(net418),
    .A2(net608),
    .A1(\inter_bp.report_shift_reg[11] ));
 sg13g2_inv_1 _3144_ (.Y(_0168_),
    .A(net419));
 sg13g2_a22oi_1 _3145_ (.Y(_1125_),
    .B1(net588),
    .B2(net431),
    .A2(net608),
    .A1(\inter_bp.report_shift_reg[12] ));
 sg13g2_inv_1 _3146_ (.Y(_0169_),
    .A(net432));
 sg13g2_a22oi_1 _3147_ (.Y(_1126_),
    .B1(net587),
    .B2(net447),
    .A2(net606),
    .A1(net376));
 sg13g2_inv_1 _3148_ (.Y(_0170_),
    .A(_1126_));
 sg13g2_a22oi_1 _3149_ (.Y(_1127_),
    .B1(net587),
    .B2(net893),
    .A2(net606),
    .A1(net403));
 sg13g2_inv_1 _3150_ (.Y(_0171_),
    .A(_1127_));
 sg13g2_a22oi_1 _3151_ (.Y(_1128_),
    .B1(net587),
    .B2(net376),
    .A2(net606),
    .A1(\inter_bp.report_shift_reg[15] ));
 sg13g2_inv_1 _3152_ (.Y(_0172_),
    .A(net377));
 sg13g2_a22oi_1 _3153_ (.Y(_1129_),
    .B1(net587),
    .B2(net403),
    .A2(net606),
    .A1(\inter_bp.report_shift_reg[16] ));
 sg13g2_inv_1 _3154_ (.Y(_0173_),
    .A(net404));
 sg13g2_a22oi_1 _3155_ (.Y(_1130_),
    .B1(net587),
    .B2(net435),
    .A2(net606),
    .A1(net374));
 sg13g2_inv_1 _3156_ (.Y(_0174_),
    .A(_1130_));
 sg13g2_a22oi_1 _3157_ (.Y(_1131_),
    .B1(net587),
    .B2(net437),
    .A2(net606),
    .A1(\inter_bp.report_shift_reg[18] ));
 sg13g2_inv_1 _3158_ (.Y(_0175_),
    .A(net438));
 sg13g2_a22oi_1 _3159_ (.Y(_1132_),
    .B1(net587),
    .B2(net374),
    .A2(net606),
    .A1(\inter_bp.report_shift_reg[19] ));
 sg13g2_inv_1 _3160_ (.Y(_0176_),
    .A(net375));
 sg13g2_mux2_1 _3161_ (.A0(net12),
    .A1(net1001),
    .S(net587),
    .X(_0177_));
 sg13g2_mux2_1 _3162_ (.A0(net13),
    .A1(net1027),
    .S(net588),
    .X(_0178_));
 sg13g2_mux2_1 _3163_ (.A0(net535),
    .A1(net257),
    .S(net747),
    .X(_0179_));
 sg13g2_mux2_1 _3164_ (.A0(net401),
    .A1(net273),
    .S(net746),
    .X(_0180_));
 sg13g2_mux2_1 _3165_ (.A0(net998),
    .A1(net410),
    .S(net747),
    .X(_0181_));
 sg13g2_mux2_1 _3166_ (.A0(net439),
    .A1(\inter_bp.report_shift_reg[3] ),
    .S(net746),
    .X(_0182_));
 sg13g2_mux2_1 _3167_ (.A0(net892),
    .A1(net858),
    .S(net747),
    .X(_0183_));
 sg13g2_mux2_1 _3168_ (.A0(net281),
    .A1(net504),
    .S(net745),
    .X(_0184_));
 sg13g2_mux2_1 _3169_ (.A0(net328),
    .A1(net426),
    .S(net746),
    .X(_0185_));
 sg13g2_mux2_1 _3170_ (.A0(net261),
    .A1(net539),
    .S(net745),
    .X(_0186_));
 sg13g2_mux2_1 _3171_ (.A0(net298),
    .A1(net386),
    .S(net746),
    .X(_0187_));
 sg13g2_mux2_1 _3172_ (.A0(net278),
    .A1(net418),
    .S(net745),
    .X(_0188_));
 sg13g2_mux2_1 _3173_ (.A0(net336),
    .A1(net431),
    .S(net746),
    .X(_0189_));
 sg13g2_mux2_1 _3174_ (.A0(net442),
    .A1(net447),
    .S(net744),
    .X(_0190_));
 sg13g2_mux2_1 _3175_ (.A0(net392),
    .A1(net893),
    .S(net744),
    .X(_0191_));
 sg13g2_mux2_1 _3176_ (.A0(net254),
    .A1(net376),
    .S(net745),
    .X(_0192_));
 sg13g2_mux2_1 _3177_ (.A0(net414),
    .A1(net403),
    .S(net744),
    .X(_0193_));
 sg13g2_mux2_1 _3178_ (.A0(net286),
    .A1(net435),
    .S(net744),
    .X(_0194_));
 sg13g2_mux2_1 _3179_ (.A0(net1003),
    .A1(net437),
    .S(net744),
    .X(_0195_));
 sg13g2_mux2_1 _3180_ (.A0(net990),
    .A1(net374),
    .S(net744),
    .X(_0196_));
 sg13g2_mux2_1 _3181_ (.A0(\inter_bp.bp_report_addr_out[18] ),
    .A1(net1001),
    .S(net744),
    .X(_0197_));
 sg13g2_mux2_1 _3182_ (.A0(net980),
    .A1(\inter_bp.report_shift_reg[19] ),
    .S(net744),
    .X(_0198_));
 sg13g2_a21oi_1 _3183_ (.A1(_0954_),
    .A2(net1064),
    .Y(_1133_),
    .B1(_0951_));
 sg13g2_a21oi_1 _3184_ (.A1(net746),
    .A2(net855),
    .Y(_1134_),
    .B1(_1102_));
 sg13g2_nand2b_1 _3185_ (.Y(_0199_),
    .B(_1134_),
    .A_N(_1133_));
 sg13g2_nor2_1 _3186_ (.A(\inter_bp.param_transmitting ),
    .B(net520),
    .Y(_1135_));
 sg13g2_and2_1 _3187_ (.A(\inter_bp.param_transmitting ),
    .B(net520),
    .X(_1136_));
 sg13g2_nor3_1 _3188_ (.A(net670),
    .B(net521),
    .C(_1136_),
    .Y(_0200_));
 sg13g2_a21oi_1 _3189_ (.A1(net1084),
    .A2(_1136_),
    .Y(_1137_),
    .B1(net670));
 sg13g2_o21ai_1 _3190_ (.B1(_1137_),
    .Y(_1138_),
    .A1(net1084),
    .A2(_1136_));
 sg13g2_inv_1 _3191_ (.Y(_0201_),
    .A(net1085));
 sg13g2_a21oi_1 _3192_ (.A1(\inter_bp.param_tx_counter[1] ),
    .A2(_1136_),
    .Y(_1139_),
    .B1(net270));
 sg13g2_and3_1 _3193_ (.X(_1140_),
    .A(net1182),
    .B(net270),
    .C(_1136_));
 sg13g2_nor3_1 _3194_ (.A(net670),
    .B(net271),
    .C(_1140_),
    .Y(_0202_));
 sg13g2_nor2_1 _3195_ (.A(net914),
    .B(_1140_),
    .Y(_1141_));
 sg13g2_and2_1 _3196_ (.A(net914),
    .B(_1140_),
    .X(_1142_));
 sg13g2_nor3_1 _3197_ (.A(net670),
    .B(net915),
    .C(_1142_),
    .Y(_0203_));
 sg13g2_a21oi_1 _3198_ (.A1(net1067),
    .A2(_1142_),
    .Y(_1143_),
    .B1(net670));
 sg13g2_o21ai_1 _3199_ (.B1(_1143_),
    .Y(_1144_),
    .A1(net1067),
    .A2(_1142_));
 sg13g2_inv_1 _3200_ (.Y(_0204_),
    .A(_1144_));
 sg13g2_nand2_1 _3201_ (.Y(_1145_),
    .A(net288),
    .B(_0948_));
 sg13g2_o21ai_1 _3202_ (.B1(_1145_),
    .Y(_0205_),
    .A1(net288),
    .A2(net591));
 sg13g2_xor2_1 _3203_ (.B(net288),
    .A(net965),
    .X(_1146_));
 sg13g2_a22oi_1 _3204_ (.Y(_1147_),
    .B1(_1146_),
    .B2(net643),
    .A2(net591),
    .A1(net965));
 sg13g2_inv_1 _3205_ (.Y(_0206_),
    .A(_1147_));
 sg13g2_a21oi_1 _3206_ (.A1(net965),
    .A2(net288),
    .Y(_1148_),
    .B1(net395));
 sg13g2_nor2_1 _3207_ (.A(net396),
    .B(_1148_),
    .Y(_1149_));
 sg13g2_a22oi_1 _3208_ (.Y(_1150_),
    .B1(_1149_),
    .B2(net643),
    .A2(net591),
    .A1(net395));
 sg13g2_inv_1 _3209_ (.Y(_0207_),
    .A(_1150_));
 sg13g2_nand2_1 _3210_ (.Y(_1151_),
    .A(net318),
    .B(_0949_));
 sg13g2_a21oi_1 _3211_ (.A1(net644),
    .A2(_1151_),
    .Y(_1152_),
    .B1(net591));
 sg13g2_a21oi_1 _3212_ (.A1(net644),
    .A2(_0949_),
    .Y(_1153_),
    .B1(net318));
 sg13g2_nor2_1 _3213_ (.A(_1152_),
    .B(net319),
    .Y(_0208_));
 sg13g2_nand4_1 _3214_ (.B(_0559_),
    .C(net644),
    .A(net318),
    .Y(_1154_),
    .D(net396));
 sg13g2_o21ai_1 _3215_ (.B1(_1154_),
    .Y(_0209_),
    .A1(_0559_),
    .A2(_1152_));
 sg13g2_nand2_1 _3216_ (.Y(_1155_),
    .A(net159),
    .B(net642));
 sg13g2_nor2b_2 _3217_ (.A(net670),
    .B_N(\inter_bp.param_transmitting ),
    .Y(_1156_));
 sg13g2_a22oi_1 _3218_ (.Y(_1157_),
    .B1(net628),
    .B2(\inter_bp.param_tx_shift_reg[2] ),
    .A2(net665),
    .A1(\bp_addr_out[0] ));
 sg13g2_nand2_1 _3219_ (.Y(_0210_),
    .A(net160),
    .B(_1157_));
 sg13g2_nand2_1 _3220_ (.Y(_1158_),
    .A(net179),
    .B(net642));
 sg13g2_a22oi_1 _3221_ (.Y(_1159_),
    .B1(net628),
    .B2(\inter_bp.param_tx_shift_reg[3] ),
    .A2(net665),
    .A1(\bp_addr_out[1] ));
 sg13g2_nand2_1 _3222_ (.Y(_0211_),
    .A(net180),
    .B(_1159_));
 sg13g2_nand2_1 _3223_ (.Y(_1160_),
    .A(net232),
    .B(net640));
 sg13g2_a22oi_1 _3224_ (.Y(_1161_),
    .B1(net629),
    .B2(\inter_bp.param_tx_shift_reg[4] ),
    .A2(net666),
    .A1(\bp_addr_out[2] ));
 sg13g2_nand2_1 _3225_ (.Y(_0212_),
    .A(_1160_),
    .B(_1161_));
 sg13g2_nand2_1 _3226_ (.Y(_1162_),
    .A(net243),
    .B(net640));
 sg13g2_a22oi_1 _3227_ (.Y(_1163_),
    .B1(net631),
    .B2(net217),
    .A2(net668),
    .A1(\bp_addr_out[3] ));
 sg13g2_nand2_1 _3228_ (.Y(_0213_),
    .A(_1162_),
    .B(_1163_));
 sg13g2_nand2_1 _3229_ (.Y(_1164_),
    .A(net301),
    .B(net641));
 sg13g2_a22oi_1 _3230_ (.Y(_1165_),
    .B1(_1156_),
    .B2(net268),
    .A2(net669),
    .A1(\bp_addr_out[4] ));
 sg13g2_nand2_1 _3231_ (.Y(_0214_),
    .A(_1164_),
    .B(_1165_));
 sg13g2_nand2_1 _3232_ (.Y(_1166_),
    .A(net100),
    .B(net631));
 sg13g2_a22oi_1 _3233_ (.Y(_1167_),
    .B1(net641),
    .B2(net217),
    .A2(net668),
    .A1(\bp_addr_out[5] ));
 sg13g2_nand2_1 _3234_ (.Y(_0215_),
    .A(_1166_),
    .B(net218));
 sg13g2_nand2_1 _3235_ (.Y(_1168_),
    .A(net268),
    .B(net641));
 sg13g2_a22oi_1 _3236_ (.Y(_1169_),
    .B1(net631),
    .B2(net245),
    .A2(net668),
    .A1(\bp_addr_out[6] ));
 sg13g2_nand2_1 _3237_ (.Y(_0216_),
    .A(_1168_),
    .B(_1169_));
 sg13g2_nand2_1 _3238_ (.Y(_1170_),
    .A(net100),
    .B(net639));
 sg13g2_a22oi_1 _3239_ (.Y(_1171_),
    .B1(net631),
    .B2(\inter_bp.param_tx_shift_reg[9] ),
    .A2(net668),
    .A1(\bp_addr_out[7] ));
 sg13g2_nand2_1 _3240_ (.Y(_0217_),
    .A(_1170_),
    .B(_1171_));
 sg13g2_nand2_1 _3241_ (.Y(_1172_),
    .A(net103),
    .B(net630));
 sg13g2_a22oi_1 _3242_ (.Y(_1173_),
    .B1(net639),
    .B2(net245),
    .A2(net669),
    .A1(\bp_addr_out[8] ));
 sg13g2_nand2_1 _3243_ (.Y(_0218_),
    .A(_1172_),
    .B(net246));
 sg13g2_nand2_1 _3244_ (.Y(_1174_),
    .A(net105),
    .B(net630));
 sg13g2_a22oi_1 _3245_ (.Y(_1175_),
    .B1(net639),
    .B2(net211),
    .A2(net667),
    .A1(\bp_addr_out[9] ));
 sg13g2_nand2_1 _3246_ (.Y(_0219_),
    .A(_1174_),
    .B(net212));
 sg13g2_nand2_1 _3247_ (.Y(_1176_),
    .A(net86),
    .B(net630));
 sg13g2_a22oi_1 _3248_ (.Y(_1177_),
    .B1(net639),
    .B2(net103),
    .A2(net668),
    .A1(\bp_addr_out[10] ));
 sg13g2_nand2_1 _3249_ (.Y(_0220_),
    .A(_1176_),
    .B(net104));
 sg13g2_nand2_1 _3250_ (.Y(_1178_),
    .A(net105),
    .B(net639));
 sg13g2_a22oi_1 _3251_ (.Y(_1179_),
    .B1(net630),
    .B2(\inter_bp.param_tx_shift_reg[13] ),
    .A2(net667),
    .A1(\bp_addr_out[11] ));
 sg13g2_nand2_1 _3252_ (.Y(_0221_),
    .A(_1178_),
    .B(_1179_));
 sg13g2_nand2_1 _3253_ (.Y(_1180_),
    .A(net80),
    .B(net631));
 sg13g2_a22oi_1 _3254_ (.Y(_1181_),
    .B1(net639),
    .B2(net86),
    .A2(net667),
    .A1(\bp_addr_out[12] ));
 sg13g2_nand2_1 _3255_ (.Y(_0222_),
    .A(_1180_),
    .B(net87));
 sg13g2_nand2_1 _3256_ (.Y(_1182_),
    .A(net60),
    .B(net631));
 sg13g2_a22oi_1 _3257_ (.Y(_1183_),
    .B1(net639),
    .B2(\inter_bp.param_tx_shift_reg[13] ),
    .A2(net668),
    .A1(\bp_addr_out[13] ));
 sg13g2_nand2_1 _3258_ (.Y(_0223_),
    .A(_1182_),
    .B(_1183_));
 sg13g2_nand2_1 _3259_ (.Y(_1184_),
    .A(net72),
    .B(net631));
 sg13g2_a22oi_1 _3260_ (.Y(_1185_),
    .B1(net638),
    .B2(net80),
    .A2(net668),
    .A1(\bp_addr_out[14] ));
 sg13g2_nand2_1 _3261_ (.Y(_0224_),
    .A(_1184_),
    .B(net81));
 sg13g2_nand2_1 _3262_ (.Y(_1186_),
    .A(net60),
    .B(net638));
 sg13g2_a22oi_1 _3263_ (.Y(_1187_),
    .B1(net627),
    .B2(net88),
    .A2(net663),
    .A1(\bp_addr_out[15] ));
 sg13g2_nand2_1 _3264_ (.Y(_0225_),
    .A(_1186_),
    .B(net89));
 sg13g2_nand2_1 _3265_ (.Y(_1188_),
    .A(net72),
    .B(net638));
 sg13g2_a22oi_1 _3266_ (.Y(_1189_),
    .B1(net625),
    .B2(\inter_bp.param_tx_shift_reg[18] ),
    .A2(net664),
    .A1(\bp_addr_out[16] ));
 sg13g2_nand2_1 _3267_ (.Y(_0226_),
    .A(_1188_),
    .B(_1189_));
 sg13g2_nand2_1 _3268_ (.Y(_1190_),
    .A(net88),
    .B(net635));
 sg13g2_a22oi_1 _3269_ (.Y(_1191_),
    .B1(net626),
    .B2(net78),
    .A2(net663),
    .A1(net102));
 sg13g2_nand2_1 _3270_ (.Y(_0227_),
    .A(_1190_),
    .B(_1191_));
 sg13g2_nand2_1 _3271_ (.Y(_1192_),
    .A(net190),
    .B(net635));
 sg13g2_a22oi_1 _3272_ (.Y(_1193_),
    .B1(net625),
    .B2(net137),
    .A2(net664),
    .A1(\bp_addr_out[18] ));
 sg13g2_nand2_1 _3273_ (.Y(_0228_),
    .A(_1192_),
    .B(_1193_));
 sg13g2_nand2_1 _3274_ (.Y(_1194_),
    .A(net78),
    .B(net635));
 sg13g2_a22oi_1 _3275_ (.Y(_1195_),
    .B1(net626),
    .B2(\inter_bp.param_tx_shift_reg[21] ),
    .A2(net663),
    .A1(\bp_addr_out[19] ));
 sg13g2_nand2_1 _3276_ (.Y(_0229_),
    .A(_1194_),
    .B(_1195_));
 sg13g2_nand2_1 _3277_ (.Y(_1196_),
    .A(net137),
    .B(net636));
 sg13g2_a22oi_1 _3278_ (.Y(_1197_),
    .B1(net625),
    .B2(\inter_bp.param_tx_shift_reg[22] ),
    .A2(net664),
    .A1(\bp_core.bp_stride_out[0] ));
 sg13g2_nand2_1 _3279_ (.Y(_0230_),
    .A(_1196_),
    .B(_1197_));
 sg13g2_nand2_1 _3280_ (.Y(_1198_),
    .A(net67),
    .B(net625));
 sg13g2_a22oi_1 _3281_ (.Y(_1199_),
    .B1(net636),
    .B2(net84),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[1] ));
 sg13g2_nand2_1 _3282_ (.Y(_0231_),
    .A(_1198_),
    .B(net85));
 sg13g2_nand2_1 _3283_ (.Y(_1200_),
    .A(net221),
    .B(net635));
 sg13g2_a22oi_1 _3284_ (.Y(_1201_),
    .B1(net626),
    .B2(net206),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[2] ));
 sg13g2_nand2_1 _3285_ (.Y(_0232_),
    .A(_1200_),
    .B(_1201_));
 sg13g2_nand2_1 _3286_ (.Y(_1202_),
    .A(net67),
    .B(net636));
 sg13g2_a22oi_1 _3287_ (.Y(_1203_),
    .B1(net625),
    .B2(\inter_bp.param_tx_shift_reg[25] ),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[3] ));
 sg13g2_nand2_1 _3288_ (.Y(_0233_),
    .A(_1202_),
    .B(_1203_));
 sg13g2_nand2_1 _3289_ (.Y(_1204_),
    .A(net162),
    .B(net630));
 sg13g2_a22oi_1 _3290_ (.Y(_1205_),
    .B1(net638),
    .B2(net206),
    .A2(net667),
    .A1(\bp_core.bp_stride_out[4] ));
 sg13g2_nand2_1 _3291_ (.Y(_0234_),
    .A(_1204_),
    .B(net207));
 sg13g2_nand2_1 _3292_ (.Y(_1206_),
    .A(net62),
    .B(net627));
 sg13g2_a22oi_1 _3293_ (.Y(_1207_),
    .B1(net636),
    .B2(\inter_bp.param_tx_shift_reg[25] ),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[5] ));
 sg13g2_nand2_1 _3294_ (.Y(_0235_),
    .A(_1206_),
    .B(_1207_));
 sg13g2_nand2_1 _3295_ (.Y(_1208_),
    .A(net162),
    .B(net638));
 sg13g2_a22oi_1 _3296_ (.Y(_1209_),
    .B1(net630),
    .B2(net129),
    .A2(net667),
    .A1(\bp_core.bp_stride_out[6] ));
 sg13g2_nand2_1 _3297_ (.Y(_0236_),
    .A(_1208_),
    .B(_1209_));
 sg13g2_nand2_1 _3298_ (.Y(_1210_),
    .A(net62),
    .B(net637));
 sg13g2_a22oi_1 _3299_ (.Y(_1211_),
    .B1(net627),
    .B2(net200),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[7] ));
 sg13g2_nand2_1 _3300_ (.Y(_0237_),
    .A(_1210_),
    .B(net201));
 sg13g2_nand2_1 _3301_ (.Y(_1212_),
    .A(net98),
    .B(net630));
 sg13g2_a22oi_1 _3302_ (.Y(_1213_),
    .B1(net638),
    .B2(net129),
    .A2(net667),
    .A1(\bp_core.bp_stride_out[8] ));
 sg13g2_nand2_1 _3303_ (.Y(_0238_),
    .A(_1212_),
    .B(net130));
 sg13g2_nand2_1 _3304_ (.Y(_1214_),
    .A(net139),
    .B(net627));
 sg13g2_a22oi_1 _3305_ (.Y(_1215_),
    .B1(net636),
    .B2(net200),
    .A2(net663),
    .A1(net202));
 sg13g2_nand2_1 _3306_ (.Y(_0239_),
    .A(_1214_),
    .B(_1215_));
 sg13g2_nand2_1 _3307_ (.Y(_1216_),
    .A(net98),
    .B(net638));
 sg13g2_a22oi_1 _3308_ (.Y(_1217_),
    .B1(net630),
    .B2(net82),
    .A2(net667),
    .A1(\bp_core.bp_stride_out[10] ));
 sg13g2_nand2_1 _3309_ (.Y(_0240_),
    .A(_1216_),
    .B(_1217_));
 sg13g2_nand2_1 _3310_ (.Y(_1218_),
    .A(net139),
    .B(net637));
 sg13g2_a22oi_1 _3311_ (.Y(_1219_),
    .B1(net627),
    .B2(net127),
    .A2(net663),
    .A1(\bp_core.bp_stride_out[11] ));
 sg13g2_nand2_1 _3312_ (.Y(_0241_),
    .A(_1218_),
    .B(_1219_));
 sg13g2_nand2_1 _3313_ (.Y(_1220_),
    .A(net82),
    .B(net638));
 sg13g2_a22oi_1 _3314_ (.Y(_1221_),
    .B1(net629),
    .B2(\inter_bp.param_tx_shift_reg[34] ),
    .A2(net667),
    .A1(\bp_core.bp_stride_out[12] ));
 sg13g2_nand2_1 _3315_ (.Y(_0242_),
    .A(_1220_),
    .B(_1221_));
 sg13g2_nand2_1 _3316_ (.Y(_1222_),
    .A(net127),
    .B(net636));
 sg13g2_a22oi_1 _3317_ (.Y(_1223_),
    .B1(net627),
    .B2(\inter_bp.param_tx_shift_reg[35] ),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[13] ));
 sg13g2_nand2_1 _3318_ (.Y(_0243_),
    .A(_1222_),
    .B(_1223_));
 sg13g2_nand2_1 _3319_ (.Y(_1224_),
    .A(net111),
    .B(net636));
 sg13g2_a22oi_1 _3320_ (.Y(_1225_),
    .B1(net627),
    .B2(net92),
    .A2(net663),
    .A1(\bp_core.bp_stride_out[14] ));
 sg13g2_nand2_1 _3321_ (.Y(_0244_),
    .A(_1224_),
    .B(_1225_));
 sg13g2_nand2_1 _3322_ (.Y(_1226_),
    .A(net188),
    .B(net625));
 sg13g2_a22oi_1 _3323_ (.Y(_1227_),
    .B1(net635),
    .B2(\inter_bp.param_tx_shift_reg[35] ),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[15] ));
 sg13g2_nand2_1 _3324_ (.Y(_0245_),
    .A(_1226_),
    .B(_1227_));
 sg13g2_nand2_1 _3325_ (.Y(_1228_),
    .A(net92),
    .B(net637));
 sg13g2_a22oi_1 _3326_ (.Y(_1229_),
    .B1(net625),
    .B2(\inter_bp.param_tx_shift_reg[38] ),
    .A2(net662),
    .A1(\bp_core.bp_stride_out[16] ));
 sg13g2_nand2_1 _3327_ (.Y(_0246_),
    .A(_1228_),
    .B(_1229_));
 sg13g2_nand2_1 _3328_ (.Y(_1230_),
    .A(net175),
    .B(net625));
 sg13g2_a22oi_1 _3329_ (.Y(_1231_),
    .B1(net635),
    .B2(\inter_bp.param_tx_shift_reg[37] ),
    .A2(net664),
    .A1(\bp_core.bp_stride_out[17] ));
 sg13g2_nand2_1 _3330_ (.Y(_0247_),
    .A(_1230_),
    .B(_1231_));
 sg13g2_nand2_1 _3331_ (.Y(_1232_),
    .A(net96),
    .B(net635));
 sg13g2_a22oi_1 _3332_ (.Y(_1233_),
    .B1(net626),
    .B2(\inter_bp.param_tx_shift_reg[40] ),
    .A2(net664),
    .A1(\bp_core.bp_stride_out[18] ));
 sg13g2_nand2_1 _3333_ (.Y(_0248_),
    .A(_1232_),
    .B(_1233_));
 sg13g2_nand2_1 _3334_ (.Y(_1234_),
    .A(net390),
    .B(net628));
 sg13g2_a22oi_1 _3335_ (.Y(_1235_),
    .B1(net635),
    .B2(net175),
    .A2(net664),
    .A1(\bp_core.bp_stride_out[19] ));
 sg13g2_nand2_1 _3336_ (.Y(_0249_),
    .A(_1234_),
    .B(_1235_));
 sg13g2_nand2_1 _3337_ (.Y(_1236_),
    .A(net90),
    .B(net628));
 sg13g2_a22oi_1 _3338_ (.Y(_1237_),
    .B1(net637),
    .B2(net143),
    .A2(net666),
    .A1(\bp_core.bp_lambda_out[0] ));
 sg13g2_nand2_1 _3339_ (.Y(_0250_),
    .A(_1236_),
    .B(net144));
 sg13g2_nand2_1 _3340_ (.Y(_1238_),
    .A(net94),
    .B(net628));
 sg13g2_a22oi_1 _3341_ (.Y(_1239_),
    .B1(net640),
    .B2(\inter_bp.param_tx_shift_reg[41] ),
    .A2(net665),
    .A1(\bp_core.bp_lambda_out[1] ));
 sg13g2_nand2_1 _3342_ (.Y(_0251_),
    .A(_1238_),
    .B(_1239_));
 sg13g2_nand2_1 _3343_ (.Y(_1240_),
    .A(net90),
    .B(net637));
 sg13g2_a22oi_1 _3344_ (.Y(_1241_),
    .B1(net628),
    .B2(\inter_bp.param_tx_shift_reg[44] ),
    .A2(net666),
    .A1(\bp_core.bp_lambda_out[2] ));
 sg13g2_nand2_1 _3345_ (.Y(_0252_),
    .A(_1240_),
    .B(_1241_));
 sg13g2_nand2_1 _3346_ (.Y(_1242_),
    .A(net94),
    .B(net640));
 sg13g2_a22oi_1 _3347_ (.Y(_1243_),
    .B1(net629),
    .B2(net135),
    .A2(net665),
    .A1(\bp_core.bp_lambda_out[3] ));
 sg13g2_nand2_1 _3348_ (.Y(_0253_),
    .A(_1242_),
    .B(net136));
 sg13g2_nand2_1 _3349_ (.Y(_1244_),
    .A(net213),
    .B(net640));
 sg13g2_a22oi_1 _3350_ (.Y(_1245_),
    .B1(net628),
    .B2(\inter_bp.param_tx_shift_reg[46] ),
    .A2(net665),
    .A1(\bp_core.bp_lambda_out[4] ));
 sg13g2_nand2_1 _3351_ (.Y(_0254_),
    .A(_1244_),
    .B(_1245_));
 sg13g2_nand2_1 _3352_ (.Y(_1246_),
    .A(net135),
    .B(net640));
 sg13g2_a22oi_1 _3353_ (.Y(_1247_),
    .B1(net628),
    .B2(net196),
    .A2(net665),
    .A1(\bp_core.bp_lambda_out[5] ));
 sg13g2_nand2_1 _3354_ (.Y(_0255_),
    .A(_1246_),
    .B(net197));
 sg13g2_a22oi_1 _3355_ (.Y(_1248_),
    .B1(net640),
    .B2(net320),
    .A2(net665),
    .A1(\bp_core.bp_lambda_out[6] ));
 sg13g2_inv_1 _3356_ (.Y(_0256_),
    .A(net321));
 sg13g2_a22oi_1 _3357_ (.Y(_1249_),
    .B1(net640),
    .B2(net196),
    .A2(net665),
    .A1(net234));
 sg13g2_inv_1 _3358_ (.Y(_0257_),
    .A(_1249_));
 sg13g2_nor2_1 _3359_ (.A(\inter_bp.report_transmitting ),
    .B(net555),
    .Y(_1250_));
 sg13g2_and2_1 _3360_ (.A(\inter_bp.report_transmitting ),
    .B(net555),
    .X(_1251_));
 sg13g2_nor3_1 _3361_ (.A(net660),
    .B(net556),
    .C(_1251_),
    .Y(_0258_));
 sg13g2_a21oi_1 _3362_ (.A1(net1079),
    .A2(_1251_),
    .Y(_1252_),
    .B1(net660));
 sg13g2_o21ai_1 _3363_ (.B1(_1252_),
    .Y(_1253_),
    .A1(net1079),
    .A2(_1251_));
 sg13g2_inv_1 _3364_ (.Y(_0259_),
    .A(net1080));
 sg13g2_a21oi_1 _3365_ (.A1(\inter_bp.report_tx_counter[1] ),
    .A2(_1251_),
    .Y(_1254_),
    .B1(net325));
 sg13g2_and3_1 _3366_ (.X(_1255_),
    .A(\inter_bp.report_tx_counter[1] ),
    .B(net325),
    .C(_1251_));
 sg13g2_nor3_1 _3367_ (.A(net660),
    .B(net326),
    .C(_1255_),
    .Y(_0260_));
 sg13g2_nor2_1 _3368_ (.A(net1007),
    .B(_1255_),
    .Y(_1256_));
 sg13g2_and2_1 _3369_ (.A(net1007),
    .B(_1255_),
    .X(_1257_));
 sg13g2_nor3_1 _3370_ (.A(net660),
    .B(net1008),
    .C(_1257_),
    .Y(_0261_));
 sg13g2_a21oi_1 _3371_ (.A1(net1040),
    .A2(_1257_),
    .Y(_1258_),
    .B1(net660));
 sg13g2_o21ai_1 _3372_ (.B1(_1258_),
    .Y(_1259_),
    .A1(net1040),
    .A2(_1257_));
 sg13g2_inv_1 _3373_ (.Y(_0262_),
    .A(net1041));
 sg13g2_nor2b_2 _3374_ (.A(net660),
    .B_N(\inter_bp.report_transmitting ),
    .Y(_1260_));
 sg13g2_nand2_1 _3375_ (.Y(_1261_),
    .A(net182),
    .B(net634));
 sg13g2_a22oi_1 _3376_ (.Y(_1262_),
    .B1(net624),
    .B2(\inter_bp.report_tx_shift_reg[2] ),
    .A2(net661),
    .A1(\bp_core.bp_report_addr_out[0] ));
 sg13g2_nand2_1 _3377_ (.Y(_0263_),
    .A(net183),
    .B(_1262_));
 sg13g2_nand2_1 _3378_ (.Y(_1263_),
    .A(net247),
    .B(net661));
 sg13g2_a22oi_1 _3379_ (.Y(_1264_),
    .B1(net624),
    .B2(net185),
    .A2(net634),
    .A1(\inter_bp.report_tx_shift_reg[1] ));
 sg13g2_nand2_1 _3380_ (.Y(_0264_),
    .A(net248),
    .B(_1264_));
 sg13g2_nand2_1 _3381_ (.Y(_1265_),
    .A(net164),
    .B(net661));
 sg13g2_a22oi_1 _3382_ (.Y(_1266_),
    .B1(net624),
    .B2(\inter_bp.report_tx_shift_reg[4] ),
    .A2(net634),
    .A1(\inter_bp.report_tx_shift_reg[2] ));
 sg13g2_nand2_1 _3383_ (.Y(_0265_),
    .A(net165),
    .B(_1266_));
 sg13g2_nand2_1 _3384_ (.Y(_1267_),
    .A(net185),
    .B(net634));
 sg13g2_a22oi_1 _3385_ (.Y(_1268_),
    .B1(_1260_),
    .B2(net69),
    .A2(net661),
    .A1(\bp_core.bp_report_addr_out[3] ));
 sg13g2_nand2_1 _3386_ (.Y(_0266_),
    .A(net186),
    .B(_1268_));
 sg13g2_nand2_1 _3387_ (.Y(_1269_),
    .A(net115),
    .B(net661));
 sg13g2_a22oi_1 _3388_ (.Y(_1270_),
    .B1(_1260_),
    .B2(\inter_bp.report_tx_shift_reg[6] ),
    .A2(net634),
    .A1(\inter_bp.report_tx_shift_reg[4] ));
 sg13g2_nand2_1 _3389_ (.Y(_0267_),
    .A(net116),
    .B(_1270_));
 sg13g2_nand2_1 _3390_ (.Y(_1271_),
    .A(net69),
    .B(_1048_));
 sg13g2_a22oi_1 _3391_ (.Y(_1272_),
    .B1(net624),
    .B2(\inter_bp.report_tx_shift_reg[7] ),
    .A2(net659),
    .A1(\bp_core.bp_report_addr_out[5] ));
 sg13g2_nand2_1 _3392_ (.Y(_0268_),
    .A(net70),
    .B(_1272_));
 sg13g2_nand2_1 _3393_ (.Y(_1273_),
    .A(net208),
    .B(net661));
 sg13g2_a22oi_1 _3394_ (.Y(_1274_),
    .B1(_1260_),
    .B2(\inter_bp.report_tx_shift_reg[8] ),
    .A2(net634),
    .A1(\inter_bp.report_tx_shift_reg[6] ));
 sg13g2_nand2_1 _3395_ (.Y(_0269_),
    .A(net209),
    .B(_1274_));
 sg13g2_nand2_1 _3396_ (.Y(_1275_),
    .A(net124),
    .B(net659));
 sg13g2_a22oi_1 _3397_ (.Y(_1276_),
    .B1(net623),
    .B2(\inter_bp.report_tx_shift_reg[9] ),
    .A2(net633),
    .A1(\inter_bp.report_tx_shift_reg[7] ));
 sg13g2_nand2_1 _3398_ (.Y(_0270_),
    .A(net125),
    .B(_1276_));
 sg13g2_nand2_1 _3399_ (.Y(_1277_),
    .A(net74),
    .B(net659));
 sg13g2_a22oi_1 _3400_ (.Y(_1278_),
    .B1(net624),
    .B2(\inter_bp.report_tx_shift_reg[10] ),
    .A2(net633),
    .A1(\inter_bp.report_tx_shift_reg[8] ));
 sg13g2_nand2_1 _3401_ (.Y(_0271_),
    .A(net75),
    .B(_1278_));
 sg13g2_nand2_1 _3402_ (.Y(_1279_),
    .A(net145),
    .B(net658));
 sg13g2_a22oi_1 _3403_ (.Y(_1280_),
    .B1(net624),
    .B2(net118),
    .A2(net633),
    .A1(\inter_bp.report_tx_shift_reg[9] ));
 sg13g2_nand2_1 _3404_ (.Y(_0272_),
    .A(net146),
    .B(_1280_));
 sg13g2_nand2_1 _3405_ (.Y(_1281_),
    .A(net64),
    .B(net659));
 sg13g2_a22oi_1 _3406_ (.Y(_1282_),
    .B1(net624),
    .B2(\inter_bp.report_tx_shift_reg[12] ),
    .A2(net633),
    .A1(\inter_bp.report_tx_shift_reg[10] ));
 sg13g2_nand2_1 _3407_ (.Y(_0273_),
    .A(net65),
    .B(_1282_));
 sg13g2_nand2_1 _3408_ (.Y(_1283_),
    .A(net118),
    .B(net632));
 sg13g2_a22oi_1 _3409_ (.Y(_1284_),
    .B1(net623),
    .B2(net109),
    .A2(net658),
    .A1(\bp_core.bp_report_addr_out[11] ));
 sg13g2_nand2_1 _3410_ (.Y(_0274_),
    .A(_1283_),
    .B(_1284_));
 sg13g2_nand2_1 _3411_ (.Y(_1285_),
    .A(net203),
    .B(net658));
 sg13g2_a22oi_1 _3412_ (.Y(_1286_),
    .B1(net623),
    .B2(\inter_bp.report_tx_shift_reg[14] ),
    .A2(net632),
    .A1(\inter_bp.report_tx_shift_reg[12] ));
 sg13g2_nand2_1 _3413_ (.Y(_0275_),
    .A(net204),
    .B(_1286_));
 sg13g2_nand2_1 _3414_ (.Y(_1287_),
    .A(net109),
    .B(net632));
 sg13g2_a22oi_1 _3415_ (.Y(_1288_),
    .B1(net623),
    .B2(\inter_bp.report_tx_shift_reg[15] ),
    .A2(net658),
    .A1(\bp_core.bp_report_addr_out[13] ));
 sg13g2_nand2_1 _3416_ (.Y(_0276_),
    .A(_1287_),
    .B(_1288_));
 sg13g2_nand2_1 _3417_ (.Y(_1289_),
    .A(net275),
    .B(net658));
 sg13g2_a22oi_1 _3418_ (.Y(_1290_),
    .B1(net623),
    .B2(net133),
    .A2(net632),
    .A1(\inter_bp.report_tx_shift_reg[14] ));
 sg13g2_nand2_1 _3419_ (.Y(_0277_),
    .A(net276),
    .B(_1290_));
 sg13g2_nand2_1 _3420_ (.Y(_1291_),
    .A(net150),
    .B(net632));
 sg13g2_a22oi_1 _3421_ (.Y(_1292_),
    .B1(net623),
    .B2(\inter_bp.report_tx_shift_reg[17] ),
    .A2(net658),
    .A1(\bp_core.bp_report_addr_out[15] ));
 sg13g2_nand2_1 _3422_ (.Y(_0278_),
    .A(_1291_),
    .B(_1292_));
 sg13g2_nand2_1 _3423_ (.Y(_1293_),
    .A(net133),
    .B(net632));
 sg13g2_a22oi_1 _3424_ (.Y(_1294_),
    .B1(net623),
    .B2(\inter_bp.report_tx_shift_reg[18] ),
    .A2(net658),
    .A1(\bp_core.bp_report_addr_out[16] ));
 sg13g2_nand2_1 _3425_ (.Y(_0279_),
    .A(_1293_),
    .B(_1294_));
 sg13g2_nand2_1 _3426_ (.Y(_1295_),
    .A(net156),
    .B(net658));
 sg13g2_a22oi_1 _3427_ (.Y(_1296_),
    .B1(net623),
    .B2(\inter_bp.report_tx_shift_reg[19] ),
    .A2(net632),
    .A1(\inter_bp.report_tx_shift_reg[17] ));
 sg13g2_nand2_1 _3428_ (.Y(_0280_),
    .A(net157),
    .B(_1296_));
 sg13g2_a22oi_1 _3429_ (.Y(_1297_),
    .B1(net632),
    .B2(net284),
    .A2(net659),
    .A1(\bp_core.bp_report_addr_out[18] ));
 sg13g2_inv_1 _3430_ (.Y(_0281_),
    .A(net285));
 sg13g2_a22oi_1 _3431_ (.Y(_1298_),
    .B1(net633),
    .B2(net259),
    .A2(net659),
    .A1(\bp_core.bp_report_addr_out[19] ));
 sg13g2_inv_1 _3432_ (.Y(_0282_),
    .A(net260));
 sg13g2_nor3_1 _3433_ (.A(\bp_core.params_module.state[3] ),
    .B(net731),
    .C(\bp_core.params_module.state[1] ),
    .Y(_1299_));
 sg13g2_o21ai_1 _3434_ (.B1(_0835_),
    .Y(_1300_),
    .A1(\bp_core.params_module.state[0] ),
    .A2(_1299_));
 sg13g2_nand3_1 _3435_ (.B(_0834_),
    .C(_1300_),
    .A(_0831_),
    .Y(_1301_));
 sg13g2_nor2_1 _3436_ (.A(_0524_),
    .B(_1301_),
    .Y(_1302_));
 sg13g2_o21ai_1 _3437_ (.B1(_0719_),
    .Y(_1303_),
    .A1(net59),
    .A2(net734));
 sg13g2_nor2_1 _3438_ (.A(_1301_),
    .B(_1303_),
    .Y(_1304_));
 sg13g2_nor2_1 _3439_ (.A(net1149),
    .B(_1304_),
    .Y(_1305_));
 sg13g2_nor2_1 _3440_ (.A(_1302_),
    .B(_1305_),
    .Y(_0283_));
 sg13g2_nor2_1 _3441_ (.A(net738),
    .B(_1302_),
    .Y(_1306_));
 sg13g2_nand2b_1 _3442_ (.Y(_1307_),
    .B(_1303_),
    .A_N(_1301_));
 sg13g2_inv_1 _3443_ (.Y(_1308_),
    .A(_1307_));
 sg13g2_nand2_1 _3444_ (.Y(_1309_),
    .A(net738),
    .B(net1155));
 sg13g2_nand2_1 _3445_ (.Y(_1310_),
    .A(net738),
    .B(_1302_));
 sg13g2_inv_1 _3446_ (.Y(_1311_),
    .A(_1310_));
 sg13g2_nor3_1 _3447_ (.A(_1306_),
    .B(_1308_),
    .C(_1311_),
    .Y(_0284_));
 sg13g2_nor2_1 _3448_ (.A(net1147),
    .B(_1311_),
    .Y(_1312_));
 sg13g2_a21oi_1 _3449_ (.A1(net1147),
    .A2(_1311_),
    .Y(_1313_),
    .B1(_1308_));
 sg13g2_nor2b_1 _3450_ (.A(net1148),
    .B_N(_1313_),
    .Y(_0285_));
 sg13g2_nand2b_2 _3451_ (.Y(_1314_),
    .B(net1147),
    .A_N(\bp_core.params_module.counter[3] ));
 sg13g2_nor2_2 _3452_ (.A(_1309_),
    .B(_1314_),
    .Y(_1315_));
 sg13g2_a22oi_1 _3453_ (.Y(_1316_),
    .B1(_1315_),
    .B2(_1304_),
    .A2(_1313_),
    .A1(net1097));
 sg13g2_inv_1 _3454_ (.Y(_0286_),
    .A(_1316_));
 sg13g2_nand3_1 _3455_ (.B(net996),
    .C(net230),
    .A(net10),
    .Y(_1317_));
 sg13g2_a22oi_1 _3456_ (.Y(_0287_),
    .B1(_0946_),
    .B2(_1317_),
    .A2(_0558_),
    .A1(net890));
 sg13g2_mux2_1 _3457_ (.A0(net1000),
    .A1(net4),
    .S(_0826_),
    .X(_0288_));
 sg13g2_nor2_1 _3458_ (.A(net423),
    .B(_0826_),
    .Y(_1318_));
 sg13g2_a21oi_1 _3459_ (.A1(net5),
    .A2(_0826_),
    .Y(_0289_),
    .B1(net424));
 sg13g2_nor2_1 _3460_ (.A(net420),
    .B(_0826_),
    .Y(_1319_));
 sg13g2_a21oi_1 _3461_ (.A1(net6),
    .A2(_0826_),
    .Y(_0290_),
    .B1(net421));
 sg13g2_a21oi_1 _3462_ (.A1(_0526_),
    .A2(_0098_),
    .Y(_1320_),
    .B1(_0715_));
 sg13g2_nand2_2 _3463_ (.Y(_1321_),
    .A(_0836_),
    .B(_1320_));
 sg13g2_inv_2 _3464_ (.Y(_1322_),
    .A(_1321_));
 sg13g2_nor3_2 _3465_ (.A(net738),
    .B(_0524_),
    .C(_1314_),
    .Y(_1323_));
 sg13g2_o21ai_1 _3466_ (.B1(_1322_),
    .Y(_1324_),
    .A1(_0721_),
    .A2(_1323_));
 sg13g2_nand2_2 _3467_ (.Y(_1325_),
    .A(net731),
    .B(net4));
 sg13g2_o21ai_1 _3468_ (.B1(net657),
    .Y(_1326_),
    .A1(net729),
    .A2(_0610_));
 sg13g2_mux2_1 _3469_ (.A0(_1326_),
    .A1(net1154),
    .S(_1324_),
    .X(_0291_));
 sg13g2_nand2_2 _3470_ (.Y(_1327_),
    .A(net5),
    .B(net732));
 sg13g2_o21ai_1 _3471_ (.B1(_1327_),
    .Y(_1328_),
    .A1(net736),
    .A2(_0612_));
 sg13g2_mux2_1 _3472_ (.A0(_1328_),
    .A1(net1175),
    .S(_1324_),
    .X(_0292_));
 sg13g2_nand2_2 _3473_ (.Y(_1329_),
    .A(net6),
    .B(net732));
 sg13g2_o21ai_1 _3474_ (.B1(net655),
    .Y(_1330_),
    .A1(net729),
    .A2(_0614_));
 sg13g2_mux2_1 _3475_ (.A0(_1330_),
    .A1(net1164),
    .S(_1324_),
    .X(_0293_));
 sg13g2_nand2_2 _3476_ (.Y(_1331_),
    .A(net7),
    .B(net731));
 sg13g2_o21ai_1 _3477_ (.B1(_1331_),
    .Y(_1332_),
    .A1(net736),
    .A2(_0616_));
 sg13g2_mux2_1 _3478_ (.A0(_1332_),
    .A1(net1171),
    .S(_1324_),
    .X(_0294_));
 sg13g2_nand2_2 _3479_ (.Y(_1333_),
    .A(net732),
    .B(net8));
 sg13g2_o21ai_1 _3480_ (.B1(net653),
    .Y(_1334_),
    .A1(net729),
    .A2(_0618_));
 sg13g2_mux2_1 _3481_ (.A0(_1334_),
    .A1(net202),
    .S(_1324_),
    .X(_0295_));
 sg13g2_o21ai_1 _3482_ (.B1(_1322_),
    .Y(_1335_),
    .A1(_0718_),
    .A2(_0721_));
 sg13g2_o21ai_1 _3483_ (.B1(net657),
    .Y(_1336_),
    .A1(net731),
    .A2(_0638_));
 sg13g2_mux2_1 _3484_ (.A0(_1336_),
    .A1(net1160),
    .S(_1335_),
    .X(_0296_));
 sg13g2_a21oi_1 _3485_ (.A1(_0526_),
    .A2(net1123),
    .Y(_1337_),
    .B1(_1335_));
 sg13g2_a22oi_1 _3486_ (.Y(_0297_),
    .B1(_1337_),
    .B2(net656),
    .A2(_1335_),
    .A1(_0652_));
 sg13g2_o21ai_1 _3487_ (.B1(net655),
    .Y(_1338_),
    .A1(net731),
    .A2(_0640_));
 sg13g2_mux2_1 _3488_ (.A0(_1338_),
    .A1(net1172),
    .S(_1335_),
    .X(_0298_));
 sg13g2_o21ai_1 _3489_ (.B1(net654),
    .Y(_1339_),
    .A1(net731),
    .A2(_0642_));
 sg13g2_mux2_1 _3490_ (.A0(_1339_),
    .A1(net1177),
    .S(_1335_),
    .X(_0299_));
 sg13g2_o21ai_1 _3491_ (.B1(net653),
    .Y(_1340_),
    .A1(net731),
    .A2(_0644_));
 sg13g2_mux2_1 _3492_ (.A0(_1340_),
    .A1(net1168),
    .S(_1335_),
    .X(_0300_));
 sg13g2_nand2_1 _3493_ (.Y(_1341_),
    .A(\bp_core.params_module.counter[1] ),
    .B(_0524_));
 sg13g2_nor2_2 _3494_ (.A(_1314_),
    .B(_1341_),
    .Y(_1342_));
 sg13g2_o21ai_1 _3495_ (.B1(_1322_),
    .Y(_1343_),
    .A1(_0526_),
    .A2(_1342_));
 sg13g2_o21ai_1 _3496_ (.B1(net657),
    .Y(_1344_),
    .A1(net729),
    .A2(_0620_));
 sg13g2_mux2_1 _3497_ (.A0(_1344_),
    .A1(net1128),
    .S(_1343_),
    .X(_0301_));
 sg13g2_nand2_1 _3498_ (.Y(_1345_),
    .A(_0526_),
    .B(net512));
 sg13g2_nor2b_1 _3499_ (.A(_1343_),
    .B_N(net656),
    .Y(_1346_));
 sg13g2_a22oi_1 _3500_ (.Y(_0302_),
    .B1(_1345_),
    .B2(_1346_),
    .A2(_1343_),
    .A1(_0539_));
 sg13g2_o21ai_1 _3501_ (.B1(net655),
    .Y(_1347_),
    .A1(net729),
    .A2(_0622_));
 sg13g2_mux2_1 _3502_ (.A0(_1347_),
    .A1(net1162),
    .S(_1343_),
    .X(_0303_));
 sg13g2_o21ai_1 _3503_ (.B1(net654),
    .Y(_1348_),
    .A1(net728),
    .A2(_0624_));
 sg13g2_mux2_1 _3504_ (.A0(_1348_),
    .A1(net1167),
    .S(_1343_),
    .X(_0304_));
 sg13g2_o21ai_1 _3505_ (.B1(net653),
    .Y(_1349_),
    .A1(net728),
    .A2(_0626_));
 sg13g2_mux2_1 _3506_ (.A0(_1349_),
    .A1(net1144),
    .S(_1343_),
    .X(_0305_));
 sg13g2_nor2_2 _3507_ (.A(_0722_),
    .B(_1321_),
    .Y(_1350_));
 sg13g2_o21ai_1 _3508_ (.B1(net657),
    .Y(_1351_),
    .A1(net733),
    .A2(_0646_));
 sg13g2_mux2_1 _3509_ (.A0(net1158),
    .A1(_1351_),
    .S(_1350_),
    .X(_0306_));
 sg13g2_o21ai_1 _3510_ (.B1(net656),
    .Y(_1352_),
    .A1(net734),
    .A2(_0648_));
 sg13g2_mux2_1 _3511_ (.A0(net399),
    .A1(_1352_),
    .S(_1350_),
    .X(_0307_));
 sg13g2_o21ai_1 _3512_ (.B1(net655),
    .Y(_1353_),
    .A1(net732),
    .A2(_0650_));
 sg13g2_mux2_1 _3513_ (.A0(net234),
    .A1(_1353_),
    .S(_1350_),
    .X(_0308_));
 sg13g2_nand3_1 _3514_ (.B(_0822_),
    .C(_1052_),
    .A(_0820_),
    .Y(_1354_));
 sg13g2_o21ai_1 _3515_ (.B1(net722),
    .Y(_1355_),
    .A1(\bp_core.addr_reg[0] ),
    .A2(\bp_core.bp_stride_out[0] ));
 sg13g2_nand2b_1 _3516_ (.Y(_1356_),
    .B(_0730_),
    .A_N(_1355_));
 sg13g2_o21ai_1 _3517_ (.B1(_1356_),
    .Y(_1357_),
    .A1(_0527_),
    .A2(net722));
 sg13g2_mux2_1 _3518_ (.A0(_1357_),
    .A1(net1059),
    .S(net568),
    .X(_0309_));
 sg13g2_a21oi_1 _3519_ (.A1(_0730_),
    .A2(_0731_),
    .Y(_1358_),
    .B1(net720));
 sg13g2_o21ai_1 _3520_ (.B1(_1358_),
    .Y(_1359_),
    .A1(_0730_),
    .A2(_0731_));
 sg13g2_o21ai_1 _3521_ (.B1(_1359_),
    .Y(_1360_),
    .A1(_0528_),
    .A2(net726));
 sg13g2_mux2_1 _3522_ (.A0(_1360_),
    .A1(net1032),
    .S(net568),
    .X(_0310_));
 sg13g2_nand2b_1 _3523_ (.Y(_1361_),
    .B(net1142),
    .A_N(_0732_));
 sg13g2_nand2b_1 _3524_ (.Y(_1362_),
    .B(_0732_),
    .A_N(_0737_));
 sg13g2_nand3_1 _3525_ (.B(_1361_),
    .C(_1362_),
    .A(net726),
    .Y(_1363_));
 sg13g2_o21ai_1 _3526_ (.B1(_1363_),
    .Y(_1364_),
    .A1(_0529_),
    .A2(net726));
 sg13g2_mux2_1 _3527_ (.A0(_1364_),
    .A1(net1023),
    .S(net566),
    .X(_0311_));
 sg13g2_nand3_1 _3528_ (.B(_0736_),
    .C(_1362_),
    .A(_0735_),
    .Y(_1365_));
 sg13g2_a21o_1 _3529_ (.A2(_1362_),
    .A1(_0736_),
    .B1(_0735_),
    .X(_1366_));
 sg13g2_nand3_1 _3530_ (.B(_1365_),
    .C(_1366_),
    .A(net726),
    .Y(_1367_));
 sg13g2_o21ai_1 _3531_ (.B1(_1367_),
    .Y(_1368_),
    .A1(_0530_),
    .A2(net726));
 sg13g2_mux2_1 _3532_ (.A0(_1368_),
    .A1(net1102),
    .S(net566),
    .X(_0312_));
 sg13g2_nand2b_1 _3533_ (.Y(_1369_),
    .B(_0749_),
    .A_N(_0740_));
 sg13g2_nand2b_2 _3534_ (.Y(_1370_),
    .B(_0740_),
    .A_N(_0749_));
 sg13g2_nand3_1 _3535_ (.B(_1369_),
    .C(_1370_),
    .A(net726),
    .Y(_1371_));
 sg13g2_o21ai_1 _3536_ (.B1(_1371_),
    .Y(_1372_),
    .A1(_0531_),
    .A2(net726));
 sg13g2_mux2_1 _3537_ (.A0(_1372_),
    .A1(net1056),
    .S(net566),
    .X(_0313_));
 sg13g2_nand3_1 _3538_ (.B(_0748_),
    .C(_1370_),
    .A(_0747_),
    .Y(_1373_));
 sg13g2_a21o_1 _3539_ (.A2(_1370_),
    .A1(_0748_),
    .B1(_0747_),
    .X(_1374_));
 sg13g2_nand3_1 _3540_ (.B(_1373_),
    .C(_1374_),
    .A(net726),
    .Y(_1375_));
 sg13g2_o21ai_1 _3541_ (.B1(_1375_),
    .Y(_1376_),
    .A1(_0532_),
    .A2(net727));
 sg13g2_mux2_1 _3542_ (.A0(_1376_),
    .A1(net1095),
    .S(net566),
    .X(_0314_));
 sg13g2_a21oi_1 _3543_ (.A1(_0751_),
    .A2(_1370_),
    .Y(_1377_),
    .B1(_0746_));
 sg13g2_or2_1 _3544_ (.X(_1378_),
    .B(_1377_),
    .A(_0744_));
 sg13g2_nand2_1 _3545_ (.Y(_1379_),
    .A(_0744_),
    .B(_1377_));
 sg13g2_nand3_1 _3546_ (.B(_1378_),
    .C(_1379_),
    .A(net724),
    .Y(_1380_));
 sg13g2_o21ai_1 _3547_ (.B1(_1380_),
    .Y(_1381_),
    .A1(_0533_),
    .A2(net723));
 sg13g2_mux2_1 _3548_ (.A0(_1381_),
    .A1(net1112),
    .S(net566),
    .X(_0315_));
 sg13g2_nand3_1 _3549_ (.B(_0743_),
    .C(_1379_),
    .A(_0742_),
    .Y(_1382_));
 sg13g2_a21o_1 _3550_ (.A2(_1379_),
    .A1(_0743_),
    .B1(_0742_),
    .X(_1383_));
 sg13g2_nand3_1 _3551_ (.B(_1382_),
    .C(_1383_),
    .A(net724),
    .Y(_1384_));
 sg13g2_o21ai_1 _3552_ (.B1(_1384_),
    .Y(_1385_),
    .A1(_0534_),
    .A2(net724));
 sg13g2_mux2_1 _3553_ (.A0(_1385_),
    .A1(net1089),
    .S(net567),
    .X(_0316_));
 sg13g2_a21oi_1 _3554_ (.A1(_0757_),
    .A2(_0778_),
    .Y(_1386_),
    .B1(net718));
 sg13g2_o21ai_1 _3555_ (.B1(_1386_),
    .Y(_1387_),
    .A1(_0757_),
    .A2(_0778_));
 sg13g2_o21ai_1 _3556_ (.B1(_1387_),
    .Y(_1388_),
    .A1(_0535_),
    .A2(net723));
 sg13g2_mux2_1 _3557_ (.A0(_1388_),
    .A1(net1073),
    .S(net567),
    .X(_0317_));
 sg13g2_a21oi_1 _3558_ (.A1(_0757_),
    .A2(_0778_),
    .Y(_1389_),
    .B1(_0776_));
 sg13g2_nand2b_1 _3559_ (.Y(_1390_),
    .B(_0781_),
    .A_N(_1389_));
 sg13g2_nand2b_1 _3560_ (.Y(_1391_),
    .B(_1389_),
    .A_N(_0781_));
 sg13g2_nand3_1 _3561_ (.B(_1390_),
    .C(_1391_),
    .A(net724),
    .Y(_1392_));
 sg13g2_o21ai_1 _3562_ (.B1(_1392_),
    .Y(_1393_),
    .A1(_0536_),
    .A2(net724));
 sg13g2_mux2_1 _3563_ (.A0(_1393_),
    .A1(net1091),
    .S(net566),
    .X(_0318_));
 sg13g2_and2_1 _3564_ (.A(_0779_),
    .B(_1389_),
    .X(_1394_));
 sg13g2_o21ai_1 _3565_ (.B1(_0774_),
    .Y(_1395_),
    .A1(_0780_),
    .A2(_1394_));
 sg13g2_or3_1 _3566_ (.A(_0774_),
    .B(_0780_),
    .C(_1394_),
    .X(_1396_));
 sg13g2_nand3_1 _3567_ (.B(_1395_),
    .C(_1396_),
    .A(net723),
    .Y(_1397_));
 sg13g2_o21ai_1 _3568_ (.B1(_1397_),
    .Y(_1398_),
    .A1(_0537_),
    .A2(net723));
 sg13g2_mux2_1 _3569_ (.A0(_1398_),
    .A1(net1072),
    .S(net567),
    .X(_0319_));
 sg13g2_nand3_1 _3570_ (.B(_0773_),
    .C(_1396_),
    .A(_0772_),
    .Y(_1399_));
 sg13g2_a21o_1 _3571_ (.A2(_1396_),
    .A1(_0773_),
    .B1(_0772_),
    .X(_1400_));
 sg13g2_nand3_1 _3572_ (.B(_1399_),
    .C(_1400_),
    .A(net723),
    .Y(_1401_));
 sg13g2_o21ai_1 _3573_ (.B1(_1401_),
    .Y(_1402_),
    .A1(_0538_),
    .A2(net723));
 sg13g2_mux2_1 _3574_ (.A0(_1402_),
    .A1(net1081),
    .S(net567),
    .X(_0320_));
 sg13g2_o21ai_1 _3575_ (.B1(_0786_),
    .Y(_1403_),
    .A1(_0756_),
    .A2(_0782_));
 sg13g2_a21oi_1 _3576_ (.A1(_0770_),
    .A2(_1403_),
    .Y(_1404_),
    .B1(net719));
 sg13g2_dfrbpq_1 _3577_ (.RESET_B(net777),
    .D(net398),
    .Q(\bp_addr_in[0] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _3578_ (.RESET_B(net824),
    .D(_0055_),
    .Q(\bp_addr_in[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _3579_ (.RESET_B(net811),
    .D(_0056_),
    .Q(\bp_addr_in[2] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _3580_ (.RESET_B(net825),
    .D(_0057_),
    .Q(\bp_addr_in[3] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _3581_ (.RESET_B(net811),
    .D(_0058_),
    .Q(\bp_addr_in[4] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _3582_ (.RESET_B(net820),
    .D(_0059_),
    .Q(\bp_addr_in[5] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3583_ (.RESET_B(net819),
    .D(_0060_),
    .Q(\bp_addr_in[6] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _3584_ (.RESET_B(net820),
    .D(_0061_),
    .Q(\bp_addr_in[7] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3585_ (.RESET_B(net819),
    .D(_0062_),
    .Q(\bp_addr_in[8] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _3586_ (.RESET_B(net818),
    .D(_0063_),
    .Q(\bp_addr_in[9] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _3587_ (.RESET_B(net818),
    .D(_0045_),
    .Q(\bp_addr_in[10] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _3588_ (.RESET_B(net818),
    .D(_0046_),
    .Q(\bp_addr_in[11] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _3589_ (.RESET_B(net818),
    .D(_0047_),
    .Q(\bp_addr_in[12] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _3590_ (.RESET_B(net810),
    .D(_0048_),
    .Q(\bp_addr_in[13] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _3591_ (.RESET_B(net810),
    .D(_0049_),
    .Q(\bp_addr_in[14] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _3592_ (.RESET_B(net773),
    .D(_0050_),
    .Q(\bp_addr_in[15] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _3593_ (.RESET_B(net770),
    .D(net941),
    .Q(\bp_addr_in[16] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _3594_ (.RESET_B(net769),
    .D(_0052_),
    .Q(\bp_addr_in[17] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _3595_ (.RESET_B(net770),
    .D(_0053_),
    .Q(\bp_addr_in[18] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _3596_ (.RESET_B(net769),
    .D(_0054_),
    .Q(\bp_addr_in[19] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _3597_ (.RESET_B(net775),
    .D(_0072_),
    .Q(\bp_core.bp_param_valid_in ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _3598_ (.RESET_B(net774),
    .D(_0106_),
    .Q(\inter_bp.param_shift_reg[0] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _3599_ (.RESET_B(net820),
    .D(_0107_),
    .Q(\inter_bp.param_shift_reg[1] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _3600_ (.RESET_B(net811),
    .D(_0108_),
    .Q(\inter_bp.param_shift_reg[2] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _3601_ (.RESET_B(net820),
    .D(_0109_),
    .Q(\inter_bp.param_shift_reg[3] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _3602_ (.RESET_B(net812),
    .D(_0110_),
    .Q(\inter_bp.param_shift_reg[4] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _3603_ (.RESET_B(net818),
    .D(_0111_),
    .Q(\inter_bp.param_shift_reg[5] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _3604_ (.RESET_B(net811),
    .D(_0112_),
    .Q(\inter_bp.param_shift_reg[6] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _3605_ (.RESET_B(net818),
    .D(_0113_),
    .Q(\inter_bp.param_shift_reg[7] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _3606_ (.RESET_B(net810),
    .D(_0114_),
    .Q(\inter_bp.param_shift_reg[8] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _3607_ (.RESET_B(net819),
    .D(_0115_),
    .Q(\inter_bp.param_shift_reg[9] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _3608_ (.RESET_B(net812),
    .D(_0116_),
    .Q(\inter_bp.param_shift_reg[10] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _3609_ (.RESET_B(net810),
    .D(_0117_),
    .Q(\inter_bp.param_shift_reg[11] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _3610_ (.RESET_B(net810),
    .D(_0118_),
    .Q(\inter_bp.param_shift_reg[12] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _3611_ (.RESET_B(net810),
    .D(_0119_),
    .Q(\inter_bp.param_shift_reg[13] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _3612_ (.RESET_B(net773),
    .D(_0120_),
    .Q(\inter_bp.param_shift_reg[14] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _3613_ (.RESET_B(net770),
    .D(_0121_),
    .Q(\inter_bp.param_shift_reg[15] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _3614_ (.RESET_B(net769),
    .D(_0122_),
    .Q(\inter_bp.param_shift_reg[16] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _3615_ (.RESET_B(net769),
    .D(_0123_),
    .Q(\inter_bp.param_shift_reg[17] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _3616_ (.RESET_B(net770),
    .D(_0124_),
    .Q(\inter_bp.param_shift_reg[18] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _3617_ (.RESET_B(net760),
    .D(_0125_),
    .Q(\inter_bp.param_shift_reg[19] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _3618_ (.RESET_B(net773),
    .D(_0126_),
    .Q(\inter_bp.param_shift_reg[20] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _3619_ (.RESET_B(net760),
    .D(_0127_),
    .Q(\inter_bp.param_shift_reg[21] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _3620_ (.RESET_B(net807),
    .D(_0128_),
    .Q(\inter_bp.param_shift_reg[22] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _3621_ (.RESET_B(net760),
    .D(_0129_),
    .Q(\inter_bp.param_shift_reg[23] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _3622_ (.RESET_B(net807),
    .D(_0130_),
    .Q(\inter_bp.param_shift_reg[24] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _3623_ (.RESET_B(net759),
    .D(_0131_),
    .Q(\inter_bp.param_shift_reg[25] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _3624_ (.RESET_B(net807),
    .D(_0132_),
    .Q(\inter_bp.param_shift_reg[26] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _3625_ (.RESET_B(net759),
    .D(_0133_),
    .Q(\inter_bp.param_shift_reg[27] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _3626_ (.RESET_B(net773),
    .D(_0134_),
    .Q(\inter_bp.param_shift_reg[28] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _3627_ (.RESET_B(net758),
    .D(_0135_),
    .Q(\inter_bp.param_shift_reg[29] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _3628_ (.RESET_B(net773),
    .D(_0136_),
    .Q(\inter_bp.param_shift_reg[30] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _3629_ (.RESET_B(net757),
    .D(_0137_),
    .Q(\inter_bp.param_shift_reg[31] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _3630_ (.RESET_B(net769),
    .D(_0138_),
    .Q(\inter_bp.param_shift_reg[32] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _3631_ (.RESET_B(net758),
    .D(_0139_),
    .Q(\inter_bp.param_shift_reg[33] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _3632_ (.RESET_B(net771),
    .D(_0140_),
    .Q(\inter_bp.param_shift_reg[34] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _3633_ (.RESET_B(net758),
    .D(_0141_),
    .Q(\inter_bp.param_shift_reg[35] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _3634_ (.RESET_B(net771),
    .D(_0142_),
    .Q(\inter_bp.param_shift_reg[36] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _3635_ (.RESET_B(net758),
    .D(_0143_),
    .Q(\inter_bp.param_shift_reg[37] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _3636_ (.RESET_B(net761),
    .D(_0144_),
    .Q(\inter_bp.param_shift_reg[38] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _3637_ (.RESET_B(net762),
    .D(_0145_),
    .Q(\inter_bp.param_shift_reg[39] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _3638_ (.RESET_B(net766),
    .D(_0146_),
    .Q(\inter_bp.param_shift_reg[40] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _3639_ (.RESET_B(net765),
    .D(_0147_),
    .Q(\inter_bp.param_shift_reg[41] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _3640_ (.RESET_B(net766),
    .D(_0148_),
    .Q(\inter_bp.param_shift_reg[42] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _3641_ (.RESET_B(net762),
    .D(_0149_),
    .Q(\inter_bp.param_shift_reg[43] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _3642_ (.RESET_B(net764),
    .D(_0150_),
    .Q(\inter_bp.param_shift_reg[44] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _3643_ (.RESET_B(net763),
    .D(_0151_),
    .Q(\inter_bp.param_shift_reg[45] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _3644_ (.RESET_B(net763),
    .D(_0152_),
    .Q(\inter_bp.param_shift_reg[46] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _3645_ (.RESET_B(net763),
    .D(_0153_),
    .Q(\inter_bp.param_shift_reg[47] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _3646_ (.RESET_B(net791),
    .D(_0096_),
    .Q(\inter_bp.report_rx_done ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _3647_ (.RESET_B(net790),
    .D(net309),
    .Q(\inter_bp.report_rx_counter[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _3648_ (.RESET_B(net790),
    .D(_0155_),
    .Q(\inter_bp.report_rx_counter[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _3649_ (.RESET_B(net790),
    .D(_0156_),
    .Q(\inter_bp.report_rx_counter[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _3650_ (.RESET_B(net790),
    .D(net450),
    .Q(\inter_bp.report_rx_counter[3] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _3651_ (.RESET_B(net790),
    .D(net324),
    .Q(\inter_bp.report_rx_counter[4] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _3652_ (.RESET_B(net775),
    .D(net946),
    .Q(\bp_core.bp_lambda_in[0] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _3653_ (.RESET_B(net766),
    .D(net350),
    .Q(\bp_core.bp_lambda_in[1] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _3654_ (.RESET_B(net767),
    .D(_0066_),
    .Q(\bp_core.bp_lambda_in[2] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _3655_ (.RESET_B(net762),
    .D(net863),
    .Q(\bp_core.bp_lambda_in[3] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _3656_ (.RESET_B(net766),
    .D(_0068_),
    .Q(\bp_core.bp_lambda_in[4] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _3657_ (.RESET_B(net767),
    .D(net887),
    .Q(\bp_core.bp_lambda_in[5] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _3658_ (.RESET_B(net767),
    .D(net993),
    .Q(\bp_core.bp_lambda_in[6] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _3659_ (.RESET_B(net767),
    .D(_0071_),
    .Q(\bp_core.bp_lambda_in[7] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _3660_ (.RESET_B(net791),
    .D(net11),
    .Q(\inter_bp.from_left_report_valid_prev ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3661_ (.RESET_B(net762),
    .D(net10),
    .Q(\inter_bp.from_left_param_valid_prev ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _3662_ (.RESET_B(net790),
    .D(_0159_),
    .Q(\inter_bp.report_shift_reg[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _3663_ (.RESET_B(net788),
    .D(_0160_),
    .Q(\inter_bp.report_shift_reg[1] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _3664_ (.RESET_B(net790),
    .D(_0161_),
    .Q(\inter_bp.report_shift_reg[2] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _3665_ (.RESET_B(net788),
    .D(_0162_),
    .Q(\inter_bp.report_shift_reg[3] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3666_ (.RESET_B(net788),
    .D(_0163_),
    .Q(\inter_bp.report_shift_reg[4] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _3667_ (.RESET_B(net782),
    .D(_0164_),
    .Q(\inter_bp.report_shift_reg[5] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3668_ (.RESET_B(net788),
    .D(_0165_),
    .Q(\inter_bp.report_shift_reg[6] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _3669_ (.RESET_B(net782),
    .D(_0166_),
    .Q(\inter_bp.report_shift_reg[7] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3670_ (.RESET_B(net788),
    .D(_0167_),
    .Q(\inter_bp.report_shift_reg[8] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _3671_ (.RESET_B(net782),
    .D(_0168_),
    .Q(\inter_bp.report_shift_reg[9] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3672_ (.RESET_B(net782),
    .D(_0169_),
    .Q(\inter_bp.report_shift_reg[10] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3673_ (.RESET_B(net782),
    .D(_0170_),
    .Q(\inter_bp.report_shift_reg[11] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _3674_ (.RESET_B(net780),
    .D(_0171_),
    .Q(\inter_bp.report_shift_reg[12] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _3675_ (.RESET_B(net782),
    .D(_0172_),
    .Q(\inter_bp.report_shift_reg[13] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _3676_ (.RESET_B(net780),
    .D(_0173_),
    .Q(\inter_bp.report_shift_reg[14] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _3677_ (.RESET_B(net780),
    .D(_0174_),
    .Q(\inter_bp.report_shift_reg[15] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _3678_ (.RESET_B(net780),
    .D(_0175_),
    .Q(\inter_bp.report_shift_reg[16] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _3679_ (.RESET_B(net780),
    .D(_0176_),
    .Q(\inter_bp.report_shift_reg[17] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _3680_ (.RESET_B(net780),
    .D(_0177_),
    .Q(\inter_bp.report_shift_reg[18] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _3681_ (.RESET_B(net782),
    .D(_0178_),
    .Q(\inter_bp.report_shift_reg[19] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _3682_ (.RESET_B(net790),
    .D(_0179_),
    .Q(\inter_bp.bp_report_addr_out[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _3683_ (.RESET_B(net788),
    .D(net402),
    .Q(\inter_bp.bp_report_addr_out[1] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _3684_ (.RESET_B(net788),
    .D(_0181_),
    .Q(\inter_bp.bp_report_addr_out[2] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3685_ (.RESET_B(net788),
    .D(net440),
    .Q(\inter_bp.bp_report_addr_out[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3686_ (.RESET_B(net789),
    .D(_0183_),
    .Q(\inter_bp.bp_report_addr_out[4] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3687_ (.RESET_B(net783),
    .D(_0184_),
    .Q(\inter_bp.bp_report_addr_out[5] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3688_ (.RESET_B(net789),
    .D(_0185_),
    .Q(\inter_bp.bp_report_addr_out[6] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _3689_ (.RESET_B(net783),
    .D(_0186_),
    .Q(\inter_bp.bp_report_addr_out[7] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3690_ (.RESET_B(net789),
    .D(_0187_),
    .Q(\inter_bp.bp_report_addr_out[8] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _3691_ (.RESET_B(net783),
    .D(_0188_),
    .Q(\inter_bp.bp_report_addr_out[9] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3692_ (.RESET_B(net783),
    .D(_0189_),
    .Q(\inter_bp.bp_report_addr_out[10] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _3693_ (.RESET_B(net780),
    .D(_0190_),
    .Q(\inter_bp.bp_report_addr_out[11] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _3694_ (.RESET_B(net780),
    .D(_0191_),
    .Q(\inter_bp.bp_report_addr_out[12] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _3695_ (.RESET_B(net782),
    .D(_0192_),
    .Q(\inter_bp.bp_report_addr_out[13] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _3696_ (.RESET_B(net781),
    .D(_0193_),
    .Q(\inter_bp.bp_report_addr_out[14] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _3697_ (.RESET_B(net781),
    .D(net436),
    .Q(\inter_bp.bp_report_addr_out[15] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _3698_ (.RESET_B(net781),
    .D(_0195_),
    .Q(\inter_bp.bp_report_addr_out[16] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _3699_ (.RESET_B(net781),
    .D(_0196_),
    .Q(\inter_bp.bp_report_addr_out[17] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3700_ (.RESET_B(net781),
    .D(net1002),
    .Q(\inter_bp.bp_report_addr_out[18] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _3701_ (.RESET_B(net781),
    .D(net981),
    .Q(\inter_bp.bp_report_addr_out[19] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3702_ (.RESET_B(net791),
    .D(_0199_),
    .Q(\inter_bp.report_receiving ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3703_ (.RESET_B(net763),
    .D(net522),
    .Q(\inter_bp.param_tx_counter[0] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _3704_ (.RESET_B(net763),
    .D(_0201_),
    .Q(\inter_bp.param_tx_counter[1] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _3705_ (.RESET_B(net763),
    .D(net272),
    .Q(\inter_bp.param_tx_counter[2] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _3706_ (.RESET_B(net763),
    .D(net916),
    .Q(\inter_bp.param_tx_counter[3] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _3707_ (.RESET_B(net763),
    .D(_0204_),
    .Q(\inter_bp.param_tx_counter[4] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _3708_ (.RESET_B(net757),
    .D(net289),
    .Q(\inter_bp.param_rx_counter[0] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _3709_ (.RESET_B(net757),
    .D(_0206_),
    .Q(\inter_bp.param_rx_counter[1] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _3710_ (.RESET_B(net757),
    .D(_0207_),
    .Q(\inter_bp.param_rx_counter[2] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _3711_ (.RESET_B(net757),
    .D(_0208_),
    .Q(\inter_bp.param_rx_counter[3] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _3712_ (.RESET_B(net757),
    .D(_0209_),
    .Q(\inter_bp.param_rx_counter[4] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _3713_ (.RESET_B(net789),
    .D(net747),
    .Q(\inter_bp.bp_report_valid_out ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3714_ (.RESET_B(net796),
    .D(net58),
    .Q(\inter_bp.serialize_param_valid_prev ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _3715_ (.RESET_B(net764),
    .D(net1069),
    .Q(\inter_bp.param_transmitting ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _3716_ (.RESET_B(net762),
    .D(net231),
    .Q(\inter_bp.param_rx_done ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _3717_ (.RESET_B(net794),
    .D(net161),
    .Q(\inter_bp.param_tx_shift_reg[0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _3718_ (.RESET_B(net793),
    .D(net181),
    .Q(\inter_bp.param_tx_shift_reg[1] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _3719_ (.RESET_B(net829),
    .D(net233),
    .Q(\inter_bp.param_tx_shift_reg[2] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _3720_ (.RESET_B(net828),
    .D(net244),
    .Q(\inter_bp.param_tx_shift_reg[3] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _3721_ (.RESET_B(net834),
    .D(net302),
    .Q(\inter_bp.param_tx_shift_reg[4] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _3722_ (.RESET_B(net833),
    .D(_0215_),
    .Q(\inter_bp.param_tx_shift_reg[5] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _3723_ (.RESET_B(net836),
    .D(net269),
    .Q(\inter_bp.param_tx_shift_reg[6] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _3724_ (.RESET_B(net836),
    .D(net101),
    .Q(\inter_bp.param_tx_shift_reg[7] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _3725_ (.RESET_B(net836),
    .D(_0218_),
    .Q(\inter_bp.param_tx_shift_reg[8] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _3726_ (.RESET_B(net824),
    .D(_0219_),
    .Q(\inter_bp.param_tx_shift_reg[9] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _3727_ (.RESET_B(net825),
    .D(_0220_),
    .Q(\inter_bp.param_tx_shift_reg[10] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3728_ (.RESET_B(net824),
    .D(net106),
    .Q(\inter_bp.param_tx_shift_reg[11] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _3729_ (.RESET_B(net824),
    .D(_0222_),
    .Q(\inter_bp.param_tx_shift_reg[12] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3730_ (.RESET_B(net824),
    .D(net61),
    .Q(\inter_bp.param_tx_shift_reg[13] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3731_ (.RESET_B(net824),
    .D(_0224_),
    .Q(\inter_bp.param_tx_shift_reg[14] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3732_ (.RESET_B(net822),
    .D(_0225_),
    .Q(\inter_bp.param_tx_shift_reg[15] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3733_ (.RESET_B(net821),
    .D(net73),
    .Q(\inter_bp.param_tx_shift_reg[16] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _3734_ (.RESET_B(net814),
    .D(_0227_),
    .Q(\inter_bp.param_tx_shift_reg[17] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _3735_ (.RESET_B(net814),
    .D(net191),
    .Q(\inter_bp.param_tx_shift_reg[18] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _3736_ (.RESET_B(net814),
    .D(net79),
    .Q(\inter_bp.param_tx_shift_reg[19] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _3737_ (.RESET_B(net813),
    .D(net138),
    .Q(\inter_bp.param_tx_shift_reg[20] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _3738_ (.RESET_B(net813),
    .D(_0231_),
    .Q(\inter_bp.param_tx_shift_reg[21] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _3739_ (.RESET_B(net814),
    .D(net222),
    .Q(\inter_bp.param_tx_shift_reg[22] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _3740_ (.RESET_B(net813),
    .D(net68),
    .Q(\inter_bp.param_tx_shift_reg[23] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _3741_ (.RESET_B(net815),
    .D(_0234_),
    .Q(\inter_bp.param_tx_shift_reg[24] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _3742_ (.RESET_B(net813),
    .D(net63),
    .Q(\inter_bp.param_tx_shift_reg[25] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _3743_ (.RESET_B(net821),
    .D(net163),
    .Q(\inter_bp.param_tx_shift_reg[26] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _3744_ (.RESET_B(net815),
    .D(_0237_),
    .Q(\inter_bp.param_tx_shift_reg[27] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _3745_ (.RESET_B(net821),
    .D(_0238_),
    .Q(\inter_bp.param_tx_shift_reg[28] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _3746_ (.RESET_B(net815),
    .D(_0239_),
    .Q(\inter_bp.param_tx_shift_reg[29] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _3747_ (.RESET_B(net821),
    .D(net99),
    .Q(\inter_bp.param_tx_shift_reg[30] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _3748_ (.RESET_B(net815),
    .D(net140),
    .Q(\inter_bp.param_tx_shift_reg[31] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _3749_ (.RESET_B(net815),
    .D(net83),
    .Q(\inter_bp.param_tx_shift_reg[32] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _3750_ (.RESET_B(net815),
    .D(net128),
    .Q(\inter_bp.param_tx_shift_reg[33] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _3751_ (.RESET_B(net815),
    .D(net112),
    .Q(\inter_bp.param_tx_shift_reg[34] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _3752_ (.RESET_B(net814),
    .D(net189),
    .Q(\inter_bp.param_tx_shift_reg[35] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _3753_ (.RESET_B(net813),
    .D(net93),
    .Q(\inter_bp.param_tx_shift_reg[36] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _3754_ (.RESET_B(net813),
    .D(net176),
    .Q(\inter_bp.param_tx_shift_reg[37] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _3755_ (.RESET_B(net813),
    .D(net97),
    .Q(\inter_bp.param_tx_shift_reg[38] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _3756_ (.RESET_B(net777),
    .D(net391),
    .Q(\inter_bp.param_tx_shift_reg[39] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _3757_ (.RESET_B(net826),
    .D(_0250_),
    .Q(\inter_bp.param_tx_shift_reg[40] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _3758_ (.RESET_B(net826),
    .D(net95),
    .Q(\inter_bp.param_tx_shift_reg[41] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _3759_ (.RESET_B(net826),
    .D(net91),
    .Q(\inter_bp.param_tx_shift_reg[42] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _3760_ (.RESET_B(net827),
    .D(_0253_),
    .Q(\inter_bp.param_tx_shift_reg[43] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _3761_ (.RESET_B(net826),
    .D(net214),
    .Q(\inter_bp.param_tx_shift_reg[44] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _3762_ (.RESET_B(net827),
    .D(_0255_),
    .Q(\inter_bp.param_tx_shift_reg[45] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _3763_ (.RESET_B(net826),
    .D(_0256_),
    .Q(\inter_bp.param_tx_shift_reg[46] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _3764_ (.RESET_B(net827),
    .D(_0257_),
    .Q(\inter_bp.param_tx_shift_reg[47] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _3765_ (.RESET_B(net793),
    .D(net557),
    .Q(\inter_bp.report_tx_counter[0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_2 _3766_ (.RESET_B(net793),
    .D(_0259_),
    .Q(\inter_bp.report_tx_counter[1] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3767_ (.RESET_B(net793),
    .D(net327),
    .Q(\inter_bp.report_tx_counter[2] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3768_ (.RESET_B(net793),
    .D(net1009),
    .Q(\inter_bp.report_tx_counter[3] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3769_ (.RESET_B(net793),
    .D(_0262_),
    .Q(\inter_bp.report_tx_counter[4] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3770_ (.RESET_B(net773),
    .D(net1015),
    .Q(\bp_core.bp_stride_in[0] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _3771_ (.RESET_B(net769),
    .D(net857),
    .Q(\bp_core.bp_stride_in[1] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _3772_ (.RESET_B(net807),
    .D(net564),
    .Q(\bp_core.bp_stride_in[2] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _3773_ (.RESET_B(net760),
    .D(_0086_),
    .Q(\bp_core.bp_stride_in[3] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _3774_ (.RESET_B(net807),
    .D(_0087_),
    .Q(\bp_core.bp_stride_in[4] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _3775_ (.RESET_B(net760),
    .D(_0088_),
    .Q(\bp_core.bp_stride_in[5] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _3776_ (.RESET_B(net807),
    .D(net872),
    .Q(\bp_core.bp_stride_in[6] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _3777_ (.RESET_B(net760),
    .D(_0090_),
    .Q(\bp_core.bp_stride_in[7] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _3778_ (.RESET_B(net808),
    .D(_0091_),
    .Q(\bp_core.bp_stride_in[8] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _3779_ (.RESET_B(net761),
    .D(net962),
    .Q(\bp_core.bp_stride_in[9] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _3780_ (.RESET_B(net774),
    .D(_0074_),
    .Q(\bp_core.bp_stride_in[10] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _3781_ (.RESET_B(net766),
    .D(net428),
    .Q(\bp_core.bp_stride_in[11] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _3782_ (.RESET_B(net774),
    .D(_0076_),
    .Q(\bp_core.bp_stride_in[12] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _3783_ (.RESET_B(net761),
    .D(_0077_),
    .Q(\bp_core.bp_stride_in[13] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _3784_ (.RESET_B(net772),
    .D(_0078_),
    .Q(\bp_core.bp_stride_in[14] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _3785_ (.RESET_B(net761),
    .D(_0079_),
    .Q(\bp_core.bp_stride_in[15] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _3786_ (.RESET_B(net771),
    .D(_0080_),
    .Q(\bp_core.bp_stride_in[16] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _3787_ (.RESET_B(net766),
    .D(_0081_),
    .Q(\bp_core.bp_stride_in[17] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _3788_ (.RESET_B(net771),
    .D(_0082_),
    .Q(\bp_core.bp_stride_in[18] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _3789_ (.RESET_B(net766),
    .D(_0083_),
    .Q(\bp_core.bp_stride_in[19] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _3790_ (.RESET_B(net801),
    .D(net57),
    .Q(\inter_bp.serialize_report_valid_prev ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _3791_ (.RESET_B(net766),
    .D(net969),
    .Q(\inter_bp.param_pending ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _3792_ (.RESET_B(net794),
    .D(_0097_),
    .Q(\inter_bp.report_transmitting ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3793_ (.RESET_B(net793),
    .D(net184),
    .Q(\inter_bp.report_tx_shift_reg[0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _3794_ (.RESET_B(net793),
    .D(net249),
    .Q(\inter_bp.report_tx_shift_reg[1] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _3795_ (.RESET_B(net794),
    .D(net166),
    .Q(\inter_bp.report_tx_shift_reg[2] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3796_ (.RESET_B(net792),
    .D(net187),
    .Q(\inter_bp.report_tx_shift_reg[3] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _3797_ (.RESET_B(net794),
    .D(net117),
    .Q(\inter_bp.report_tx_shift_reg[4] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _3798_ (.RESET_B(net792),
    .D(net71),
    .Q(\inter_bp.report_tx_shift_reg[5] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _3799_ (.RESET_B(net794),
    .D(net210),
    .Q(\inter_bp.report_tx_shift_reg[6] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3800_ (.RESET_B(net785),
    .D(net126),
    .Q(\inter_bp.report_tx_shift_reg[7] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3801_ (.RESET_B(net792),
    .D(net76),
    .Q(\inter_bp.report_tx_shift_reg[8] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3802_ (.RESET_B(net785),
    .D(net147),
    .Q(\inter_bp.report_tx_shift_reg[9] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _3803_ (.RESET_B(net787),
    .D(net66),
    .Q(\inter_bp.report_tx_shift_reg[10] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _3804_ (.RESET_B(net785),
    .D(net119),
    .Q(\inter_bp.report_tx_shift_reg[11] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _3805_ (.RESET_B(net787),
    .D(net205),
    .Q(\inter_bp.report_tx_shift_reg[12] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _3806_ (.RESET_B(net785),
    .D(net110),
    .Q(\inter_bp.report_tx_shift_reg[13] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _3807_ (.RESET_B(net797),
    .D(net277),
    .Q(\inter_bp.report_tx_shift_reg[14] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _3808_ (.RESET_B(net787),
    .D(net151),
    .Q(\inter_bp.report_tx_shift_reg[15] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3809_ (.RESET_B(net797),
    .D(net134),
    .Q(\inter_bp.report_tx_shift_reg[16] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _3810_ (.RESET_B(net786),
    .D(net158),
    .Q(\inter_bp.report_tx_shift_reg[17] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3811_ (.RESET_B(net796),
    .D(_0281_),
    .Q(\inter_bp.report_tx_shift_reg[18] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _3812_ (.RESET_B(net786),
    .D(_0282_),
    .Q(\inter_bp.report_tx_shift_reg[19] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _3813_ (.RESET_B(net798),
    .D(_0283_),
    .Q(\bp_core.params_module.counter[0] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _3814_ (.RESET_B(net798),
    .D(_0284_),
    .Q(\bp_core.params_module.counter[1] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _3815_ (.RESET_B(net798),
    .D(_0285_),
    .Q(\bp_core.params_module.counter[2] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _3816_ (.RESET_B(net778),
    .D(_0286_),
    .Q(\bp_core.params_module.counter[3] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _3817_ (.RESET_B(net762),
    .D(net997),
    .Q(\inter_bp.param_receiving ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _3818_ (.RESET_B(net798),
    .D(_0103_),
    .Q(_0098_),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _3819_ (.RESET_B(net798),
    .D(_0000_),
    .Q(\bp_core.params_module.state[1] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _3820_ (.RESET_B(net798),
    .D(_0001_),
    .Q(\bp_core.params_module.state[2] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _3821_ (.RESET_B(net796),
    .D(_0002_),
    .Q(\bp_core.params_module.state[3] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _3822_ (.RESET_B(net803),
    .D(_0288_),
    .Q(\bp_core.threshold_reg[5] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3823_ (.RESET_B(net803),
    .D(net425),
    .Q(_0099_),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3824_ (.RESET_B(net803),
    .D(net422),
    .Q(_0100_),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _3825_ (.RESET_B(net808),
    .D(_0291_),
    .Q(\bp_core.bp_stride_out[5] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _3826_ (.RESET_B(net808),
    .D(net1176),
    .Q(\bp_core.bp_stride_out[6] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _3827_ (.RESET_B(net808),
    .D(_0293_),
    .Q(\bp_core.bp_stride_out[7] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _3828_ (.RESET_B(net809),
    .D(_0294_),
    .Q(\bp_core.bp_stride_out[8] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _3829_ (.RESET_B(net808),
    .D(_0295_),
    .Q(\bp_core.bp_stride_out[9] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _3830_ (.RESET_B(net778),
    .D(net1161),
    .Q(\bp_core.bp_lambda_out[0] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _3831_ (.RESET_B(net778),
    .D(net1124),
    .Q(\bp_core.bp_lambda_out[1] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _3832_ (.RESET_B(net796),
    .D(_0298_),
    .Q(\bp_core.bp_lambda_out[2] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _3833_ (.RESET_B(net776),
    .D(net1178),
    .Q(\bp_core.bp_lambda_out[3] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _3834_ (.RESET_B(net775),
    .D(_0300_),
    .Q(\bp_core.bp_lambda_out[4] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _3835_ (.RESET_B(net813),
    .D(_0301_),
    .Q(\bp_core.bp_stride_out[10] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _3836_ (.RESET_B(net777),
    .D(net513),
    .Q(\bp_core.bp_stride_out[11] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _3837_ (.RESET_B(net777),
    .D(_0303_),
    .Q(\bp_core.bp_stride_out[12] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _3838_ (.RESET_B(net777),
    .D(_0304_),
    .Q(\bp_core.bp_stride_out[13] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _3839_ (.RESET_B(net777),
    .D(_0305_),
    .Q(\bp_core.bp_stride_out[14] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _3840_ (.RESET_B(net826),
    .D(net1159),
    .Q(\bp_core.bp_lambda_out[5] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _3841_ (.RESET_B(net826),
    .D(_0307_),
    .Q(\bp_core.bp_lambda_out[6] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _3842_ (.RESET_B(net826),
    .D(_0308_),
    .Q(\bp_core.bp_lambda_out[7] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _3843_ (.RESET_B(net829),
    .D(net1060),
    .Q(\bp_addr_out[0] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _3844_ (.RESET_B(net827),
    .D(_0310_),
    .Q(\bp_addr_out[1] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _3845_ (.RESET_B(net828),
    .D(_0311_),
    .Q(\bp_addr_out[2] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _3846_ (.RESET_B(net828),
    .D(net1103),
    .Q(\bp_addr_out[3] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _3847_ (.RESET_B(net828),
    .D(_0313_),
    .Q(\bp_addr_out[4] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _3848_ (.RESET_B(net833),
    .D(net1096),
    .Q(\bp_addr_out[5] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _3849_ (.RESET_B(net833),
    .D(net1113),
    .Q(\bp_addr_out[6] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3850_ (.RESET_B(net836),
    .D(net1090),
    .Q(\bp_addr_out[7] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3851_ (.RESET_B(net833),
    .D(net1074),
    .Q(\bp_addr_out[8] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3852_ (.RESET_B(net824),
    .D(_0318_),
    .Q(\bp_addr_out[9] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3853_ (.RESET_B(net822),
    .D(_0319_),
    .Q(\bp_addr_out[10] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _3854_ (.RESET_B(net822),
    .D(net1082),
    .Q(\bp_addr_out[11] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _3855_ (.RESET_B(net822),
    .D(net1078),
    .Q(\bp_addr_out[12] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _3856_ (.RESET_B(net822),
    .D(net1088),
    .Q(\bp_addr_out[13] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _3857_ (.RESET_B(net816),
    .D(net1105),
    .Q(\bp_addr_out[14] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _3858_ (.RESET_B(net814),
    .D(net1048),
    .Q(\bp_addr_out[15] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _3859_ (.RESET_B(net778),
    .D(net1020),
    .Q(\bp_addr_out[16] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _3860_ (.RESET_B(net814),
    .D(_0326_),
    .Q(\bp_addr_out[17] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _3861_ (.RESET_B(net778),
    .D(net1066),
    .Q(\bp_addr_out[18] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _3862_ (.RESET_B(net778),
    .D(net1039),
    .Q(\bp_addr_out[19] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _3863_ (.RESET_B(net797),
    .D(net59),
    .Q(\bp_core.bp_param_output_valid ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _3864_ (.RESET_B(net797),
    .D(net199),
    .Q(\bp_core.bp_param_valid_out ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _3865_ (.RESET_B(net777),
    .D(_0330_),
    .Q(\bp_core.bp_stride_out[15] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _3866_ (.RESET_B(net775),
    .D(_0331_),
    .Q(\bp_core.bp_stride_out[16] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _3867_ (.RESET_B(net775),
    .D(_0332_),
    .Q(\bp_core.bp_stride_out[17] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _3868_ (.RESET_B(net775),
    .D(_0333_),
    .Q(\bp_core.bp_stride_out[18] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _3869_ (.RESET_B(net777),
    .D(_0334_),
    .Q(\bp_core.bp_stride_out[19] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _3870_ (.RESET_B(net797),
    .D(net460),
    .Q(\bp_core.bp_param_output_data[0] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _3871_ (.RESET_B(net802),
    .D(net291),
    .Q(\bp_core.bp_param_output_data[1] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _3872_ (.RESET_B(net797),
    .D(net953),
    .Q(\bp_core.bp_param_output_data[2] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _3873_ (.RESET_B(net799),
    .D(net297),
    .Q(\bp_core.bp_param_output_data[3] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _3874_ (.RESET_B(net797),
    .D(net960),
    .Q(\bp_core.bp_param_output_data[4] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _3875_ (.RESET_B(net799),
    .D(net924),
    .Q(\bp_core.params_module.params_ready ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _3876_ (.RESET_B(net799),
    .D(\bp_core.params_module.state[0] ),
    .Q(\bp_core.params_done ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _3877_ (.RESET_B(net774),
    .D(net1025),
    .Q(\bp_core.params_addr[15] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _3878_ (.RESET_B(net771),
    .D(net975),
    .Q(\bp_core.params_addr[16] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _3879_ (.RESET_B(net771),
    .D(_0342_),
    .Q(\bp_core.params_addr[17] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _3880_ (.RESET_B(net775),
    .D(net878),
    .Q(\bp_core.params_addr[18] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _3881_ (.RESET_B(net771),
    .D(_0344_),
    .Q(\bp_core.params_addr[19] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _3882_ (.RESET_B(net831),
    .D(net251),
    .Q(\bp_core.data_reg[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3883_ (.RESET_B(net830),
    .D(net413),
    .Q(\bp_core.data_reg[1] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3884_ (.RESET_B(net830),
    .D(net365),
    .Q(\bp_core.data_reg[2] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3885_ (.RESET_B(net830),
    .D(_0348_),
    .Q(\bp_core.data_reg[3] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3886_ (.RESET_B(net831),
    .D(net348),
    .Q(\bp_core.data_reg[4] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3887_ (.RESET_B(net803),
    .D(net361),
    .Q(\bp_core.data_reg[5] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3888_ (.RESET_B(net804),
    .D(_0351_),
    .Q(\bp_core.data_reg[6] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _3889_ (.RESET_B(net802),
    .D(net385),
    .Q(\bp_core.data_reg[7] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _3890_ (.RESET_B(net827),
    .D(net1135),
    .Q(\bp_core.addr_reg[0] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _3891_ (.RESET_B(net827),
    .D(_0354_),
    .Q(\bp_core.addr_reg[1] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _3892_ (.RESET_B(net828),
    .D(_0355_),
    .Q(\bp_core.addr_reg[2] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _3893_ (.RESET_B(net828),
    .D(net1107),
    .Q(\bp_core.addr_reg[3] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _3894_ (.RESET_B(net828),
    .D(_0357_),
    .Q(\bp_core.addr_reg[4] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _3895_ (.RESET_B(net833),
    .D(_0358_),
    .Q(\bp_core.addr_reg[5] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3896_ (.RESET_B(net833),
    .D(_0359_),
    .Q(\bp_core.addr_reg[6] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3897_ (.RESET_B(net833),
    .D(net1131),
    .Q(\bp_core.addr_reg[7] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3898_ (.RESET_B(net833),
    .D(_0361_),
    .Q(\bp_core.addr_reg[8] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _3899_ (.RESET_B(net822),
    .D(_0362_),
    .Q(\bp_core.addr_reg[9] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _3900_ (.RESET_B(net823),
    .D(net1062),
    .Q(\bp_core.addr_reg[10] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _3901_ (.RESET_B(net822),
    .D(net1116),
    .Q(\bp_core.addr_reg[11] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _3902_ (.RESET_B(net822),
    .D(_0365_),
    .Q(\bp_core.addr_reg[12] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _3903_ (.RESET_B(net816),
    .D(_0366_),
    .Q(\bp_core.addr_reg[13] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _3904_ (.RESET_B(net828),
    .D(_0367_),
    .Q(\bp_core.addr_reg[14] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _3905_ (.RESET_B(net827),
    .D(_0368_),
    .Q(\bp_core.addr_reg[15] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _3906_ (.RESET_B(net776),
    .D(_0369_),
    .Q(\bp_core.addr_reg[16] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _3907_ (.RESET_B(net776),
    .D(_0370_),
    .Q(\bp_core.addr_reg[17] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _3908_ (.RESET_B(net776),
    .D(net483),
    .Q(\bp_core.addr_reg[18] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _3909_ (.RESET_B(net796),
    .D(_0372_),
    .Q(\bp_core.addr_reg[19] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _3910_ (.RESET_B(net798),
    .D(_0037_),
    .Q(\bp_core.params_module.start_load ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _3911_ (.RESET_B(net801),
    .D(net455),
    .Q(\bp_core.busy_out ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _3912_ (.RESET_B(net838),
    .D(_0374_),
    .Q(\bp_core.init_counter[0] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _3913_ (.RESET_B(net839),
    .D(_0375_),
    .Q(\bp_core.init_counter[1] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _3914_ (.RESET_B(net839),
    .D(_0376_),
    .Q(\bp_core.init_counter[2] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _3915_ (.RESET_B(net839),
    .D(_0377_),
    .Q(\bp_core.init_counter[3] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_2 _3916_ (.RESET_B(net835),
    .D(_0378_),
    .Q(\bp_core.init_counter[4] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _3917_ (.RESET_B(net835),
    .D(_0379_),
    .Q(\bp_core.init_counter[5] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _3918_ (.RESET_B(net837),
    .D(_0380_),
    .Q(\bp_core.init_counter[6] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _3919_ (.RESET_B(net836),
    .D(_0381_),
    .Q(\bp_core.init_counter[7] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_2 _3920_ (.RESET_B(net836),
    .D(_0382_),
    .Q(\bp_core.init_counter[8] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _3921_ (.RESET_B(net836),
    .D(net481),
    .Q(\bp_core.init_counter[9] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _3922_ (.RESET_B(net834),
    .D(_0384_),
    .Q(\bp_core.init_counter[10] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_2 _3923_ (.RESET_B(net834),
    .D(_0385_),
    .Q(\bp_core.init_counter[11] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _3924_ (.RESET_B(net834),
    .D(_0386_),
    .Q(\bp_core.init_counter[12] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _3925_ (.RESET_B(net834),
    .D(_0387_),
    .Q(\bp_core.init_counter[13] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _3926_ (.RESET_B(net832),
    .D(_0388_),
    .Q(\bp_core.init_counter[14] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _3927_ (.RESET_B(net831),
    .D(net370),
    .Q(\bp_core.init_counter[15] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _3928_ (.RESET_B(net801),
    .D(net354),
    .Q(\bp_core.status_out[0] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _3929_ (.RESET_B(net801),
    .D(net383),
    .Q(\bp_core.status_out[1] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _3930_ (.RESET_B(net801),
    .D(_0040_),
    .Q(\bp_core.status_out[2] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _3931_ (.RESET_B(net801),
    .D(net352),
    .Q(\bp_core.status_out[3] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _3932_ (.RESET_B(net801),
    .D(_0042_),
    .Q(\bp_core.status_out[4] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _3933_ (.RESET_B(net798),
    .D(_0036_),
    .Q(\bp_core.bp_param_ack_out ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _3934_ (.RESET_B(net801),
    .D(_0043_),
    .Q(\bp_core.valid_out ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _3935_ (.RESET_B(net803),
    .D(_0390_),
    .Q(\bp_core.threshold_load_counter ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _3936_ (.RESET_B(net832),
    .D(net880),
    .Q(\bp_core.ram_we ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _3937_ (.RESET_B(net799),
    .D(_0035_),
    .Q(\bp_core.params_forward ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _3938_ (.RESET_B(net805),
    .D(net345),
    .Q(\bp_core.bp_report_addr_out[0] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3939_ (.RESET_B(net792),
    .D(_0025_),
    .Q(\bp_core.bp_report_addr_out[1] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3940_ (.RESET_B(net805),
    .D(_0026_),
    .Q(\bp_core.bp_report_addr_out[2] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3941_ (.RESET_B(net792),
    .D(net848),
    .Q(\bp_core.bp_report_addr_out[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3942_ (.RESET_B(net792),
    .D(_0028_),
    .Q(\bp_core.bp_report_addr_out[4] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3943_ (.RESET_B(net785),
    .D(net283),
    .Q(\bp_core.bp_report_addr_out[5] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3944_ (.RESET_B(net792),
    .D(net330),
    .Q(\bp_core.bp_report_addr_out[6] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3945_ (.RESET_B(net785),
    .D(net263),
    .Q(\bp_core.bp_report_addr_out[7] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3946_ (.RESET_B(net792),
    .D(net300),
    .Q(\bp_core.bp_report_addr_out[8] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _3947_ (.RESET_B(net786),
    .D(net280),
    .Q(\bp_core.bp_report_addr_out[9] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _3948_ (.RESET_B(net785),
    .D(net338),
    .Q(\bp_core.bp_report_addr_out[10] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _3949_ (.RESET_B(net786),
    .D(net443),
    .Q(\bp_core.bp_report_addr_out[11] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3950_ (.RESET_B(net786),
    .D(net393),
    .Q(\bp_core.bp_report_addr_out[12] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _3951_ (.RESET_B(net785),
    .D(net256),
    .Q(\bp_core.bp_report_addr_out[13] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3952_ (.RESET_B(net786),
    .D(net415),
    .Q(\bp_core.bp_report_addr_out[14] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _3953_ (.RESET_B(net786),
    .D(net287),
    .Q(\bp_core.bp_report_addr_out[15] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3954_ (.RESET_B(net796),
    .D(net343),
    .Q(\bp_core.bp_report_addr_out[16] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _3955_ (.RESET_B(net786),
    .D(net933),
    .Q(\bp_core.bp_report_addr_out[17] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _3956_ (.RESET_B(net796),
    .D(net973),
    .Q(\bp_core.bp_report_addr_out[18] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _3957_ (.RESET_B(net796),
    .D(_0024_),
    .Q(\bp_core.bp_report_addr_out[19] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _3958_ (.RESET_B(net805),
    .D(_0034_),
    .Q(\bp_core.bp_report_valid_out ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _3959_ (.RESET_B(net832),
    .D(_1799_[0]),
    .Q(\bp_core.ram_start ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _3960_ (.RESET_B(net831),
    .D(net358),
    .Q(\bp_core.ram_wdata[0] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _3961_ (.RESET_B(net830),
    .D(net457),
    .Q(\bp_core.ram_wdata[1] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3962_ (.RESET_B(net830),
    .D(_0394_),
    .Q(\bp_core.ram_wdata[2] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _3963_ (.RESET_B(net830),
    .D(_0395_),
    .Q(\bp_core.ram_wdata[3] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _3964_ (.RESET_B(net830),
    .D(_0396_),
    .Q(\bp_core.ram_wdata[4] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _3965_ (.RESET_B(net830),
    .D(net311),
    .Q(\bp_core.ram_wdata[5] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _3966_ (.RESET_B(net831),
    .D(_0398_),
    .Q(\bp_core.ram_wdata[6] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _3967_ (.RESET_B(net831),
    .D(net356),
    .Q(\bp_core.ram_wdata[7] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _3968_ (.RESET_B(net838),
    .D(net220),
    .Q(\bp_core.ram_addr[0] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _3969_ (.RESET_B(net839),
    .D(net149),
    .Q(\bp_core.ram_addr[1] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _3970_ (.RESET_B(net838),
    .D(net114),
    .Q(\bp_core.ram_addr[2] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _3971_ (.RESET_B(net839),
    .D(net153),
    .Q(\bp_core.ram_addr[3] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _3972_ (.RESET_B(net838),
    .D(net170),
    .Q(\bp_core.ram_addr[4] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _3973_ (.RESET_B(net835),
    .D(net155),
    .Q(\bp_core.ram_addr[5] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _3974_ (.RESET_B(net835),
    .D(net121),
    .Q(\bp_core.ram_addr[6] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _3975_ (.RESET_B(net835),
    .D(net123),
    .Q(\bp_core.ram_addr[7] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _3976_ (.RESET_B(net835),
    .D(net108),
    .Q(\bp_core.ram_addr[8] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _3977_ (.RESET_B(net835),
    .D(net193),
    .Q(\bp_core.ram_addr[9] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _3978_ (.RESET_B(net835),
    .D(net178),
    .Q(\bp_core.ram_addr[10] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _3979_ (.RESET_B(net834),
    .D(net195),
    .Q(\bp_core.ram_addr[11] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _3980_ (.RESET_B(net834),
    .D(net174),
    .Q(\bp_core.ram_addr[12] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _3981_ (.RESET_B(net838),
    .D(net132),
    .Q(\bp_core.ram_addr[13] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _3982_ (.RESET_B(net832),
    .D(net142),
    .Q(\bp_core.ram_addr[14] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _3983_ (.RESET_B(net832),
    .D(net172),
    .Q(\bp_core.ram_addr[15] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _3984_ (.RESET_B(net803),
    .D(_0416_),
    .Q(\bp_core.threshold_reg[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3985_ (.RESET_B(net804),
    .D(_0417_),
    .Q(\bp_core.threshold_reg[1] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _3986_ (.RESET_B(net804),
    .D(net517),
    .Q(\bp_core.threshold_reg[2] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _3987_ (.RESET_B(net803),
    .D(_0419_),
    .Q(_0101_),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3988_ (.RESET_B(net803),
    .D(_0420_),
    .Q(\bp_core.threshold_reg[4] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _3989_ (.RESET_B(net802),
    .D(net865),
    .Q(\bp_core.initialized ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _3990_ (.RESET_B(net808),
    .D(_0422_),
    .Q(\bp_core.bp_stride_out[0] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _3991_ (.RESET_B(net808),
    .D(net1139),
    .Q(\bp_core.bp_stride_out[1] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _3992_ (.RESET_B(net809),
    .D(_0424_),
    .Q(\bp_core.bp_stride_out[2] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _3993_ (.RESET_B(net808),
    .D(_0425_),
    .Q(\bp_core.bp_stride_out[3] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _3994_ (.RESET_B(net809),
    .D(_0426_),
    .Q(\bp_core.bp_stride_out[4] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _3995_ (.RESET_B(net47),
    .D(_0427_),
    .Q(\spi_ctrl.addr[0] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _3996_ (.RESET_B(net46),
    .D(net307),
    .Q(\spi_ctrl.addr[1] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _3997_ (.RESET_B(net45),
    .D(_0429_),
    .Q(\spi_ctrl.addr[2] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _3998_ (.RESET_B(net44),
    .D(net314),
    .Q(\spi_ctrl.addr[3] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _3999_ (.RESET_B(net43),
    .D(_0431_),
    .Q(\spi_ctrl.addr[4] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _4000_ (.RESET_B(net42),
    .D(_0432_),
    .Q(\spi_ctrl.addr[5] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4001_ (.RESET_B(net41),
    .D(_0433_),
    .Q(\spi_ctrl.addr[6] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4002_ (.RESET_B(net40),
    .D(_0434_),
    .Q(\spi_ctrl.addr[7] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4003_ (.RESET_B(net39),
    .D(_0435_),
    .Q(\spi_ctrl.addr[8] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4004_ (.RESET_B(net38),
    .D(_0436_),
    .Q(\spi_ctrl.addr[9] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4005_ (.RESET_B(net37),
    .D(_0437_),
    .Q(\spi_ctrl.addr[10] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _4006_ (.RESET_B(net36),
    .D(net340),
    .Q(\spi_ctrl.addr[11] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _4007_ (.RESET_B(net35),
    .D(net379),
    .Q(\spi_ctrl.addr[12] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _4008_ (.RESET_B(net34),
    .D(net240),
    .Q(\spi_ctrl.addr[13] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4009_ (.RESET_B(net33),
    .D(net237),
    .Q(\spi_ctrl.addr[14] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4010_ (.RESET_B(net32),
    .D(net253),
    .Q(\spi_ctrl.addr[15] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _4011_ (.RESET_B(net819),
    .D(_0443_),
    .Q(\bp_core.params_addr[10] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4012_ (.RESET_B(net819),
    .D(_0444_),
    .Q(\bp_core.params_addr[11] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4013_ (.RESET_B(net819),
    .D(_0445_),
    .Q(\bp_core.params_addr[12] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4014_ (.RESET_B(net811),
    .D(_0446_),
    .Q(\bp_core.params_addr[13] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4015_ (.RESET_B(net811),
    .D(_0447_),
    .Q(\bp_core.params_addr[14] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _4016_ (.RESET_B(net821),
    .D(_0448_),
    .Q(\bp_core.params_addr[5] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4017_ (.RESET_B(net821),
    .D(_0449_),
    .Q(\bp_core.params_addr[6] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4018_ (.RESET_B(net821),
    .D(_0450_),
    .Q(\bp_core.params_addr[7] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _4019_ (.RESET_B(net823),
    .D(_0451_),
    .Q(\bp_core.params_addr[8] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _4020_ (.RESET_B(net823),
    .D(net958),
    .Q(\bp_core.params_addr[9] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_2 _4021_ (.RESET_B(net802),
    .D(_0104_),
    .Q(_0102_),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _4022_ (.RESET_B(net831),
    .D(_0005_),
    .Q(\bp_core.state[1] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4023_ (.RESET_B(net799),
    .D(net964),
    .Q(\bp_core.state[2] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _4024_ (.RESET_B(net804),
    .D(_0007_),
    .Q(\bp_core.state[3] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _4025_ (.RESET_B(net799),
    .D(net944),
    .Q(\bp_core.state[4] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _4026_ (.RESET_B(net799),
    .D(_0009_),
    .Q(\bp_core.state[5] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _4027_ (.RESET_B(net802),
    .D(net293),
    .Q(\bp_core.state[6] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4028_ (.RESET_B(net832),
    .D(_0011_),
    .Q(\bp_core.state[7] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _4029_ (.RESET_B(net799),
    .D(net168),
    .Q(\bp_core.state[8] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _4030_ (.RESET_B(net802),
    .D(_0013_),
    .Q(\bp_core.state[9] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _4031_ (.RESET_B(net802),
    .D(net216),
    .Q(\bp_core.state[10] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4032_ (.RESET_B(net802),
    .D(net930),
    .Q(\bp_core.state[11] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _4033_ (.RESET_B(net778),
    .D(net434),
    .Q(\bp_core.params_addr[0] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _4034_ (.RESET_B(net821),
    .D(net1017),
    .Q(\bp_core.params_addr[1] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _4035_ (.RESET_B(net816),
    .D(net956),
    .Q(\bp_core.params_addr[2] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _4036_ (.RESET_B(net815),
    .D(_0456_),
    .Q(\bp_core.params_addr[3] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _4037_ (.RESET_B(net816),
    .D(net987),
    .Q(\bp_core.params_addr[4] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _4038_ (.RESET_B(net31),
    .D(net381),
    .Q(\spi_ctrl.bits_remaining[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4039_ (.RESET_B(net30),
    .D(_0459_),
    .Q(\spi_ctrl.bits_remaining[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4040_ (.RESET_B(net29),
    .D(net226),
    .Q(\spi_ctrl.bits_remaining[2] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4041_ (.RESET_B(net28),
    .D(_0461_),
    .Q(\spi_ctrl.bits_remaining[3] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _4042_ (.RESET_B(net27),
    .D(_0462_),
    .Q(\spi_ctrl.fsm_state[0] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _4043_ (.RESET_B(net26),
    .D(_0463_),
    .Q(\spi_ctrl.fsm_state[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _4044_ (.RESET_B(net25),
    .D(net407),
    .Q(\spi_ctrl.writing ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _4045_ (.RESET_B(net24),
    .D(net1071),
    .Q(\bp_core.ram_rdata[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _4046_ (.RESET_B(net23),
    .D(net869),
    .Q(\bp_core.ram_rdata[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _4047_ (.RESET_B(net22),
    .D(net417),
    .Q(\bp_core.ram_rdata[2] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _4048_ (.RESET_B(net21),
    .D(net389),
    .Q(\bp_core.ram_rdata[3] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _4049_ (.RESET_B(net20),
    .D(net224),
    .Q(\bp_core.ram_rdata[4] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _4050_ (.RESET_B(net19),
    .D(net267),
    .Q(\bp_core.ram_rdata[5] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _4051_ (.RESET_B(net18),
    .D(net228),
    .Q(\bp_core.ram_rdata[6] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _4052_ (.RESET_B(net17),
    .D(net332),
    .Q(\bp_core.ram_rdata[7] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _4053_ (.RESET_B(net16),
    .D(net9),
    .Q(\spi_ctrl.spi_miso_buf ),
    .CLK(net55));
 sg13g2_dfrbpq_1 _4054_ (.RESET_B(net774),
    .D(_0473_),
    .Q(\inter_bp.param_pending_reg[0] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _4055_ (.RESET_B(net824),
    .D(_0474_),
    .Q(\inter_bp.param_pending_reg[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _4056_ (.RESET_B(net811),
    .D(net491),
    .Q(\inter_bp.param_pending_reg[2] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4057_ (.RESET_B(net820),
    .D(net895),
    .Q(\inter_bp.param_pending_reg[3] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _4058_ (.RESET_B(net811),
    .D(net511),
    .Q(\inter_bp.param_pending_reg[4] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4059_ (.RESET_B(net825),
    .D(net554),
    .Q(\inter_bp.param_pending_reg[5] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4060_ (.RESET_B(net820),
    .D(_0479_),
    .Q(\inter_bp.param_pending_reg[6] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4061_ (.RESET_B(net825),
    .D(net852),
    .Q(\inter_bp.param_pending_reg[7] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4062_ (.RESET_B(net820),
    .D(net532),
    .Q(\inter_bp.param_pending_reg[8] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _4063_ (.RESET_B(net819),
    .D(net861),
    .Q(\inter_bp.param_pending_reg[9] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4064_ (.RESET_B(net818),
    .D(net843),
    .Q(\inter_bp.param_pending_reg[10] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _4065_ (.RESET_B(net818),
    .D(net524),
    .Q(\inter_bp.param_pending_reg[11] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4066_ (.RESET_B(net812),
    .D(net471),
    .Q(\inter_bp.param_pending_reg[12] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _4067_ (.RESET_B(net810),
    .D(_0486_),
    .Q(\inter_bp.param_pending_reg[13] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_1 _4068_ (.RESET_B(net810),
    .D(net901),
    .Q(\inter_bp.param_pending_reg[14] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4069_ (.RESET_B(net773),
    .D(net876),
    .Q(\inter_bp.param_pending_reg[15] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _4070_ (.RESET_B(net770),
    .D(net846),
    .Q(\inter_bp.param_pending_reg[16] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _4071_ (.RESET_B(net769),
    .D(net477),
    .Q(\inter_bp.param_pending_reg[17] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _4072_ (.RESET_B(net770),
    .D(_0491_),
    .Q(\inter_bp.param_pending_reg[18] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _4073_ (.RESET_B(net769),
    .D(net561),
    .Q(\inter_bp.param_pending_reg[19] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _4074_ (.RESET_B(net774),
    .D(net479),
    .Q(\inter_bp.param_pending_reg[20] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4075_ (.RESET_B(net760),
    .D(net489),
    .Q(\inter_bp.param_pending_reg[21] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _4076_ (.RESET_B(net807),
    .D(_0495_),
    .Q(\inter_bp.param_pending_reg[22] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4077_ (.RESET_B(net760),
    .D(net475),
    .Q(\inter_bp.param_pending_reg[23] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _4078_ (.RESET_B(net809),
    .D(net552),
    .Q(\inter_bp.param_pending_reg[24] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4079_ (.RESET_B(net759),
    .D(_0498_),
    .Q(\inter_bp.param_pending_reg[25] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _4080_ (.RESET_B(net809),
    .D(_0499_),
    .Q(\inter_bp.param_pending_reg[26] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_1 _4081_ (.RESET_B(net759),
    .D(_0500_),
    .Q(\inter_bp.param_pending_reg[27] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _4082_ (.RESET_B(net807),
    .D(net519),
    .Q(\inter_bp.param_pending_reg[28] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _4083_ (.RESET_B(net757),
    .D(net528),
    .Q(\inter_bp.param_pending_reg[29] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4084_ (.RESET_B(net773),
    .D(_0503_),
    .Q(\inter_bp.param_pending_reg[30] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _4085_ (.RESET_B(net761),
    .D(_0504_),
    .Q(\inter_bp.param_pending_reg[31] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _4086_ (.RESET_B(net774),
    .D(net465),
    .Q(\inter_bp.param_pending_reg[32] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _4087_ (.RESET_B(net761),
    .D(net469),
    .Q(\inter_bp.param_pending_reg[33] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4088_ (.RESET_B(net772),
    .D(net501),
    .Q(\inter_bp.param_pending_reg[34] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _4089_ (.RESET_B(net757),
    .D(net508),
    .Q(\inter_bp.param_pending_reg[35] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4090_ (.RESET_B(net771),
    .D(net467),
    .Q(\inter_bp.param_pending_reg[36] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _4091_ (.RESET_B(net758),
    .D(net547),
    .Q(\inter_bp.param_pending_reg[37] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _4092_ (.RESET_B(net761),
    .D(_0511_),
    .Q(\inter_bp.param_pending_reg[38] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _4093_ (.RESET_B(net765),
    .D(net544),
    .Q(\inter_bp.param_pending_reg[39] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4094_ (.RESET_B(net775),
    .D(net884),
    .Q(\inter_bp.param_pending_reg[40] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _4095_ (.RESET_B(net762),
    .D(_0514_),
    .Q(\inter_bp.param_pending_reg[41] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4096_ (.RESET_B(net767),
    .D(net874),
    .Q(\inter_bp.param_pending_reg[42] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4097_ (.RESET_B(net762),
    .D(net538),
    .Q(\inter_bp.param_pending_reg[43] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _4098_ (.RESET_B(net767),
    .D(net497),
    .Q(\inter_bp.param_pending_reg[44] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4099_ (.RESET_B(net764),
    .D(net559),
    .Q(\inter_bp.param_pending_reg[45] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _4100_ (.RESET_B(net764),
    .D(net503),
    .Q(\inter_bp.param_pending_reg[46] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _4101_ (.RESET_B(net764),
    .D(net542),
    .Q(\inter_bp.param_pending_reg[47] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_tiehi _4052__17 (.L_HI(net17));
 sg13g2_tiehi _4051__18 (.L_HI(net18));
 sg13g2_tiehi _4050__19 (.L_HI(net19));
 sg13g2_tiehi _4049__20 (.L_HI(net20));
 sg13g2_tiehi _4048__21 (.L_HI(net21));
 sg13g2_tiehi _4047__22 (.L_HI(net22));
 sg13g2_tiehi _4046__23 (.L_HI(net23));
 sg13g2_tiehi _4045__24 (.L_HI(net24));
 sg13g2_tiehi _4044__25 (.L_HI(net25));
 sg13g2_tiehi _4043__26 (.L_HI(net26));
 sg13g2_tiehi _4042__27 (.L_HI(net27));
 sg13g2_tiehi _4041__28 (.L_HI(net28));
 sg13g2_tiehi _4040__29 (.L_HI(net29));
 sg13g2_tiehi _4039__30 (.L_HI(net30));
 sg13g2_tiehi _4038__31 (.L_HI(net31));
 sg13g2_tiehi _4010__32 (.L_HI(net32));
 sg13g2_tiehi _4009__33 (.L_HI(net33));
 sg13g2_tiehi _4008__34 (.L_HI(net34));
 sg13g2_tiehi _4007__35 (.L_HI(net35));
 sg13g2_tiehi _4006__36 (.L_HI(net36));
 sg13g2_tiehi _4005__37 (.L_HI(net37));
 sg13g2_tiehi _4004__38 (.L_HI(net38));
 sg13g2_tiehi _4003__39 (.L_HI(net39));
 sg13g2_tiehi _4002__40 (.L_HI(net40));
 sg13g2_tiehi _4001__41 (.L_HI(net41));
 sg13g2_tiehi _4000__42 (.L_HI(net42));
 sg13g2_tiehi _3999__43 (.L_HI(net43));
 sg13g2_tiehi _3998__44 (.L_HI(net44));
 sg13g2_tiehi _3997__45 (.L_HI(net45));
 sg13g2_tiehi _3996__46 (.L_HI(net46));
 sg13g2_tiehi _3995__47 (.L_HI(net47));
 sg13g2_tiehi tt_um_swenson_cqs_48 (.L_HI(net48));
 sg13g2_tiehi tt_um_swenson_cqs_49 (.L_HI(net49));
 sg13g2_tiehi tt_um_swenson_cqs_50 (.L_HI(net50));
 sg13g2_tiehi tt_um_swenson_cqs_51 (.L_HI(net51));
 sg13g2_tiehi tt_um_swenson_cqs_52 (.L_HI(net52));
 sg13g2_tiehi tt_um_swenson_cqs_53 (.L_HI(net53));
 sg13g2_tiehi tt_um_swenson_cqs_54 (.L_HI(net54));
 sg13g2_inv_1 _2363__1 (.Y(net55),
    .A(clknet_1_1__leaf_clk));
 sg13g2_tielo tt_um_swenson_cqs_15 (.L_LO(net15));
 sg13g2_tiehi _4053__16 (.L_HI(net16));
 sg13g2_buf_2 _4143_ (.A(spi_cs),
    .X(uio_out[0]));
 sg13g2_buf_1 _4144_ (.A(net56),
    .X(uio_out[1]));
 sg13g2_buf_2 _4145_ (.A(\spi_ctrl.spi_mosi ),
    .X(uio_out[2]));
 sg13g2_buf_1 _4146_ (.A(\inter_bp.param_transmitting ),
    .X(uio_out[4]));
 sg13g2_buf_1 _4147_ (.A(\inter_bp.report_transmitting ),
    .X(uio_out[5]));
 sg13g2_buf_1 _4148_ (.A(\bp_core.busy_out ),
    .X(uo_out[0]));
 sg13g2_buf_1 _4149_ (.A(\bp_core.bp_report_valid_out ),
    .X(uo_out[2]));
 sg13g2_buf_8 fanout566 (.A(_1354_),
    .X(net566));
 sg13g2_buf_8 fanout567 (.A(net568),
    .X(net567));
 sg13g2_buf_8 fanout568 (.A(_1354_),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(net571),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(net571),
    .X(net570));
 sg13g2_buf_8 fanout571 (.A(_0974_),
    .X(net571));
 sg13g2_buf_8 fanout572 (.A(net573),
    .X(net572));
 sg13g2_buf_8 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_8 fanout574 (.A(net578),
    .X(net574));
 sg13g2_buf_8 fanout575 (.A(net578),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(net577),
    .X(net576));
 sg13g2_buf_1 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(_0971_),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(net580),
    .X(net579));
 sg13g2_buf_1 fanout580 (.A(_1744_),
    .X(net580));
 sg13g2_buf_8 fanout581 (.A(net583),
    .X(net581));
 sg13g2_buf_1 fanout582 (.A(net583),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(_1692_),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(net586),
    .X(net584));
 sg13g2_buf_1 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(_1584_),
    .X(net586));
 sg13g2_buf_8 fanout587 (.A(net588),
    .X(net587));
 sg13g2_buf_8 fanout588 (.A(net590),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_1103_),
    .X(net590));
 sg13g2_buf_8 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(net596),
    .X(net592));
 sg13g2_buf_8 fanout593 (.A(net594),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net596),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(net596),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(_1054_),
    .X(net596));
 sg13g2_buf_8 fanout597 (.A(net599),
    .X(net597));
 sg13g2_buf_1 fanout598 (.A(net599),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(_1054_),
    .X(net599));
 sg13g2_buf_8 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(net605),
    .X(net601));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_8 fanout603 (.A(net604),
    .X(net603));
 sg13g2_buf_8 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_1041_),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(net608),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_8 fanout608 (.A(_0953_),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(_0817_),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(_0817_),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_8 fanout613 (.A(_1691_),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(_1583_),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(net622),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(net621),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(net620),
    .X(net618));
 sg13g2_buf_1 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(net621),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(_1549_),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(_1260_),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(net626),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(net627),
    .X(net626));
 sg13g2_buf_8 fanout627 (.A(net629),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(_1156_),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(net631),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(_1156_),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(net633),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(_1048_),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(net636),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(net637),
    .X(net636));
 sg13g2_buf_8 fanout637 (.A(net641),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_8 fanout639 (.A(net641),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net641),
    .X(net640));
 sg13g2_buf_8 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(_1043_),
    .X(net642));
 sg13g2_buf_8 fanout643 (.A(net646),
    .X(net643));
 sg13g2_buf_8 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_8 fanout645 (.A(net646),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(net648),
    .X(net646));
 sg13g2_buf_8 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_8 fanout648 (.A(_0947_),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net651),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_0947_),
    .X(net650));
 sg13g2_buf_8 fanout651 (.A(_0947_),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(_0813_),
    .X(net652));
 sg13g2_buf_8 fanout653 (.A(_1333_),
    .X(net653));
 sg13g2_buf_8 fanout654 (.A(_1331_),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(_1329_),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(_1327_),
    .X(net656));
 sg13g2_buf_8 fanout657 (.A(_1325_),
    .X(net657));
 sg13g2_buf_8 fanout658 (.A(net659),
    .X(net658));
 sg13g2_buf_8 fanout659 (.A(_1047_),
    .X(net659));
 sg13g2_buf_8 fanout660 (.A(net661),
    .X(net660));
 sg13g2_buf_8 fanout661 (.A(_1047_),
    .X(net661));
 sg13g2_buf_8 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_8 fanout663 (.A(net664),
    .X(net663));
 sg13g2_buf_8 fanout664 (.A(net666),
    .X(net664));
 sg13g2_buf_8 fanout665 (.A(net666),
    .X(net665));
 sg13g2_buf_8 fanout666 (.A(net669),
    .X(net666));
 sg13g2_buf_8 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(net669),
    .X(net668));
 sg13g2_buf_8 fanout669 (.A(_1042_),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(_1042_),
    .X(net670));
 sg13g2_buf_8 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_1 fanout673 (.A(_1037_),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_1036_),
    .X(net675));
 sg13g2_buf_8 fanout676 (.A(net679),
    .X(net676));
 sg13g2_buf_8 fanout677 (.A(net679),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(net679),
    .X(net678));
 sg13g2_buf_8 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_8 fanout680 (.A(_0944_),
    .X(net680));
 sg13g2_buf_8 fanout681 (.A(net682),
    .X(net681));
 sg13g2_buf_8 fanout682 (.A(net683),
    .X(net682));
 sg13g2_buf_8 fanout683 (.A(_0944_),
    .X(net683));
 sg13g2_buf_8 fanout684 (.A(net687),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(net687),
    .X(net685));
 sg13g2_buf_1 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_8 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(_0843_),
    .X(net688));
 sg13g2_buf_8 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_8 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_8 fanout691 (.A(_0843_),
    .X(net691));
 sg13g2_buf_8 fanout692 (.A(net694),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(net694),
    .X(net693));
 sg13g2_buf_8 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_8 fanout695 (.A(_0842_),
    .X(net695));
 sg13g2_buf_8 fanout696 (.A(net697),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(net698),
    .X(net697));
 sg13g2_buf_8 fanout698 (.A(_0842_),
    .X(net698));
 sg13g2_buf_8 fanout699 (.A(net701),
    .X(net699));
 sg13g2_buf_8 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_8 fanout701 (.A(net705),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(net704),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(net704),
    .X(net703));
 sg13g2_buf_8 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_8 fanout705 (.A(net708),
    .X(net705));
 sg13g2_buf_8 fanout706 (.A(net708),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(net708),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(net715),
    .X(net708));
 sg13g2_buf_8 fanout709 (.A(net715),
    .X(net709));
 sg13g2_buf_2 fanout710 (.A(net715),
    .X(net710));
 sg13g2_buf_8 fanout711 (.A(net713),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(net713),
    .X(net712));
 sg13g2_buf_8 fanout713 (.A(net714),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(net715),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(_0841_),
    .X(net715));
 sg13g2_buf_8 fanout716 (.A(_0818_),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(net720),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(net719),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(_0547_),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(net727),
    .X(net721));
 sg13g2_buf_1 fanout722 (.A(net727),
    .X(net722));
 sg13g2_buf_8 fanout723 (.A(net725),
    .X(net723));
 sg13g2_buf_1 fanout724 (.A(net725),
    .X(net724));
 sg13g2_buf_8 fanout725 (.A(net727),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(net727),
    .X(net726));
 sg13g2_buf_8 fanout727 (.A(net1100),
    .X(net727));
 sg13g2_buf_8 fanout728 (.A(net730),
    .X(net728));
 sg13g2_buf_8 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(net737),
    .X(net730));
 sg13g2_buf_8 fanout731 (.A(net734),
    .X(net731));
 sg13g2_buf_1 fanout732 (.A(net734),
    .X(net732));
 sg13g2_buf_8 fanout733 (.A(net734),
    .X(net733));
 sg13g2_buf_8 fanout734 (.A(net737),
    .X(net734));
 sg13g2_buf_8 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_8 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_8 fanout737 (.A(\bp_core.params_module.state[2] ),
    .X(net737));
 sg13g2_buf_8 fanout738 (.A(net1180),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_1 fanout740 (.A(net743),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(net742),
    .X(net741));
 sg13g2_buf_8 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(\inter_bp.bp_report_valid_out ),
    .X(net743));
 sg13g2_buf_8 fanout744 (.A(net748),
    .X(net744));
 sg13g2_buf_1 fanout745 (.A(net748),
    .X(net745));
 sg13g2_buf_8 fanout746 (.A(net748),
    .X(net746));
 sg13g2_buf_1 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_8 fanout748 (.A(net458),
    .X(net748));
 sg13g2_buf_8 fanout749 (.A(net750),
    .X(net749));
 sg13g2_buf_8 fanout750 (.A(_0710_),
    .X(net750));
 sg13g2_buf_8 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(net753),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_8 fanout754 (.A(_0710_),
    .X(net754));
 sg13g2_buf_8 fanout755 (.A(_0709_),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(net3),
    .X(net756));
 sg13g2_buf_8 fanout757 (.A(net759),
    .X(net757));
 sg13g2_buf_8 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_8 fanout759 (.A(net768),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(net768),
    .X(net760));
 sg13g2_buf_8 fanout761 (.A(net768),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(net765),
    .X(net762));
 sg13g2_buf_8 fanout763 (.A(net765),
    .X(net763));
 sg13g2_buf_8 fanout764 (.A(net765),
    .X(net764));
 sg13g2_buf_8 fanout765 (.A(net768),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(net768),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(net768),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(net806),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net772),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(net772),
    .X(net770));
 sg13g2_buf_8 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(net779),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(net774),
    .X(net773));
 sg13g2_buf_8 fanout774 (.A(net779),
    .X(net774));
 sg13g2_buf_8 fanout775 (.A(net779),
    .X(net775));
 sg13g2_buf_1 fanout776 (.A(net779),
    .X(net776));
 sg13g2_buf_8 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_8 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(net806),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net784),
    .X(net780));
 sg13g2_buf_8 fanout781 (.A(net784),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(net784),
    .X(net782));
 sg13g2_buf_1 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(net795),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(net787),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net795),
    .X(net786));
 sg13g2_buf_8 fanout787 (.A(net795),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net791),
    .X(net788));
 sg13g2_buf_1 fanout789 (.A(net791),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_8 fanout791 (.A(net795),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(net794),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net794),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_8 fanout795 (.A(net806),
    .X(net795));
 sg13g2_buf_8 fanout796 (.A(net800),
    .X(net796));
 sg13g2_buf_8 fanout797 (.A(net800),
    .X(net797));
 sg13g2_buf_8 fanout798 (.A(net800),
    .X(net798));
 sg13g2_buf_8 fanout799 (.A(net800),
    .X(net799));
 sg13g2_buf_8 fanout800 (.A(net806),
    .X(net800));
 sg13g2_buf_8 fanout801 (.A(net805),
    .X(net801));
 sg13g2_buf_8 fanout802 (.A(net804),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(net804),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(net805),
    .X(net804));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805));
 sg13g2_buf_8 fanout806 (.A(net841),
    .X(net806));
 sg13g2_buf_8 fanout807 (.A(net809),
    .X(net807));
 sg13g2_buf_8 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_8 fanout809 (.A(net817),
    .X(net809));
 sg13g2_buf_8 fanout810 (.A(net812),
    .X(net810));
 sg13g2_buf_8 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_8 fanout812 (.A(net817),
    .X(net812));
 sg13g2_buf_8 fanout813 (.A(net814),
    .X(net813));
 sg13g2_buf_8 fanout814 (.A(net817),
    .X(net814));
 sg13g2_buf_8 fanout815 (.A(net816),
    .X(net815));
 sg13g2_buf_8 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_8 fanout817 (.A(net841),
    .X(net817));
 sg13g2_buf_8 fanout818 (.A(net819),
    .X(net818));
 sg13g2_buf_8 fanout819 (.A(net820),
    .X(net819));
 sg13g2_buf_8 fanout820 (.A(net825),
    .X(net820));
 sg13g2_buf_8 fanout821 (.A(net823),
    .X(net821));
 sg13g2_buf_8 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_8 fanout823 (.A(net825),
    .X(net823));
 sg13g2_buf_8 fanout824 (.A(net825),
    .X(net824));
 sg13g2_buf_8 fanout825 (.A(net841),
    .X(net825));
 sg13g2_buf_8 fanout826 (.A(net827),
    .X(net826));
 sg13g2_buf_8 fanout827 (.A(net829),
    .X(net827));
 sg13g2_buf_8 fanout828 (.A(net829),
    .X(net828));
 sg13g2_buf_8 fanout829 (.A(net840),
    .X(net829));
 sg13g2_buf_8 fanout830 (.A(net831),
    .X(net830));
 sg13g2_buf_8 fanout831 (.A(net832),
    .X(net831));
 sg13g2_buf_8 fanout832 (.A(net840),
    .X(net832));
 sg13g2_buf_8 fanout833 (.A(net837),
    .X(net833));
 sg13g2_buf_8 fanout834 (.A(net837),
    .X(net834));
 sg13g2_buf_8 fanout835 (.A(net836),
    .X(net835));
 sg13g2_buf_8 fanout836 (.A(net837),
    .X(net836));
 sg13g2_buf_8 fanout837 (.A(net840),
    .X(net837));
 sg13g2_buf_8 fanout838 (.A(net840),
    .X(net838));
 sg13g2_buf_8 fanout839 (.A(net840),
    .X(net839));
 sg13g2_buf_8 fanout840 (.A(net841),
    .X(net840));
 sg13g2_buf_8 fanout841 (.A(rst_n),
    .X(net841));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_2 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tielo tt_um_swenson_cqs_14 (.L_LO(net14));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_8 clkbuf_leaf_0_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_1_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_2_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_3_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_4_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_5_clk_regs (.A(clknet_4_1_0_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_6_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_7_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_8_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_9_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_10_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_11_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_12_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_13_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_14_clk_regs (.A(clknet_4_4_0_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_15_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_16_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_17_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_18_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_19_clk_regs (.A(clknet_4_5_0_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_20_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_21_clk_regs (.A(clknet_4_6_0_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_22_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_23_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_24_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_25_clk_regs (.A(clknet_4_7_0_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_26_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_27_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_28_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_29_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_30_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_31_clk_regs (.A(clknet_4_13_0_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_32_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_33_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_34_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_35_clk_regs (.A(clknet_4_15_0_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_36_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_37_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_38_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_39_clk_regs (.A(clknet_4_14_0_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_40_clk_regs (.A(clknet_4_12_0_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_41_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_42_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_43_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_44_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_45_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_46_clk_regs (.A(clknet_4_11_0_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_47_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_48_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_49_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_50_clk_regs (.A(clknet_4_10_0_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_51_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_52_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_53_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_54_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_55_clk_regs (.A(clknet_4_8_0_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_56_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_57_clk_regs (.A(clknet_4_9_0_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_58_clk_regs (.A(clknet_4_3_0_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_59_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_60_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_61_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_62_clk_regs (.A(clknet_4_2_0_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_63_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_64_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_65_clk_regs (.A(clknet_4_0_0_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_buf_8 clkload0 (.A(clknet_4_1_0_clk_regs));
 sg13g2_buf_8 clkload1 (.A(clknet_4_2_0_clk_regs));
 sg13g2_buf_8 clkload2 (.A(clknet_4_3_0_clk_regs));
 sg13g2_buf_8 clkload3 (.A(clknet_4_4_0_clk_regs));
 sg13g2_buf_8 clkload4 (.A(clknet_4_5_0_clk_regs));
 sg13g2_buf_8 clkload5 (.A(clknet_4_6_0_clk_regs));
 sg13g2_buf_8 clkload6 (.A(clknet_4_7_0_clk_regs));
 sg13g2_buf_8 clkload7 (.A(clknet_4_9_0_clk_regs));
 sg13g2_buf_8 clkload8 (.A(clknet_4_10_0_clk_regs));
 sg13g2_buf_8 clkload9 (.A(clknet_4_11_0_clk_regs));
 sg13g2_buf_8 clkload10 (.A(clknet_4_12_0_clk_regs));
 sg13g2_buf_8 clkload11 (.A(clknet_4_13_0_clk_regs));
 sg13g2_buf_8 clkload12 (.A(clknet_4_14_0_clk_regs));
 sg13g2_buf_8 clkload13 (.A(clknet_4_15_0_clk_regs));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_65_clk_regs));
 sg13g2_buf_8 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\bp_core.bp_report_valid_out ),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold2 (.A(\bp_core.bp_param_valid_out ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold3 (.A(\bp_core.params_module.state[3] ),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold4 (.A(\inter_bp.param_tx_shift_reg[15] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0223_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold6 (.A(\inter_bp.param_tx_shift_reg[27] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0235_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold8 (.A(\bp_core.bp_report_addr_out[10] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold9 (.A(_1281_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0273_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold11 (.A(\inter_bp.param_tx_shift_reg[23] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0233_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold13 (.A(\inter_bp.report_tx_shift_reg[5] ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold14 (.A(_1271_),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0268_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold16 (.A(\inter_bp.param_tx_shift_reg[16] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0226_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold18 (.A(\bp_core.bp_report_addr_out[8] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold19 (.A(_1277_),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold20 (.A(_0271_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0098_),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold22 (.A(\inter_bp.param_tx_shift_reg[19] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0229_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold24 (.A(\inter_bp.param_tx_shift_reg[14] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold25 (.A(_1185_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold26 (.A(\inter_bp.param_tx_shift_reg[32] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0242_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold28 (.A(\inter_bp.param_tx_shift_reg[21] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold29 (.A(_1199_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold30 (.A(\inter_bp.param_tx_shift_reg[12] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold31 (.A(_1181_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold32 (.A(\inter_bp.param_tx_shift_reg[17] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold33 (.A(_1187_),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold34 (.A(\inter_bp.param_tx_shift_reg[42] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0252_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold36 (.A(\inter_bp.param_tx_shift_reg[36] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0246_),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold38 (.A(\inter_bp.param_tx_shift_reg[43] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0251_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold40 (.A(\inter_bp.param_tx_shift_reg[38] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0248_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold42 (.A(\inter_bp.param_tx_shift_reg[30] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0240_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold44 (.A(\inter_bp.param_tx_shift_reg[7] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0217_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold46 (.A(\bp_addr_out[17] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold47 (.A(\inter_bp.param_tx_shift_reg[10] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold48 (.A(_1177_),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold49 (.A(\inter_bp.param_tx_shift_reg[11] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0221_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold51 (.A(\bp_core.ram_addr[8] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold52 (.A(_0408_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold53 (.A(\inter_bp.report_tx_shift_reg[13] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0276_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold55 (.A(\inter_bp.param_tx_shift_reg[34] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0244_),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold57 (.A(\bp_core.ram_addr[2] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold58 (.A(_0402_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold59 (.A(\bp_core.bp_report_addr_out[4] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold60 (.A(_1269_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0267_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold62 (.A(\inter_bp.report_tx_shift_reg[11] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0274_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold64 (.A(\bp_core.ram_addr[6] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0406_),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold66 (.A(\bp_core.ram_addr[7] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0407_),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold68 (.A(\bp_core.bp_report_addr_out[7] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold69 (.A(_1275_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0270_),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold71 (.A(\inter_bp.param_tx_shift_reg[33] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0243_),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold73 (.A(\inter_bp.param_tx_shift_reg[28] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold74 (.A(_1213_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold75 (.A(\bp_core.ram_addr[13] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0413_),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold77 (.A(\inter_bp.report_tx_shift_reg[16] ),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0279_),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold79 (.A(\inter_bp.param_tx_shift_reg[45] ),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold80 (.A(_1243_),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold81 (.A(\inter_bp.param_tx_shift_reg[20] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold82 (.A(_0230_),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold83 (.A(\inter_bp.param_tx_shift_reg[31] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0241_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold85 (.A(\bp_core.ram_addr[14] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0414_),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold87 (.A(\inter_bp.param_tx_shift_reg[40] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold88 (.A(_1237_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold89 (.A(\bp_core.bp_report_addr_out[9] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold90 (.A(_1279_),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold91 (.A(_0272_),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold92 (.A(\bp_core.ram_addr[1] ),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold93 (.A(_0401_),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold94 (.A(\inter_bp.report_tx_shift_reg[15] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0278_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold96 (.A(\bp_core.ram_addr[3] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0403_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold98 (.A(\bp_core.ram_addr[5] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0405_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold100 (.A(\bp_core.bp_report_addr_out[17] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold101 (.A(_1295_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold102 (.A(_0280_),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold103 (.A(\inter_bp.param_tx_shift_reg[0] ),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold104 (.A(_1155_),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0210_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold106 (.A(\inter_bp.param_tx_shift_reg[26] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold107 (.A(_0236_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold108 (.A(\bp_core.bp_report_addr_out[2] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold109 (.A(_1265_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold110 (.A(_0265_),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold111 (.A(\bp_core.params_module.params_ready ),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0012_),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold113 (.A(\bp_core.ram_addr[4] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0404_),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold115 (.A(\bp_core.ram_addr[15] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0415_),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold117 (.A(\bp_core.ram_addr[12] ),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0412_),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold119 (.A(\inter_bp.param_tx_shift_reg[39] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold120 (.A(_0247_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold121 (.A(\bp_core.ram_addr[10] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold122 (.A(_0410_),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold123 (.A(\inter_bp.param_tx_shift_reg[1] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold124 (.A(_1158_),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0211_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold126 (.A(\inter_bp.report_tx_shift_reg[0] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold127 (.A(_1261_),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold128 (.A(_0263_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold129 (.A(\inter_bp.report_tx_shift_reg[3] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold130 (.A(_1267_),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0266_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold132 (.A(\inter_bp.param_tx_shift_reg[37] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0245_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold134 (.A(\inter_bp.param_tx_shift_reg[18] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0228_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold136 (.A(\bp_core.ram_addr[9] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0409_),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold138 (.A(\bp_core.ram_addr[11] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0411_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold140 (.A(\inter_bp.param_tx_shift_reg[47] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold141 (.A(_1247_),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold142 (.A(\bp_core.params_module.state[1] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0329_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold144 (.A(\inter_bp.param_tx_shift_reg[29] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold145 (.A(_1211_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold146 (.A(\bp_core.bp_stride_out[9] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold147 (.A(\bp_core.bp_report_addr_out[12] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold148 (.A(_1285_),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0275_),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold150 (.A(\inter_bp.param_tx_shift_reg[24] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold151 (.A(_1205_),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold152 (.A(\bp_core.bp_report_addr_out[6] ),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold153 (.A(_1273_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0269_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold155 (.A(\inter_bp.param_tx_shift_reg[9] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold156 (.A(_1175_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold157 (.A(\inter_bp.param_tx_shift_reg[44] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold158 (.A(_0254_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold159 (.A(\bp_core.state[10] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold160 (.A(_0003_),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold161 (.A(\inter_bp.param_tx_shift_reg[5] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold162 (.A(_1167_),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold163 (.A(\bp_core.ram_addr[0] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0400_),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold165 (.A(\inter_bp.param_tx_shift_reg[22] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0232_),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold167 (.A(\bp_core.ram_wdata[4] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold168 (.A(_0469_),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold169 (.A(\spi_ctrl.bits_remaining[2] ),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold170 (.A(_0460_),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold171 (.A(\bp_core.ram_wdata[6] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0471_),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold173 (.A(\inter_bp.param_rx_counter[4] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0950_),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0094_),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold176 (.A(\inter_bp.param_tx_shift_reg[2] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0212_),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold178 (.A(\bp_core.bp_lambda_out[7] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold179 (.A(\spi_ctrl.addr[14] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold180 (.A(_1707_),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold181 (.A(_0441_),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold182 (.A(\spi_ctrl.addr[13] ),
    .X(net238));
 sg13g2_dlygate4sd3_1 hold183 (.A(_1706_),
    .X(net239));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0440_),
    .X(net240));
 sg13g2_dlygate4sd3_1 hold185 (.A(\bp_core.params_done ),
    .X(net241));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0701_),
    .X(net242));
 sg13g2_dlygate4sd3_1 hold187 (.A(\inter_bp.param_tx_shift_reg[3] ),
    .X(net243));
 sg13g2_dlygate4sd3_1 hold188 (.A(_0213_),
    .X(net244));
 sg13g2_dlygate4sd3_1 hold189 (.A(\inter_bp.param_tx_shift_reg[8] ),
    .X(net245));
 sg13g2_dlygate4sd3_1 hold190 (.A(_1173_),
    .X(net246));
 sg13g2_dlygate4sd3_1 hold191 (.A(\bp_core.bp_report_addr_out[1] ),
    .X(net247));
 sg13g2_dlygate4sd3_1 hold192 (.A(_1263_),
    .X(net248));
 sg13g2_dlygate4sd3_1 hold193 (.A(_0264_),
    .X(net249));
 sg13g2_dlygate4sd3_1 hold194 (.A(\bp_core.data_reg[0] ),
    .X(net250));
 sg13g2_dlygate4sd3_1 hold195 (.A(_0345_),
    .X(net251));
 sg13g2_dlygate4sd3_1 hold196 (.A(\spi_ctrl.addr[15] ),
    .X(net252));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0442_),
    .X(net253));
 sg13g2_dlygate4sd3_1 hold198 (.A(\inter_bp.bp_report_addr_out[13] ),
    .X(net254));
 sg13g2_dlygate4sd3_1 hold199 (.A(_1012_),
    .X(net255));
 sg13g2_dlygate4sd3_1 hold200 (.A(_0018_),
    .X(net256));
 sg13g2_dlygate4sd3_1 hold201 (.A(\inter_bp.report_shift_reg[0] ),
    .X(net257));
 sg13g2_dlygate4sd3_1 hold202 (.A(_1115_),
    .X(net258));
 sg13g2_dlygate4sd3_1 hold203 (.A(\inter_bp.report_tx_shift_reg[19] ),
    .X(net259));
 sg13g2_dlygate4sd3_1 hold204 (.A(_1298_),
    .X(net260));
 sg13g2_dlygate4sd3_1 hold205 (.A(\inter_bp.bp_report_addr_out[7] ),
    .X(net261));
 sg13g2_dlygate4sd3_1 hold206 (.A(_1000_),
    .X(net262));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0031_),
    .X(net263));
 sg13g2_dlygate4sd3_1 hold208 (.A(\spi_ctrl.addr[4] ),
    .X(net264));
 sg13g2_dlygate4sd3_1 hold209 (.A(_1697_),
    .X(net265));
 sg13g2_dlygate4sd3_1 hold210 (.A(\bp_core.ram_wdata[5] ),
    .X(net266));
 sg13g2_dlygate4sd3_1 hold211 (.A(_0470_),
    .X(net267));
 sg13g2_dlygate4sd3_1 hold212 (.A(\inter_bp.param_tx_shift_reg[6] ),
    .X(net268));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0216_),
    .X(net269));
 sg13g2_dlygate4sd3_1 hold214 (.A(\inter_bp.param_tx_counter[2] ),
    .X(net270));
 sg13g2_dlygate4sd3_1 hold215 (.A(_1139_),
    .X(net271));
 sg13g2_dlygate4sd3_1 hold216 (.A(_0202_),
    .X(net272));
 sg13g2_dlygate4sd3_1 hold217 (.A(\inter_bp.report_shift_reg[1] ),
    .X(net273));
 sg13g2_dlygate4sd3_1 hold218 (.A(_1116_),
    .X(net274));
 sg13g2_dlygate4sd3_1 hold219 (.A(\bp_core.bp_report_addr_out[14] ),
    .X(net275));
 sg13g2_dlygate4sd3_1 hold220 (.A(_1289_),
    .X(net276));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0277_),
    .X(net277));
 sg13g2_dlygate4sd3_1 hold222 (.A(\inter_bp.bp_report_addr_out[9] ),
    .X(net278));
 sg13g2_dlygate4sd3_1 hold223 (.A(_1004_),
    .X(net279));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0033_),
    .X(net280));
 sg13g2_dlygate4sd3_1 hold225 (.A(\inter_bp.bp_report_addr_out[5] ),
    .X(net281));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0996_),
    .X(net282));
 sg13g2_dlygate4sd3_1 hold227 (.A(_0029_),
    .X(net283));
 sg13g2_dlygate4sd3_1 hold228 (.A(\inter_bp.report_tx_shift_reg[18] ),
    .X(net284));
 sg13g2_dlygate4sd3_1 hold229 (.A(_1297_),
    .X(net285));
 sg13g2_dlygate4sd3_1 hold230 (.A(\inter_bp.bp_report_addr_out[15] ),
    .X(net286));
 sg13g2_dlygate4sd3_1 hold231 (.A(_0020_),
    .X(net287));
 sg13g2_dlygate4sd3_1 hold232 (.A(\inter_bp.param_rx_counter[0] ),
    .X(net288));
 sg13g2_dlygate4sd3_1 hold233 (.A(_0205_),
    .X(net289));
 sg13g2_dlygate4sd3_1 hold234 (.A(\bp_core.bp_param_output_data[1] ),
    .X(net290));
 sg13g2_dlygate4sd3_1 hold235 (.A(_0336_),
    .X(net291));
 sg13g2_dlygate4sd3_1 hold236 (.A(\bp_core.threshold_load_counter ),
    .X(net292));
 sg13g2_dlygate4sd3_1 hold237 (.A(_0010_),
    .X(net293));
 sg13g2_dlygate4sd3_1 hold238 (.A(\spi_ctrl.addr[9] ),
    .X(net294));
 sg13g2_dlygate4sd3_1 hold239 (.A(_1702_),
    .X(net295));
 sg13g2_dlygate4sd3_1 hold240 (.A(\bp_core.bp_param_output_data[3] ),
    .X(net296));
 sg13g2_dlygate4sd3_1 hold241 (.A(_0338_),
    .X(net297));
 sg13g2_dlygate4sd3_1 hold242 (.A(\inter_bp.bp_report_addr_out[8] ),
    .X(net298));
 sg13g2_dlygate4sd3_1 hold243 (.A(_1002_),
    .X(net299));
 sg13g2_dlygate4sd3_1 hold244 (.A(_0032_),
    .X(net300));
 sg13g2_dlygate4sd3_1 hold245 (.A(\inter_bp.param_tx_shift_reg[4] ),
    .X(net301));
 sg13g2_dlygate4sd3_1 hold246 (.A(_0214_),
    .X(net302));
 sg13g2_dlygate4sd3_1 hold247 (.A(\spi_ctrl.addr[2] ),
    .X(net303));
 sg13g2_dlygate4sd3_1 hold248 (.A(_1695_),
    .X(net304));
 sg13g2_dlygate4sd3_1 hold249 (.A(\spi_ctrl.addr[1] ),
    .X(net305));
 sg13g2_dlygate4sd3_1 hold250 (.A(_1694_),
    .X(net306));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0428_),
    .X(net307));
 sg13g2_dlygate4sd3_1 hold252 (.A(\inter_bp.report_rx_counter[0] ),
    .X(net308));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0154_),
    .X(net309));
 sg13g2_dlygate4sd3_1 hold254 (.A(\bp_core.state[3] ),
    .X(net310));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0397_),
    .X(net311));
 sg13g2_dlygate4sd3_1 hold256 (.A(\spi_ctrl.addr[10] ),
    .X(net312));
 sg13g2_dlygate4sd3_1 hold257 (.A(\spi_ctrl.addr[3] ),
    .X(net313));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0430_),
    .X(net314));
 sg13g2_dlygate4sd3_1 hold259 (.A(\spi_ctrl.addr[5] ),
    .X(net315));
 sg13g2_dlygate4sd3_1 hold260 (.A(\spi_ctrl.addr[7] ),
    .X(net316));
 sg13g2_dlygate4sd3_1 hold261 (.A(_1700_),
    .X(net317));
 sg13g2_dlygate4sd3_1 hold262 (.A(\inter_bp.param_rx_counter[3] ),
    .X(net318));
 sg13g2_dlygate4sd3_1 hold263 (.A(_1153_),
    .X(net319));
 sg13g2_dlygate4sd3_1 hold264 (.A(\inter_bp.param_tx_shift_reg[46] ),
    .X(net320));
 sg13g2_dlygate4sd3_1 hold265 (.A(_1248_),
    .X(net321));
 sg13g2_dlygate4sd3_1 hold266 (.A(\inter_bp.report_rx_counter[4] ),
    .X(net322));
 sg13g2_dlygate4sd3_1 hold267 (.A(_1113_),
    .X(net323));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0158_),
    .X(net324));
 sg13g2_dlygate4sd3_1 hold269 (.A(\inter_bp.report_tx_counter[2] ),
    .X(net325));
 sg13g2_dlygate4sd3_1 hold270 (.A(_1254_),
    .X(net326));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0260_),
    .X(net327));
 sg13g2_dlygate4sd3_1 hold272 (.A(\inter_bp.bp_report_addr_out[6] ),
    .X(net328));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0998_),
    .X(net329));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0030_),
    .X(net330));
 sg13g2_dlygate4sd3_1 hold275 (.A(\bp_core.ram_rdata[6] ),
    .X(net331));
 sg13g2_dlygate4sd3_1 hold276 (.A(_0472_),
    .X(net332));
 sg13g2_dlygate4sd3_1 hold277 (.A(\bp_core.addr_reg[2] ),
    .X(net333));
 sg13g2_dlygate4sd3_1 hold278 (.A(_0986_),
    .X(net334));
 sg13g2_dlygate4sd3_1 hold279 (.A(\bp_core.threshold_reg[0] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold280 (.A(\inter_bp.bp_report_addr_out[10] ),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold281 (.A(_1006_),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold282 (.A(_0015_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold283 (.A(\spi_ctrl.addr[11] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0438_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold285 (.A(\bp_core.data_reg[6] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold286 (.A(\bp_core.bp_report_addr_out[16] ),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0021_),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold288 (.A(\bp_core.bp_report_addr_out[0] ),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0014_),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold290 (.A(\spi_ctrl.addr[6] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold291 (.A(\bp_core.data_reg[4] ),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0349_),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold293 (.A(\inter_bp.param_shift_reg[41] ),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0065_),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold295 (.A(\bp_core.status_out[3] ),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold296 (.A(_0041_),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold297 (.A(\bp_core.status_out[0] ),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold298 (.A(_0038_),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold299 (.A(\bp_core.ram_wdata[7] ),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0399_),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold301 (.A(\bp_core.ram_wdata[0] ),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0392_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0102_),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold304 (.A(\bp_core.data_reg[5] ),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold305 (.A(_0350_),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold306 (.A(\spi_ctrl.addr[8] ),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold307 (.A(\bp_core.ram_rdata[4] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold308 (.A(\bp_core.data_reg[2] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold309 (.A(_0347_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold310 (.A(\spi_ctrl.addr[0] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold311 (.A(_1693_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold312 (.A(\bp_core.init_counter[15] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold313 (.A(_1617_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0389_),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold315 (.A(\bp_core.addr_reg[4] ),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0995_),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold317 (.A(\bp_core.data_reg[3] ),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold318 (.A(\inter_bp.report_shift_reg[17] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold319 (.A(_1132_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold320 (.A(\inter_bp.report_shift_reg[13] ),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold321 (.A(_1128_),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold322 (.A(\spi_ctrl.addr[12] ),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0439_),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold324 (.A(\spi_ctrl.bits_remaining[0] ),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0458_),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold326 (.A(\bp_core.status_out[1] ),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0039_),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold328 (.A(\bp_core.data_reg[7] ),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0352_),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold330 (.A(\inter_bp.report_shift_reg[8] ),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold331 (.A(_1123_),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold332 (.A(\bp_core.ram_rdata[3] ),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold333 (.A(_0468_),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold334 (.A(\inter_bp.param_tx_shift_reg[41] ),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0249_),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold336 (.A(\inter_bp.bp_report_addr_out[12] ),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold337 (.A(_0017_),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold338 (.A(\bp_core.status_out[2] ),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold339 (.A(\inter_bp.param_rx_counter[2] ),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0949_),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold341 (.A(\inter_bp.param_shift_reg[0] ),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0044_),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold343 (.A(\bp_core.bp_lambda_out[6] ),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold344 (.A(_1541_),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold345 (.A(\inter_bp.bp_report_addr_out[1] ),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0180_),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold347 (.A(\inter_bp.report_shift_reg[14] ),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold348 (.A(_1129_),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold349 (.A(\bp_core.status_out[4] ),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold350 (.A(\spi_ctrl.writing ),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0464_),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold352 (.A(\inter_bp.param_shift_reg[1] ),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold353 (.A(_1056_),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold354 (.A(\inter_bp.report_shift_reg[2] ),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold355 (.A(_1117_),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold356 (.A(\bp_core.data_reg[1] ),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold357 (.A(_0346_),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold358 (.A(\inter_bp.bp_report_addr_out[14] ),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold359 (.A(_0019_),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold360 (.A(\bp_core.ram_rdata[2] ),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold361 (.A(_0467_),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold362 (.A(\inter_bp.report_shift_reg[9] ),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold363 (.A(_1124_),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0100_),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold365 (.A(_1319_),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold366 (.A(_0290_),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0099_),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold368 (.A(_1318_),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0289_),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold370 (.A(\inter_bp.report_shift_reg[6] ),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold371 (.A(\inter_bp.param_shift_reg[31] ),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0075_),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold373 (.A(\inter_bp.param_shift_reg[25] ),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold374 (.A(_1080_),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold375 (.A(\inter_bp.report_shift_reg[10] ),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold376 (.A(_1125_),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold377 (.A(\bp_addr_in[0] ),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0453_),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold379 (.A(\inter_bp.report_shift_reg[15] ),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0194_),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold381 (.A(\inter_bp.report_shift_reg[16] ),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold382 (.A(_1131_),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold383 (.A(\inter_bp.bp_report_addr_out[3] ),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0182_),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold385 (.A(\bp_core.ram_wdata[3] ),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold386 (.A(\inter_bp.bp_report_addr_out[11] ),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0016_),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold388 (.A(\inter_bp.param_shift_reg[22] ),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold389 (.A(_1077_),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold390 (.A(\bp_core.addr_reg[1] ),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold391 (.A(\inter_bp.report_shift_reg[11] ),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold392 (.A(\inter_bp.report_rx_counter[3] ),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold393 (.A(_1112_),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0157_),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold395 (.A(\inter_bp.param_shift_reg[27] ),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold396 (.A(_1082_),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold397 (.A(\bp_core.threshold_reg[1] ),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold398 (.A(\bp_core.busy_out ),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold399 (.A(_0373_),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold400 (.A(\bp_core.ram_wdata[1] ),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0393_),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold402 (.A(\inter_bp.report_rx_done ),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold403 (.A(\bp_core.bp_param_output_data[0] ),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0335_),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold405 (.A(\inter_bp.from_left_report_valid_prev ),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold406 (.A(\inter_bp.param_shift_reg[38] ),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold407 (.A(_1093_),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold408 (.A(\inter_bp.param_pending_reg[32] ),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0505_),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold410 (.A(\inter_bp.param_pending_reg[36] ),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0509_),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold412 (.A(\inter_bp.param_pending_reg[33] ),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0506_),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold414 (.A(\inter_bp.param_pending_reg[12] ),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0485_),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold416 (.A(\inter_bp.param_pending_reg[27] ),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold417 (.A(\inter_bp.param_pending_reg[25] ),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold418 (.A(\inter_bp.param_pending_reg[23] ),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold419 (.A(_0496_),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold420 (.A(\inter_bp.param_pending_reg[17] ),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold421 (.A(_0490_),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold422 (.A(\inter_bp.param_pending_reg[20] ),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold423 (.A(_0493_),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold424 (.A(\bp_core.init_counter[9] ),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0383_),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold426 (.A(\bp_core.addr_reg[18] ),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold427 (.A(_0371_),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold428 (.A(\inter_bp.param_shift_reg[13] ),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold429 (.A(_1068_),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold430 (.A(\inter_bp.report_shift_reg[3] ),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold431 (.A(_1118_),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold432 (.A(\inter_bp.param_pending_reg[21] ),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0494_),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold434 (.A(\inter_bp.param_pending_reg[2] ),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0475_),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold436 (.A(\bp_core.ram_wdata[2] ),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold437 (.A(\inter_bp.param_shift_reg[6] ),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold438 (.A(_1061_),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold439 (.A(\inter_bp.param_pending_reg[0] ),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold440 (.A(\inter_bp.param_pending_reg[44] ),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0517_),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold442 (.A(\inter_bp.param_shift_reg[26] ),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold443 (.A(_1081_),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold444 (.A(\inter_bp.param_pending_reg[34] ),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold445 (.A(_0507_),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold446 (.A(\inter_bp.param_pending_reg[46] ),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0519_),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold448 (.A(\inter_bp.report_shift_reg[5] ),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold449 (.A(\bp_core.state[11] ),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0832_),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold451 (.A(\inter_bp.param_pending_reg[35] ),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0508_),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold453 (.A(\inter_bp.param_pending_reg[22] ),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold454 (.A(\inter_bp.param_pending_reg[4] ),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold455 (.A(_0477_),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold456 (.A(\bp_core.bp_stride_in[11] ),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0302_),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold458 (.A(\inter_bp.param_pending_reg[6] ),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold459 (.A(\inter_bp.param_shift_reg[36] ),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold460 (.A(\bp_core.threshold_reg[2] ),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0418_),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold462 (.A(\inter_bp.param_pending_reg[28] ),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0501_),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold464 (.A(\inter_bp.param_tx_counter[0] ),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold465 (.A(_1135_),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0200_),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold467 (.A(\inter_bp.param_pending_reg[11] ),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0484_),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold469 (.A(\inter_bp.param_shift_reg[28] ),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold470 (.A(_1083_),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold471 (.A(\inter_bp.param_pending_reg[29] ),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0502_),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold473 (.A(\inter_bp.param_shift_reg[17] ),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold474 (.A(_1072_),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold475 (.A(\inter_bp.param_pending_reg[8] ),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0481_),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold477 (.A(\inter_bp.param_shift_reg[11] ),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold478 (.A(\inter_bp.param_shift_reg[4] ),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold479 (.A(\inter_bp.bp_report_addr_out[0] ),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold480 (.A(\inter_bp.param_pending_reg[31] ),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold481 (.A(\inter_bp.param_pending_reg[43] ),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold482 (.A(_0516_),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold483 (.A(\inter_bp.report_shift_reg[7] ),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0101_),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold485 (.A(\inter_bp.param_pending_reg[47] ),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0520_),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold487 (.A(\inter_bp.param_pending_reg[39] ),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0512_),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold489 (.A(\inter_bp.param_pending_reg[38] ),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold490 (.A(\inter_bp.param_pending_reg[37] ),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0510_),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold492 (.A(\bp_core.bp_stride_in[5] ),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold493 (.A(\spi_ctrl.bits_remaining[1] ),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold494 (.A(_1738_),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold495 (.A(\inter_bp.param_pending_reg[24] ),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold496 (.A(_0497_),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold497 (.A(\inter_bp.param_pending_reg[5] ),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold498 (.A(_0478_),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold499 (.A(\inter_bp.report_tx_counter[0] ),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold500 (.A(_1250_),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0258_),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold502 (.A(\inter_bp.param_pending_reg[45] ),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0518_),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold504 (.A(\inter_bp.param_pending_reg[19] ),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0492_),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold506 (.A(\inter_bp.param_pending_reg[1] ),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold507 (.A(\bp_core.bp_stride_in[2] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0085_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold509 (.A(\inter_bp.param_pending_reg[13] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold510 (.A(\inter_bp.param_pending_reg[10] ),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0483_),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold512 (.A(\bp_core.bp_stride_in[16] ),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold513 (.A(\inter_bp.param_pending_reg[16] ),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0489_),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold515 (.A(\bp_core.bp_report_addr_out[3] ),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0027_),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold517 (.A(\inter_bp.param_shift_reg[30] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold518 (.A(_1085_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold519 (.A(\inter_bp.param_pending_reg[7] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0480_),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold521 (.A(\inter_bp.param_shift_reg[12] ),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold522 (.A(_1067_),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold523 (.A(\inter_bp.report_receiving ),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold524 (.A(\inter_bp.param_shift_reg[21] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold525 (.A(_0084_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold526 (.A(\inter_bp.report_shift_reg[4] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold527 (.A(\inter_bp.param_pending_reg[30] ),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold528 (.A(\inter_bp.param_pending_reg[9] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0482_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold530 (.A(\inter_bp.param_shift_reg[43] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0067_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold532 (.A(\bp_core.initialized ),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0421_),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold534 (.A(\inter_bp.param_shift_reg[32] ),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold535 (.A(_1087_),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold536 (.A(\bp_core.ram_rdata[1] ),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold537 (.A(_0466_),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold538 (.A(\inter_bp.param_pending_reg[26] ),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold539 (.A(_0899_),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0089_),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold541 (.A(\inter_bp.param_pending_reg[42] ),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0515_),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold543 (.A(\inter_bp.param_pending_reg[15] ),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold544 (.A(_0488_),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold545 (.A(\bp_core.params_addr[18] ),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold546 (.A(_0343_),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold547 (.A(\bp_core.ram_we ),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold548 (.A(_0391_),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold549 (.A(\inter_bp.param_shift_reg[24] ),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold550 (.A(\inter_bp.param_shift_reg[19] ),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold551 (.A(\inter_bp.param_pending_reg[40] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold552 (.A(_0513_),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold553 (.A(\inter_bp.param_pending_reg[41] ),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold554 (.A(\inter_bp.param_shift_reg[45] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold555 (.A(_0069_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold556 (.A(\inter_bp.param_shift_reg[18] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold557 (.A(_1073_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold558 (.A(\inter_bp.param_rx_done ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold559 (.A(\inter_bp.param_shift_reg[10] ),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold560 (.A(\inter_bp.bp_report_addr_out[4] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold561 (.A(\inter_bp.report_shift_reg[12] ),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold562 (.A(\inter_bp.param_pending_reg[3] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold563 (.A(_0476_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold564 (.A(\inter_bp.param_pending_reg[18] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold565 (.A(_0883_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold566 (.A(\inter_bp.param_shift_reg[33] ),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold567 (.A(_1088_),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold568 (.A(\inter_bp.param_pending_reg[14] ),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold569 (.A(_0487_),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold570 (.A(\bp_addr_in[1] ),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold571 (.A(\bp_core.bp_stride_in[4] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold572 (.A(\inter_bp.param_shift_reg[3] ),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold573 (.A(_1058_),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold574 (.A(\bp_core.bp_stride_in[10] ),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold575 (.A(\inter_bp.param_shift_reg[7] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold576 (.A(_1062_),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold577 (.A(\bp_addr_in[6] ),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold578 (.A(\inter_bp.param_shift_reg[47] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold579 (.A(\bp_addr_in[17] ),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold580 (.A(\inter_bp.param_shift_reg[35] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold581 (.A(_1090_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold582 (.A(\inter_bp.param_tx_counter[3] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold583 (.A(_1141_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold584 (.A(_0203_),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold585 (.A(\inter_bp.param_shift_reg[44] ),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold586 (.A(_1099_),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold587 (.A(\bp_core.bp_lambda_in[7] ),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold588 (.A(\inter_bp.param_shift_reg[9] ),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold589 (.A(\inter_bp.param_shift_reg[34] ),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold590 (.A(\bp_core.params_module.start_load ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold591 (.A(_0830_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold592 (.A(_1800_[0]),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold593 (.A(\bp_core.bp_stride_in[12] ),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold594 (.A(\inter_bp.param_shift_reg[2] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold595 (.A(\inter_bp.param_shift_reg[5] ),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold596 (.A(\bp_core.bp_stride_in[18] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold597 (.A(\bp_core.state[5] ),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold598 (.A(_0004_),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold599 (.A(\bp_addr_in[4] ),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold600 (.A(\bp_core.addr_reg[17] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold601 (.A(_0022_),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold602 (.A(\inter_bp.param_shift_reg[8] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold603 (.A(\inter_bp.param_shift_reg[23] ),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold604 (.A(\bp_addr_in[11] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold605 (.A(\bp_addr_in[12] ),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold606 (.A(\bp_core.bp_lambda_in[4] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold607 (.A(\inter_bp.param_shift_reg[39] ),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold608 (.A(\inter_bp.param_shift_reg[16] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold609 (.A(_0051_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold610 (.A(\inter_bp.param_shift_reg[20] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold611 (.A(\bp_core.state[4] ),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold612 (.A(_0008_),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold613 (.A(\inter_bp.param_shift_reg[40] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold614 (.A(_0064_),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold615 (.A(\bp_core.bp_stride_in[8] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold616 (.A(\inter_bp.param_shift_reg[37] ),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold617 (.A(\bp_core.bp_stride_in[14] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold618 (.A(\bp_addr_in[5] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold619 (.A(\bp_core.bp_stride_in[7] ),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold620 (.A(\bp_core.bp_param_output_data[2] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold621 (.A(_0337_),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold622 (.A(\bp_core.bp_stride_in[13] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold623 (.A(\bp_core.params_addr[2] ),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold624 (.A(_0455_),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold625 (.A(\bp_core.params_addr[9] ),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold626 (.A(_0452_),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold627 (.A(\bp_core.bp_param_output_data[4] ),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold628 (.A(_0339_),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold629 (.A(\inter_bp.param_shift_reg[29] ),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold630 (.A(_0092_),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold631 (.A(\bp_core.state[2] ),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold632 (.A(_0006_),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold633 (.A(\inter_bp.param_rx_counter[1] ),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold634 (.A(\bp_addr_in[10] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold635 (.A(\bp_core.bp_stride_in[19] ),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold636 (.A(\inter_bp.param_pending ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold637 (.A(_0093_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold638 (.A(\bp_addr_in[13] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold639 (.A(\inter_bp.param_shift_reg[42] ),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold640 (.A(\bp_core.bp_report_addr_out[18] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold641 (.A(_0023_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold642 (.A(\bp_core.params_addr[16] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold643 (.A(_0341_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold644 (.A(\bp_core.params_addr[5] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold645 (.A(\bp_core.bp_stride_in[15] ),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold646 (.A(\bp_core.bp_lambda_in[2] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold647 (.A(\bp_core.params_addr[11] ),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold648 (.A(\inter_bp.bp_report_addr_out[19] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold649 (.A(_0198_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold650 (.A(\bp_core.bp_stride_in[3] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold651 (.A(\bp_addr_in[9] ),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold652 (.A(\bp_addr_in[19] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold653 (.A(\bp_core.params_addr[17] ),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold654 (.A(\bp_core.params_addr[4] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold655 (.A(_0457_),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold656 (.A(\bp_core.params_addr[10] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold657 (.A(\bp_core.params_addr[6] ),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold658 (.A(\inter_bp.bp_report_addr_out[17] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold659 (.A(\bp_addr_in[2] ),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold660 (.A(\inter_bp.param_shift_reg[46] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold661 (.A(_0070_),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold662 (.A(\bp_addr_in[3] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold663 (.A(\bp_addr_in[8] ),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold664 (.A(\inter_bp.param_receiving ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold665 (.A(_0287_),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold666 (.A(\inter_bp.bp_report_addr_out[2] ),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold667 (.A(\bp_addr_in[7] ),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold668 (.A(\bp_core.threshold_reg[5] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold669 (.A(\inter_bp.report_shift_reg[18] ),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold670 (.A(_0197_),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold671 (.A(\inter_bp.bp_report_addr_out[16] ),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold672 (.A(\inter_bp.param_shift_reg[14] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold673 (.A(\inter_bp.param_shift_reg[15] ),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold674 (.A(\bp_core.bp_stride_in[17] ),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold675 (.A(\inter_bp.report_tx_counter[3] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold676 (.A(_1256_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold677 (.A(_0261_),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold678 (.A(\bp_core.params_addr[8] ),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold679 (.A(\bp_core.params_addr[12] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold680 (.A(\bp_core.init_counter[10] ),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold681 (.A(_1607_),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold682 (.A(\bp_core.bp_stride_in[0] ),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold683 (.A(_0073_),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold684 (.A(\bp_core.params_addr[1] ),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold685 (.A(_0454_),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold686 (.A(\bp_addr_in[14] ),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold687 (.A(\bp_addr_out[16] ),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold688 (.A(_0325_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold689 (.A(\bp_core.init_counter[7] ),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold690 (.A(_1600_),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold691 (.A(\bp_addr_out[2] ),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold692 (.A(\bp_core.params_addr[15] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold693 (.A(_0340_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold694 (.A(\bp_core.params_forward ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold695 (.A(\inter_bp.report_shift_reg[19] ),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold696 (.A(\bp_core.threshold_reg[4] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold697 (.A(\bp_core.params_addr[7] ),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold698 (.A(\bp_core.init_counter[6] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold699 (.A(_1598_),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold700 (.A(\bp_addr_out[1] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold701 (.A(\bp_core.init_counter[3] ),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold702 (.A(_1591_),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold703 (.A(\bp_core.params_addr[3] ),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold704 (.A(\bp_core.params_addr[19] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold705 (.A(\bp_core.params_addr[13] ),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold706 (.A(\bp_addr_out[19] ),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold707 (.A(_0328_),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold708 (.A(\inter_bp.report_tx_counter[4] ),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold709 (.A(_1259_),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold710 (.A(\bp_core.state[9] ),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold711 (.A(\bp_addr_in[15] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold712 (.A(\bp_core.init_counter[4] ),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold713 (.A(_1593_),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold714 (.A(\bp_core.params_addr[14] ),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold715 (.A(\bp_addr_out[15] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold716 (.A(_0324_),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold717 (.A(\bp_core.init_counter[13] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold718 (.A(_1614_),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold719 (.A(\bp_core.init_counter[14] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold720 (.A(_1616_),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold721 (.A(\bp_core.init_counter[2] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold722 (.A(_1589_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold723 (.A(\bp_core.addr_reg[9] ),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold724 (.A(\bp_addr_out[4] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold725 (.A(\bp_core.init_counter[8] ),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold726 (.A(_1602_),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold727 (.A(\bp_addr_out[0] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold728 (.A(_0309_),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold729 (.A(\bp_core.addr_reg[10] ),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold730 (.A(_0363_),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold731 (.A(\inter_bp.report_rx_counter[2] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold732 (.A(_0955_),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold733 (.A(\bp_addr_out[18] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold734 (.A(_0327_),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold735 (.A(\inter_bp.param_tx_counter[4] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold736 (.A(_1046_),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold737 (.A(_0095_),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold738 (.A(\bp_core.ram_rdata[0] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold739 (.A(_0465_),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold740 (.A(\bp_addr_out[10] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold741 (.A(\bp_addr_out[8] ),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold742 (.A(_0317_),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold743 (.A(\bp_core.init_counter[12] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold744 (.A(_1612_),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold745 (.A(\bp_addr_out[12] ),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold746 (.A(_0321_),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold747 (.A(\inter_bp.report_tx_counter[1] ),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold748 (.A(_1253_),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold749 (.A(\bp_addr_out[11] ),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold750 (.A(_0320_),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold751 (.A(\inter_bp.serialize_param_valid_prev ),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold752 (.A(\inter_bp.param_tx_counter[1] ),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold753 (.A(_1138_),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold754 (.A(\inter_bp.report_rx_counter[1] ),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold755 (.A(\bp_addr_out[13] ),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold756 (.A(_0322_),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold757 (.A(\bp_addr_out[7] ),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold758 (.A(_0316_),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold759 (.A(\bp_addr_out[9] ),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold760 (.A(\bp_core.addr_reg[19] ),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold761 (.A(\bp_core.bp_stride_out[17] ),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold762 (.A(\bp_core.init_counter[11] ),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold763 (.A(\bp_addr_out[5] ),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold764 (.A(_0314_),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold765 (.A(\bp_core.params_module.counter[3] ),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold766 (.A(_0719_),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold767 (.A(_0833_),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold768 (.A(\bp_core.state[7] ),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold769 (.A(_1371_),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold770 (.A(\bp_addr_out[3] ),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold771 (.A(_0312_),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold772 (.A(\bp_addr_out[14] ),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold773 (.A(_0323_),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold774 (.A(\bp_core.addr_reg[3] ),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold775 (.A(_0356_),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold776 (.A(\bp_core.init_counter[1] ),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold777 (.A(_1586_),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold778 (.A(\bp_core.state[6] ),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold779 (.A(\bp_core.init_counter[5] ),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold780 (.A(\bp_addr_out[6] ),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold781 (.A(_0315_),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold782 (.A(\inter_bp.report_transmitting ),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold783 (.A(\bp_core.addr_reg[11] ),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold784 (.A(_0364_),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold785 (.A(\bp_core.bp_stride_out[15] ),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold786 (.A(\bp_core.addr_reg[8] ),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold787 (.A(\bp_core.addr_reg[6] ),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold788 (.A(\bp_core.addr_reg[16] ),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold789 (.A(\bp_core.bp_report_addr_out[19] ),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold790 (.A(_1032_),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold791 (.A(\bp_core.bp_lambda_in[1] ),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold792 (.A(_0297_),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold793 (.A(\bp_core.bp_param_ack_out ),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold794 (.A(\bp_core.addr_reg[13] ),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold795 (.A(\bp_core.addr_reg[12] ),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold796 (.A(\bp_core.bp_stride_out[10] ),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold797 (.A(\bp_core.addr_reg[15] ),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold798 (.A(\bp_core.addr_reg[7] ),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold799 (.A(_0360_),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold800 (.A(\bp_core.state[8] ),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold801 (.A(\bp_core.addr_reg[14] ),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold802 (.A(\bp_core.addr_reg[0] ),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold803 (.A(_0353_),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold804 (.A(\bp_core.bp_stride_out[19] ),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold805 (.A(\bp_core.bp_stride_out[0] ),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold806 (.A(\bp_core.bp_stride_out[1] ),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold807 (.A(_0423_),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold808 (.A(\bp_core.bp_param_valid_in ),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold809 (.A(\bp_core.addr_reg[2] ),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold810 (.A(_0737_),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold811 (.A(\bp_core.bp_lambda_in[6] ),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold812 (.A(\bp_core.bp_stride_out[14] ),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold813 (.A(\bp_core.bp_stride_out[16] ),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold814 (.A(\bp_core.init_counter[0] ),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold815 (.A(\bp_core.params_module.counter[2] ),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold816 (.A(_1312_),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold817 (.A(\bp_core.params_module.counter[0] ),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold818 (.A(\bp_core.bp_stride_out[18] ),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold819 (.A(\bp_core.bp_stride_out[2] ),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold820 (.A(\spi_ctrl.fsm_state[1] ),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold821 (.A(_1743_),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold822 (.A(\bp_core.bp_stride_out[5] ),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold823 (.A(\bp_core.params_module.counter[0] ),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold824 (.A(\bp_core.bp_stride_out[3] ),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold825 (.A(\bp_core.addr_reg[5] ),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold826 (.A(\bp_core.bp_lambda_out[5] ),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold827 (.A(_0306_),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold828 (.A(\bp_core.bp_lambda_out[0] ),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold829 (.A(_0296_),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold830 (.A(\bp_core.bp_stride_out[12] ),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold831 (.A(\bp_core.addr_reg[1] ),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold832 (.A(\bp_core.bp_stride_out[7] ),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold833 (.A(\bp_core.bp_stride_in[9] ),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold834 (.A(\bp_core.state[1] ),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold835 (.A(\bp_core.bp_stride_out[13] ),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold836 (.A(\bp_core.bp_lambda_out[4] ),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold837 (.A(\spi_ctrl.bits_remaining[3] ),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold838 (.A(_1741_),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold839 (.A(\bp_core.bp_stride_out[8] ),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold840 (.A(\bp_core.bp_lambda_out[2] ),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold841 (.A(\spi_ctrl.fsm_state[0] ),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold842 (.A(_1742_),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold843 (.A(\bp_core.bp_stride_out[6] ),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold844 (.A(_0292_),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold845 (.A(\bp_core.bp_lambda_out[3] ),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold846 (.A(_0299_),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold847 (.A(\bp_core.bp_stride_out[4] ),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold848 (.A(\bp_core.params_module.counter[1] ),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold849 (.A(\inter_bp.param_rx_counter[1] ),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold850 (.A(\inter_bp.param_tx_counter[1] ),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold851 (.A(\bp_core.bp_stride_out[4] ),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold852 (.A(\bp_core.bp_stride_out[13] ),
    .X(net1184));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_fill_1 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_fill_1 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_decap_8 FILLER_2_427 ();
 sg13g2_decap_8 FILLER_2_434 ();
 sg13g2_decap_8 FILLER_2_441 ();
 sg13g2_decap_8 FILLER_2_448 ();
 sg13g2_decap_8 FILLER_2_455 ();
 sg13g2_decap_8 FILLER_2_462 ();
 sg13g2_decap_8 FILLER_2_469 ();
 sg13g2_decap_8 FILLER_2_476 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_8 FILLER_2_497 ();
 sg13g2_decap_8 FILLER_2_504 ();
 sg13g2_decap_8 FILLER_2_511 ();
 sg13g2_decap_8 FILLER_2_518 ();
 sg13g2_decap_8 FILLER_2_525 ();
 sg13g2_decap_8 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_539 ();
 sg13g2_decap_8 FILLER_2_546 ();
 sg13g2_decap_8 FILLER_2_553 ();
 sg13g2_decap_8 FILLER_2_560 ();
 sg13g2_decap_8 FILLER_2_567 ();
 sg13g2_decap_8 FILLER_2_574 ();
 sg13g2_decap_8 FILLER_2_581 ();
 sg13g2_decap_8 FILLER_2_588 ();
 sg13g2_decap_8 FILLER_2_595 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_8 FILLER_2_609 ();
 sg13g2_decap_8 FILLER_2_616 ();
 sg13g2_decap_8 FILLER_2_623 ();
 sg13g2_decap_8 FILLER_2_630 ();
 sg13g2_decap_8 FILLER_2_637 ();
 sg13g2_decap_8 FILLER_2_644 ();
 sg13g2_decap_8 FILLER_2_651 ();
 sg13g2_decap_8 FILLER_2_658 ();
 sg13g2_decap_8 FILLER_2_665 ();
 sg13g2_decap_8 FILLER_2_672 ();
 sg13g2_decap_8 FILLER_2_679 ();
 sg13g2_decap_8 FILLER_2_686 ();
 sg13g2_decap_8 FILLER_2_693 ();
 sg13g2_decap_8 FILLER_2_700 ();
 sg13g2_decap_8 FILLER_2_707 ();
 sg13g2_decap_8 FILLER_2_714 ();
 sg13g2_decap_8 FILLER_2_721 ();
 sg13g2_decap_8 FILLER_2_728 ();
 sg13g2_decap_8 FILLER_2_735 ();
 sg13g2_decap_8 FILLER_2_742 ();
 sg13g2_decap_8 FILLER_2_749 ();
 sg13g2_decap_8 FILLER_2_756 ();
 sg13g2_decap_8 FILLER_2_763 ();
 sg13g2_decap_8 FILLER_2_770 ();
 sg13g2_decap_8 FILLER_2_777 ();
 sg13g2_decap_8 FILLER_2_784 ();
 sg13g2_decap_8 FILLER_2_791 ();
 sg13g2_decap_8 FILLER_2_798 ();
 sg13g2_decap_8 FILLER_2_805 ();
 sg13g2_decap_8 FILLER_2_812 ();
 sg13g2_decap_8 FILLER_2_819 ();
 sg13g2_decap_8 FILLER_2_826 ();
 sg13g2_decap_8 FILLER_2_833 ();
 sg13g2_decap_8 FILLER_2_840 ();
 sg13g2_decap_8 FILLER_2_847 ();
 sg13g2_decap_8 FILLER_2_854 ();
 sg13g2_fill_1 FILLER_2_861 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_fill_1 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_fill_1 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_decap_8 FILLER_5_427 ();
 sg13g2_decap_8 FILLER_5_434 ();
 sg13g2_decap_8 FILLER_5_441 ();
 sg13g2_decap_8 FILLER_5_448 ();
 sg13g2_decap_8 FILLER_5_455 ();
 sg13g2_decap_8 FILLER_5_462 ();
 sg13g2_decap_8 FILLER_5_469 ();
 sg13g2_decap_8 FILLER_5_476 ();
 sg13g2_decap_8 FILLER_5_483 ();
 sg13g2_decap_8 FILLER_5_490 ();
 sg13g2_decap_8 FILLER_5_497 ();
 sg13g2_decap_8 FILLER_5_504 ();
 sg13g2_decap_8 FILLER_5_511 ();
 sg13g2_decap_8 FILLER_5_518 ();
 sg13g2_decap_8 FILLER_5_525 ();
 sg13g2_decap_8 FILLER_5_532 ();
 sg13g2_decap_8 FILLER_5_539 ();
 sg13g2_decap_8 FILLER_5_546 ();
 sg13g2_decap_8 FILLER_5_553 ();
 sg13g2_decap_8 FILLER_5_560 ();
 sg13g2_decap_8 FILLER_5_567 ();
 sg13g2_decap_8 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_581 ();
 sg13g2_decap_8 FILLER_5_588 ();
 sg13g2_decap_8 FILLER_5_595 ();
 sg13g2_decap_8 FILLER_5_602 ();
 sg13g2_decap_8 FILLER_5_609 ();
 sg13g2_decap_8 FILLER_5_616 ();
 sg13g2_decap_8 FILLER_5_623 ();
 sg13g2_decap_8 FILLER_5_630 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_8 FILLER_5_672 ();
 sg13g2_decap_8 FILLER_5_679 ();
 sg13g2_decap_8 FILLER_5_686 ();
 sg13g2_decap_8 FILLER_5_693 ();
 sg13g2_decap_8 FILLER_5_700 ();
 sg13g2_decap_8 FILLER_5_707 ();
 sg13g2_decap_8 FILLER_5_714 ();
 sg13g2_decap_8 FILLER_5_721 ();
 sg13g2_decap_8 FILLER_5_728 ();
 sg13g2_decap_8 FILLER_5_735 ();
 sg13g2_decap_8 FILLER_5_742 ();
 sg13g2_decap_8 FILLER_5_749 ();
 sg13g2_decap_8 FILLER_5_756 ();
 sg13g2_decap_8 FILLER_5_763 ();
 sg13g2_decap_8 FILLER_5_770 ();
 sg13g2_decap_8 FILLER_5_777 ();
 sg13g2_decap_8 FILLER_5_784 ();
 sg13g2_decap_8 FILLER_5_791 ();
 sg13g2_decap_8 FILLER_5_798 ();
 sg13g2_decap_8 FILLER_5_805 ();
 sg13g2_decap_8 FILLER_5_812 ();
 sg13g2_decap_8 FILLER_5_819 ();
 sg13g2_decap_8 FILLER_5_826 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_decap_8 FILLER_5_847 ();
 sg13g2_decap_8 FILLER_5_854 ();
 sg13g2_fill_1 FILLER_5_861 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_fill_1 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_fill_1 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_fill_1 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_fill_1 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_decap_8 FILLER_10_406 ();
 sg13g2_decap_8 FILLER_10_413 ();
 sg13g2_decap_8 FILLER_10_420 ();
 sg13g2_decap_8 FILLER_10_427 ();
 sg13g2_decap_8 FILLER_10_434 ();
 sg13g2_decap_8 FILLER_10_441 ();
 sg13g2_decap_8 FILLER_10_448 ();
 sg13g2_decap_8 FILLER_10_455 ();
 sg13g2_decap_8 FILLER_10_462 ();
 sg13g2_decap_8 FILLER_10_469 ();
 sg13g2_decap_8 FILLER_10_476 ();
 sg13g2_decap_8 FILLER_10_483 ();
 sg13g2_decap_8 FILLER_10_490 ();
 sg13g2_decap_8 FILLER_10_497 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_8 FILLER_10_511 ();
 sg13g2_decap_8 FILLER_10_518 ();
 sg13g2_decap_8 FILLER_10_525 ();
 sg13g2_decap_8 FILLER_10_532 ();
 sg13g2_decap_8 FILLER_10_539 ();
 sg13g2_decap_8 FILLER_10_546 ();
 sg13g2_decap_8 FILLER_10_553 ();
 sg13g2_decap_8 FILLER_10_560 ();
 sg13g2_decap_8 FILLER_10_567 ();
 sg13g2_decap_8 FILLER_10_574 ();
 sg13g2_decap_8 FILLER_10_581 ();
 sg13g2_decap_8 FILLER_10_588 ();
 sg13g2_decap_8 FILLER_10_595 ();
 sg13g2_decap_8 FILLER_10_602 ();
 sg13g2_decap_8 FILLER_10_609 ();
 sg13g2_decap_8 FILLER_10_616 ();
 sg13g2_decap_8 FILLER_10_623 ();
 sg13g2_decap_8 FILLER_10_630 ();
 sg13g2_decap_8 FILLER_10_637 ();
 sg13g2_decap_8 FILLER_10_644 ();
 sg13g2_decap_8 FILLER_10_651 ();
 sg13g2_decap_8 FILLER_10_658 ();
 sg13g2_decap_8 FILLER_10_665 ();
 sg13g2_decap_8 FILLER_10_672 ();
 sg13g2_decap_8 FILLER_10_679 ();
 sg13g2_decap_8 FILLER_10_686 ();
 sg13g2_decap_8 FILLER_10_693 ();
 sg13g2_decap_8 FILLER_10_700 ();
 sg13g2_decap_8 FILLER_10_707 ();
 sg13g2_decap_8 FILLER_10_714 ();
 sg13g2_decap_8 FILLER_10_721 ();
 sg13g2_decap_8 FILLER_10_728 ();
 sg13g2_decap_8 FILLER_10_735 ();
 sg13g2_decap_8 FILLER_10_742 ();
 sg13g2_decap_8 FILLER_10_749 ();
 sg13g2_decap_8 FILLER_10_756 ();
 sg13g2_decap_8 FILLER_10_763 ();
 sg13g2_decap_8 FILLER_10_770 ();
 sg13g2_decap_8 FILLER_10_777 ();
 sg13g2_decap_8 FILLER_10_784 ();
 sg13g2_decap_8 FILLER_10_791 ();
 sg13g2_decap_8 FILLER_10_798 ();
 sg13g2_decap_8 FILLER_10_805 ();
 sg13g2_decap_8 FILLER_10_812 ();
 sg13g2_decap_8 FILLER_10_819 ();
 sg13g2_decap_8 FILLER_10_826 ();
 sg13g2_decap_8 FILLER_10_833 ();
 sg13g2_decap_8 FILLER_10_840 ();
 sg13g2_decap_8 FILLER_10_847 ();
 sg13g2_decap_8 FILLER_10_854 ();
 sg13g2_fill_1 FILLER_10_861 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_fill_1 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_decap_8 FILLER_12_427 ();
 sg13g2_decap_8 FILLER_12_434 ();
 sg13g2_decap_8 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_448 ();
 sg13g2_decap_8 FILLER_12_455 ();
 sg13g2_decap_8 FILLER_12_462 ();
 sg13g2_decap_8 FILLER_12_469 ();
 sg13g2_decap_8 FILLER_12_476 ();
 sg13g2_decap_8 FILLER_12_483 ();
 sg13g2_decap_8 FILLER_12_490 ();
 sg13g2_decap_8 FILLER_12_497 ();
 sg13g2_decap_8 FILLER_12_504 ();
 sg13g2_decap_8 FILLER_12_511 ();
 sg13g2_decap_8 FILLER_12_518 ();
 sg13g2_decap_8 FILLER_12_525 ();
 sg13g2_decap_8 FILLER_12_532 ();
 sg13g2_decap_8 FILLER_12_539 ();
 sg13g2_decap_8 FILLER_12_546 ();
 sg13g2_decap_8 FILLER_12_553 ();
 sg13g2_decap_8 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_decap_8 FILLER_12_574 ();
 sg13g2_decap_8 FILLER_12_581 ();
 sg13g2_decap_8 FILLER_12_588 ();
 sg13g2_decap_8 FILLER_12_595 ();
 sg13g2_decap_8 FILLER_12_602 ();
 sg13g2_decap_8 FILLER_12_609 ();
 sg13g2_decap_8 FILLER_12_616 ();
 sg13g2_decap_8 FILLER_12_623 ();
 sg13g2_decap_8 FILLER_12_630 ();
 sg13g2_decap_8 FILLER_12_637 ();
 sg13g2_decap_8 FILLER_12_644 ();
 sg13g2_decap_8 FILLER_12_651 ();
 sg13g2_decap_8 FILLER_12_658 ();
 sg13g2_decap_8 FILLER_12_665 ();
 sg13g2_decap_8 FILLER_12_672 ();
 sg13g2_decap_8 FILLER_12_679 ();
 sg13g2_decap_8 FILLER_12_686 ();
 sg13g2_decap_8 FILLER_12_693 ();
 sg13g2_decap_8 FILLER_12_700 ();
 sg13g2_decap_8 FILLER_12_707 ();
 sg13g2_decap_8 FILLER_12_714 ();
 sg13g2_decap_8 FILLER_12_721 ();
 sg13g2_decap_8 FILLER_12_728 ();
 sg13g2_decap_8 FILLER_12_735 ();
 sg13g2_decap_8 FILLER_12_742 ();
 sg13g2_decap_8 FILLER_12_749 ();
 sg13g2_decap_8 FILLER_12_756 ();
 sg13g2_decap_8 FILLER_12_763 ();
 sg13g2_decap_8 FILLER_12_770 ();
 sg13g2_decap_8 FILLER_12_777 ();
 sg13g2_decap_8 FILLER_12_784 ();
 sg13g2_decap_8 FILLER_12_791 ();
 sg13g2_decap_8 FILLER_12_798 ();
 sg13g2_decap_8 FILLER_12_805 ();
 sg13g2_decap_8 FILLER_12_812 ();
 sg13g2_decap_8 FILLER_12_819 ();
 sg13g2_decap_8 FILLER_12_826 ();
 sg13g2_decap_8 FILLER_12_833 ();
 sg13g2_decap_8 FILLER_12_840 ();
 sg13g2_decap_8 FILLER_12_847 ();
 sg13g2_decap_8 FILLER_12_854 ();
 sg13g2_fill_1 FILLER_12_861 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_fill_1 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_fill_1 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_decap_8 FILLER_15_406 ();
 sg13g2_decap_8 FILLER_15_413 ();
 sg13g2_decap_8 FILLER_15_420 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_8 FILLER_15_434 ();
 sg13g2_decap_8 FILLER_15_441 ();
 sg13g2_decap_8 FILLER_15_448 ();
 sg13g2_decap_8 FILLER_15_455 ();
 sg13g2_decap_8 FILLER_15_462 ();
 sg13g2_decap_8 FILLER_15_469 ();
 sg13g2_decap_8 FILLER_15_476 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_8 FILLER_15_497 ();
 sg13g2_decap_8 FILLER_15_504 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_decap_8 FILLER_15_518 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_8 FILLER_15_532 ();
 sg13g2_decap_8 FILLER_15_539 ();
 sg13g2_decap_8 FILLER_15_546 ();
 sg13g2_decap_8 FILLER_15_553 ();
 sg13g2_decap_8 FILLER_15_560 ();
 sg13g2_decap_8 FILLER_15_567 ();
 sg13g2_decap_8 FILLER_15_574 ();
 sg13g2_decap_8 FILLER_15_581 ();
 sg13g2_decap_8 FILLER_15_588 ();
 sg13g2_decap_8 FILLER_15_595 ();
 sg13g2_decap_8 FILLER_15_602 ();
 sg13g2_decap_8 FILLER_15_609 ();
 sg13g2_decap_8 FILLER_15_616 ();
 sg13g2_decap_8 FILLER_15_623 ();
 sg13g2_decap_8 FILLER_15_630 ();
 sg13g2_decap_8 FILLER_15_637 ();
 sg13g2_decap_8 FILLER_15_644 ();
 sg13g2_decap_8 FILLER_15_651 ();
 sg13g2_decap_8 FILLER_15_658 ();
 sg13g2_decap_8 FILLER_15_665 ();
 sg13g2_decap_8 FILLER_15_672 ();
 sg13g2_decap_8 FILLER_15_679 ();
 sg13g2_decap_8 FILLER_15_686 ();
 sg13g2_decap_8 FILLER_15_693 ();
 sg13g2_decap_8 FILLER_15_700 ();
 sg13g2_decap_8 FILLER_15_707 ();
 sg13g2_decap_8 FILLER_15_714 ();
 sg13g2_decap_8 FILLER_15_721 ();
 sg13g2_decap_8 FILLER_15_728 ();
 sg13g2_decap_8 FILLER_15_735 ();
 sg13g2_decap_8 FILLER_15_742 ();
 sg13g2_decap_8 FILLER_15_749 ();
 sg13g2_decap_8 FILLER_15_756 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_8 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_777 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_decap_8 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_798 ();
 sg13g2_decap_8 FILLER_15_805 ();
 sg13g2_decap_8 FILLER_15_812 ();
 sg13g2_decap_8 FILLER_15_819 ();
 sg13g2_decap_8 FILLER_15_826 ();
 sg13g2_decap_8 FILLER_15_833 ();
 sg13g2_decap_8 FILLER_15_840 ();
 sg13g2_decap_8 FILLER_15_847 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_fill_1 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_fill_1 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_fill_1 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_fill_1 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_fill_1 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_decap_8 FILLER_20_266 ();
 sg13g2_decap_8 FILLER_20_273 ();
 sg13g2_decap_8 FILLER_20_280 ();
 sg13g2_decap_8 FILLER_20_287 ();
 sg13g2_decap_8 FILLER_20_294 ();
 sg13g2_decap_8 FILLER_20_301 ();
 sg13g2_decap_8 FILLER_20_308 ();
 sg13g2_decap_8 FILLER_20_315 ();
 sg13g2_decap_8 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_decap_8 FILLER_20_406 ();
 sg13g2_decap_8 FILLER_20_413 ();
 sg13g2_decap_8 FILLER_20_420 ();
 sg13g2_decap_8 FILLER_20_427 ();
 sg13g2_decap_8 FILLER_20_434 ();
 sg13g2_decap_8 FILLER_20_441 ();
 sg13g2_decap_8 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_455 ();
 sg13g2_decap_8 FILLER_20_462 ();
 sg13g2_decap_8 FILLER_20_469 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_decap_8 FILLER_20_483 ();
 sg13g2_decap_8 FILLER_20_490 ();
 sg13g2_decap_8 FILLER_20_497 ();
 sg13g2_decap_8 FILLER_20_504 ();
 sg13g2_decap_8 FILLER_20_511 ();
 sg13g2_decap_8 FILLER_20_518 ();
 sg13g2_decap_8 FILLER_20_525 ();
 sg13g2_decap_8 FILLER_20_532 ();
 sg13g2_decap_8 FILLER_20_539 ();
 sg13g2_decap_8 FILLER_20_546 ();
 sg13g2_decap_8 FILLER_20_553 ();
 sg13g2_decap_8 FILLER_20_560 ();
 sg13g2_decap_8 FILLER_20_567 ();
 sg13g2_decap_8 FILLER_20_574 ();
 sg13g2_decap_8 FILLER_20_581 ();
 sg13g2_decap_8 FILLER_20_588 ();
 sg13g2_decap_8 FILLER_20_595 ();
 sg13g2_decap_8 FILLER_20_602 ();
 sg13g2_decap_8 FILLER_20_609 ();
 sg13g2_decap_8 FILLER_20_616 ();
 sg13g2_decap_8 FILLER_20_623 ();
 sg13g2_decap_8 FILLER_20_630 ();
 sg13g2_decap_8 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_644 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_decap_8 FILLER_20_672 ();
 sg13g2_decap_8 FILLER_20_679 ();
 sg13g2_decap_8 FILLER_20_686 ();
 sg13g2_decap_8 FILLER_20_693 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_8 FILLER_20_714 ();
 sg13g2_decap_8 FILLER_20_721 ();
 sg13g2_decap_8 FILLER_20_728 ();
 sg13g2_decap_8 FILLER_20_735 ();
 sg13g2_decap_8 FILLER_20_742 ();
 sg13g2_decap_8 FILLER_20_749 ();
 sg13g2_decap_8 FILLER_20_756 ();
 sg13g2_decap_8 FILLER_20_763 ();
 sg13g2_decap_8 FILLER_20_770 ();
 sg13g2_decap_8 FILLER_20_777 ();
 sg13g2_decap_8 FILLER_20_784 ();
 sg13g2_decap_8 FILLER_20_791 ();
 sg13g2_decap_8 FILLER_20_798 ();
 sg13g2_decap_8 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_812 ();
 sg13g2_decap_8 FILLER_20_819 ();
 sg13g2_decap_8 FILLER_20_826 ();
 sg13g2_decap_8 FILLER_20_833 ();
 sg13g2_decap_8 FILLER_20_840 ();
 sg13g2_decap_8 FILLER_20_847 ();
 sg13g2_decap_8 FILLER_20_854 ();
 sg13g2_fill_1 FILLER_20_861 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_fill_1 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_4 FILLER_22_245 ();
 sg13g2_fill_1 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_286 ();
 sg13g2_decap_8 FILLER_22_293 ();
 sg13g2_decap_8 FILLER_22_300 ();
 sg13g2_decap_8 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_314 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_fill_1 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_416 ();
 sg13g2_decap_8 FILLER_22_423 ();
 sg13g2_decap_8 FILLER_22_430 ();
 sg13g2_decap_8 FILLER_22_437 ();
 sg13g2_decap_8 FILLER_22_444 ();
 sg13g2_decap_8 FILLER_22_451 ();
 sg13g2_decap_8 FILLER_22_458 ();
 sg13g2_decap_8 FILLER_22_465 ();
 sg13g2_decap_8 FILLER_22_472 ();
 sg13g2_decap_8 FILLER_22_479 ();
 sg13g2_decap_8 FILLER_22_486 ();
 sg13g2_decap_8 FILLER_22_493 ();
 sg13g2_decap_8 FILLER_22_500 ();
 sg13g2_decap_8 FILLER_22_507 ();
 sg13g2_decap_8 FILLER_22_514 ();
 sg13g2_decap_8 FILLER_22_521 ();
 sg13g2_decap_8 FILLER_22_528 ();
 sg13g2_decap_8 FILLER_22_535 ();
 sg13g2_decap_8 FILLER_22_542 ();
 sg13g2_decap_8 FILLER_22_549 ();
 sg13g2_decap_8 FILLER_22_556 ();
 sg13g2_decap_8 FILLER_22_563 ();
 sg13g2_decap_8 FILLER_22_570 ();
 sg13g2_decap_8 FILLER_22_577 ();
 sg13g2_decap_8 FILLER_22_584 ();
 sg13g2_decap_8 FILLER_22_591 ();
 sg13g2_decap_8 FILLER_22_598 ();
 sg13g2_decap_8 FILLER_22_605 ();
 sg13g2_decap_8 FILLER_22_612 ();
 sg13g2_decap_8 FILLER_22_619 ();
 sg13g2_decap_8 FILLER_22_626 ();
 sg13g2_decap_8 FILLER_22_633 ();
 sg13g2_decap_8 FILLER_22_640 ();
 sg13g2_decap_8 FILLER_22_647 ();
 sg13g2_decap_8 FILLER_22_654 ();
 sg13g2_decap_8 FILLER_22_661 ();
 sg13g2_decap_8 FILLER_22_668 ();
 sg13g2_decap_8 FILLER_22_675 ();
 sg13g2_decap_8 FILLER_22_682 ();
 sg13g2_decap_8 FILLER_22_689 ();
 sg13g2_decap_8 FILLER_22_696 ();
 sg13g2_decap_8 FILLER_22_703 ();
 sg13g2_decap_8 FILLER_22_710 ();
 sg13g2_decap_8 FILLER_22_717 ();
 sg13g2_decap_8 FILLER_22_724 ();
 sg13g2_decap_8 FILLER_22_731 ();
 sg13g2_decap_8 FILLER_22_738 ();
 sg13g2_decap_8 FILLER_22_745 ();
 sg13g2_decap_8 FILLER_22_752 ();
 sg13g2_decap_8 FILLER_22_759 ();
 sg13g2_decap_8 FILLER_22_766 ();
 sg13g2_decap_8 FILLER_22_773 ();
 sg13g2_decap_8 FILLER_22_780 ();
 sg13g2_decap_8 FILLER_22_787 ();
 sg13g2_decap_8 FILLER_22_794 ();
 sg13g2_decap_8 FILLER_22_801 ();
 sg13g2_decap_8 FILLER_22_808 ();
 sg13g2_decap_8 FILLER_22_815 ();
 sg13g2_decap_8 FILLER_22_822 ();
 sg13g2_decap_8 FILLER_22_829 ();
 sg13g2_decap_8 FILLER_22_836 ();
 sg13g2_decap_8 FILLER_22_843 ();
 sg13g2_decap_8 FILLER_22_850 ();
 sg13g2_decap_4 FILLER_22_857 ();
 sg13g2_fill_1 FILLER_22_861 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_4 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_4 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_193 ();
 sg13g2_decap_4 FILLER_23_210 ();
 sg13g2_fill_1 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_4 FILLER_23_231 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_267 ();
 sg13g2_decap_8 FILLER_23_274 ();
 sg13g2_fill_2 FILLER_23_281 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_2 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_fill_2 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_369 ();
 sg13g2_fill_2 FILLER_23_376 ();
 sg13g2_fill_1 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_382 ();
 sg13g2_fill_1 FILLER_23_386 ();
 sg13g2_fill_2 FILLER_23_402 ();
 sg13g2_fill_2 FILLER_23_428 ();
 sg13g2_decap_8 FILLER_23_436 ();
 sg13g2_decap_4 FILLER_23_452 ();
 sg13g2_fill_1 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_decap_4 FILLER_23_508 ();
 sg13g2_fill_1 FILLER_23_512 ();
 sg13g2_decap_8 FILLER_23_523 ();
 sg13g2_decap_8 FILLER_23_530 ();
 sg13g2_decap_8 FILLER_23_537 ();
 sg13g2_fill_1 FILLER_23_544 ();
 sg13g2_decap_8 FILLER_23_554 ();
 sg13g2_decap_4 FILLER_23_561 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_fill_1 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_fill_1 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_93 ();
 sg13g2_decap_4 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_104 ();
 sg13g2_decap_4 FILLER_24_115 ();
 sg13g2_fill_2 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_fill_2 FILLER_24_228 ();
 sg13g2_fill_1 FILLER_24_230 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_fill_1 FILLER_24_282 ();
 sg13g2_decap_4 FILLER_24_365 ();
 sg13g2_fill_2 FILLER_24_369 ();
 sg13g2_fill_1 FILLER_24_399 ();
 sg13g2_fill_1 FILLER_24_456 ();
 sg13g2_fill_2 FILLER_24_489 ();
 sg13g2_fill_2 FILLER_24_582 ();
 sg13g2_decap_8 FILLER_24_597 ();
 sg13g2_decap_8 FILLER_24_604 ();
 sg13g2_decap_8 FILLER_24_611 ();
 sg13g2_decap_8 FILLER_24_618 ();
 sg13g2_decap_8 FILLER_24_625 ();
 sg13g2_decap_8 FILLER_24_632 ();
 sg13g2_decap_8 FILLER_24_639 ();
 sg13g2_decap_8 FILLER_24_646 ();
 sg13g2_decap_8 FILLER_24_653 ();
 sg13g2_decap_8 FILLER_24_660 ();
 sg13g2_decap_8 FILLER_24_667 ();
 sg13g2_decap_8 FILLER_24_674 ();
 sg13g2_decap_8 FILLER_24_681 ();
 sg13g2_decap_8 FILLER_24_688 ();
 sg13g2_decap_8 FILLER_24_695 ();
 sg13g2_decap_8 FILLER_24_702 ();
 sg13g2_decap_8 FILLER_24_709 ();
 sg13g2_decap_8 FILLER_24_716 ();
 sg13g2_decap_8 FILLER_24_723 ();
 sg13g2_decap_8 FILLER_24_730 ();
 sg13g2_decap_8 FILLER_24_737 ();
 sg13g2_decap_8 FILLER_24_744 ();
 sg13g2_decap_8 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_758 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_8 FILLER_24_772 ();
 sg13g2_decap_8 FILLER_24_779 ();
 sg13g2_decap_8 FILLER_24_786 ();
 sg13g2_decap_8 FILLER_24_793 ();
 sg13g2_decap_8 FILLER_24_800 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_8 FILLER_24_814 ();
 sg13g2_decap_8 FILLER_24_821 ();
 sg13g2_decap_8 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_24_835 ();
 sg13g2_decap_8 FILLER_24_842 ();
 sg13g2_decap_8 FILLER_24_849 ();
 sg13g2_decap_4 FILLER_24_856 ();
 sg13g2_fill_2 FILLER_24_860 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_decap_4 FILLER_25_38 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_84 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_fill_2 FILLER_25_170 ();
 sg13g2_fill_1 FILLER_25_172 ();
 sg13g2_fill_2 FILLER_25_179 ();
 sg13g2_fill_1 FILLER_25_181 ();
 sg13g2_fill_2 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_317 ();
 sg13g2_fill_2 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_360 ();
 sg13g2_fill_2 FILLER_25_382 ();
 sg13g2_fill_2 FILLER_25_399 ();
 sg13g2_fill_1 FILLER_25_428 ();
 sg13g2_fill_1 FILLER_25_476 ();
 sg13g2_fill_2 FILLER_25_486 ();
 sg13g2_fill_2 FILLER_25_516 ();
 sg13g2_decap_8 FILLER_25_527 ();
 sg13g2_fill_1 FILLER_25_534 ();
 sg13g2_decap_4 FILLER_25_569 ();
 sg13g2_fill_1 FILLER_25_573 ();
 sg13g2_decap_8 FILLER_25_618 ();
 sg13g2_decap_8 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_632 ();
 sg13g2_decap_8 FILLER_25_639 ();
 sg13g2_decap_8 FILLER_25_646 ();
 sg13g2_decap_8 FILLER_25_653 ();
 sg13g2_decap_8 FILLER_25_660 ();
 sg13g2_decap_8 FILLER_25_667 ();
 sg13g2_decap_8 FILLER_25_674 ();
 sg13g2_decap_8 FILLER_25_681 ();
 sg13g2_decap_8 FILLER_25_688 ();
 sg13g2_decap_8 FILLER_25_695 ();
 sg13g2_decap_8 FILLER_25_702 ();
 sg13g2_decap_8 FILLER_25_709 ();
 sg13g2_decap_8 FILLER_25_716 ();
 sg13g2_decap_8 FILLER_25_723 ();
 sg13g2_decap_8 FILLER_25_730 ();
 sg13g2_decap_8 FILLER_25_737 ();
 sg13g2_decap_8 FILLER_25_744 ();
 sg13g2_decap_8 FILLER_25_751 ();
 sg13g2_decap_8 FILLER_25_758 ();
 sg13g2_decap_8 FILLER_25_765 ();
 sg13g2_decap_8 FILLER_25_772 ();
 sg13g2_decap_8 FILLER_25_779 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_decap_8 FILLER_25_814 ();
 sg13g2_decap_8 FILLER_25_821 ();
 sg13g2_decap_8 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_835 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_4 FILLER_25_856 ();
 sg13g2_fill_2 FILLER_25_860 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_63 ();
 sg13g2_decap_4 FILLER_26_106 ();
 sg13g2_fill_2 FILLER_26_110 ();
 sg13g2_fill_2 FILLER_26_201 ();
 sg13g2_fill_1 FILLER_26_257 ();
 sg13g2_fill_1 FILLER_26_275 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_decap_4 FILLER_26_312 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_414 ();
 sg13g2_fill_2 FILLER_26_501 ();
 sg13g2_fill_2 FILLER_26_528 ();
 sg13g2_fill_1 FILLER_26_530 ();
 sg13g2_fill_1 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_621 ();
 sg13g2_decap_8 FILLER_26_628 ();
 sg13g2_decap_8 FILLER_26_635 ();
 sg13g2_decap_8 FILLER_26_642 ();
 sg13g2_decap_8 FILLER_26_649 ();
 sg13g2_decap_8 FILLER_26_656 ();
 sg13g2_decap_8 FILLER_26_663 ();
 sg13g2_decap_8 FILLER_26_670 ();
 sg13g2_decap_8 FILLER_26_677 ();
 sg13g2_decap_8 FILLER_26_684 ();
 sg13g2_decap_8 FILLER_26_691 ();
 sg13g2_decap_8 FILLER_26_698 ();
 sg13g2_decap_8 FILLER_26_705 ();
 sg13g2_decap_8 FILLER_26_712 ();
 sg13g2_decap_8 FILLER_26_719 ();
 sg13g2_decap_8 FILLER_26_726 ();
 sg13g2_decap_8 FILLER_26_733 ();
 sg13g2_decap_8 FILLER_26_740 ();
 sg13g2_decap_8 FILLER_26_747 ();
 sg13g2_decap_8 FILLER_26_754 ();
 sg13g2_decap_8 FILLER_26_761 ();
 sg13g2_decap_8 FILLER_26_768 ();
 sg13g2_decap_8 FILLER_26_775 ();
 sg13g2_decap_8 FILLER_26_782 ();
 sg13g2_decap_8 FILLER_26_789 ();
 sg13g2_decap_8 FILLER_26_796 ();
 sg13g2_decap_8 FILLER_26_803 ();
 sg13g2_decap_8 FILLER_26_810 ();
 sg13g2_decap_8 FILLER_26_817 ();
 sg13g2_decap_8 FILLER_26_824 ();
 sg13g2_decap_8 FILLER_26_831 ();
 sg13g2_decap_8 FILLER_26_838 ();
 sg13g2_decap_8 FILLER_26_845 ();
 sg13g2_decap_8 FILLER_26_852 ();
 sg13g2_fill_2 FILLER_26_859 ();
 sg13g2_fill_1 FILLER_26_861 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_fill_1 FILLER_27_88 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_134 ();
 sg13g2_fill_1 FILLER_27_136 ();
 sg13g2_fill_1 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_fill_1 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_decap_4 FILLER_27_332 ();
 sg13g2_fill_2 FILLER_27_336 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_decap_8 FILLER_27_358 ();
 sg13g2_fill_2 FILLER_27_377 ();
 sg13g2_fill_2 FILLER_27_392 ();
 sg13g2_fill_1 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_404 ();
 sg13g2_fill_1 FILLER_27_411 ();
 sg13g2_fill_2 FILLER_27_432 ();
 sg13g2_fill_1 FILLER_27_434 ();
 sg13g2_fill_2 FILLER_27_440 ();
 sg13g2_fill_1 FILLER_27_554 ();
 sg13g2_fill_1 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_617 ();
 sg13g2_decap_8 FILLER_27_624 ();
 sg13g2_decap_8 FILLER_27_631 ();
 sg13g2_fill_2 FILLER_27_638 ();
 sg13g2_decap_8 FILLER_27_643 ();
 sg13g2_decap_8 FILLER_27_650 ();
 sg13g2_fill_2 FILLER_27_657 ();
 sg13g2_decap_8 FILLER_27_668 ();
 sg13g2_decap_8 FILLER_27_684 ();
 sg13g2_decap_8 FILLER_27_691 ();
 sg13g2_decap_8 FILLER_27_698 ();
 sg13g2_decap_8 FILLER_27_705 ();
 sg13g2_decap_8 FILLER_27_712 ();
 sg13g2_decap_8 FILLER_27_719 ();
 sg13g2_decap_8 FILLER_27_726 ();
 sg13g2_decap_8 FILLER_27_733 ();
 sg13g2_decap_8 FILLER_27_740 ();
 sg13g2_decap_8 FILLER_27_747 ();
 sg13g2_decap_8 FILLER_27_754 ();
 sg13g2_decap_8 FILLER_27_761 ();
 sg13g2_decap_8 FILLER_27_768 ();
 sg13g2_decap_8 FILLER_27_775 ();
 sg13g2_decap_8 FILLER_27_782 ();
 sg13g2_decap_8 FILLER_27_789 ();
 sg13g2_decap_8 FILLER_27_796 ();
 sg13g2_decap_8 FILLER_27_803 ();
 sg13g2_decap_8 FILLER_27_810 ();
 sg13g2_decap_8 FILLER_27_817 ();
 sg13g2_decap_8 FILLER_27_824 ();
 sg13g2_decap_8 FILLER_27_831 ();
 sg13g2_decap_8 FILLER_27_838 ();
 sg13g2_decap_8 FILLER_27_845 ();
 sg13g2_decap_8 FILLER_27_852 ();
 sg13g2_fill_2 FILLER_27_859 ();
 sg13g2_fill_1 FILLER_27_861 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_2 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_92 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_fill_2 FILLER_28_125 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_fill_1 FILLER_28_230 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_290 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_decap_8 FILLER_28_327 ();
 sg13g2_decap_4 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_decap_4 FILLER_28_397 ();
 sg13g2_fill_1 FILLER_28_401 ();
 sg13g2_decap_4 FILLER_28_411 ();
 sg13g2_fill_1 FILLER_28_456 ();
 sg13g2_fill_2 FILLER_28_493 ();
 sg13g2_fill_1 FILLER_28_495 ();
 sg13g2_fill_2 FILLER_28_506 ();
 sg13g2_fill_1 FILLER_28_508 ();
 sg13g2_decap_8 FILLER_28_527 ();
 sg13g2_fill_2 FILLER_28_534 ();
 sg13g2_decap_4 FILLER_28_539 ();
 sg13g2_decap_4 FILLER_28_555 ();
 sg13g2_fill_1 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_563 ();
 sg13g2_decap_8 FILLER_28_576 ();
 sg13g2_fill_1 FILLER_28_583 ();
 sg13g2_fill_1 FILLER_28_624 ();
 sg13g2_decap_4 FILLER_28_630 ();
 sg13g2_decap_4 FILLER_28_695 ();
 sg13g2_decap_8 FILLER_28_712 ();
 sg13g2_decap_8 FILLER_28_719 ();
 sg13g2_decap_8 FILLER_28_726 ();
 sg13g2_decap_8 FILLER_28_733 ();
 sg13g2_decap_8 FILLER_28_740 ();
 sg13g2_decap_8 FILLER_28_747 ();
 sg13g2_decap_8 FILLER_28_754 ();
 sg13g2_decap_8 FILLER_28_761 ();
 sg13g2_decap_8 FILLER_28_768 ();
 sg13g2_decap_8 FILLER_28_775 ();
 sg13g2_decap_8 FILLER_28_782 ();
 sg13g2_decap_8 FILLER_28_789 ();
 sg13g2_decap_8 FILLER_28_796 ();
 sg13g2_decap_8 FILLER_28_803 ();
 sg13g2_decap_8 FILLER_28_810 ();
 sg13g2_decap_8 FILLER_28_817 ();
 sg13g2_decap_8 FILLER_28_824 ();
 sg13g2_decap_8 FILLER_28_831 ();
 sg13g2_decap_8 FILLER_28_838 ();
 sg13g2_decap_8 FILLER_28_845 ();
 sg13g2_decap_8 FILLER_28_852 ();
 sg13g2_fill_2 FILLER_28_859 ();
 sg13g2_fill_1 FILLER_28_861 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_82 ();
 sg13g2_fill_1 FILLER_29_86 ();
 sg13g2_fill_2 FILLER_29_124 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_fill_2 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_206 ();
 sg13g2_decap_8 FILLER_29_234 ();
 sg13g2_decap_4 FILLER_29_241 ();
 sg13g2_decap_4 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_307 ();
 sg13g2_fill_1 FILLER_29_358 ();
 sg13g2_decap_4 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_1 FILLER_29_438 ();
 sg13g2_fill_2 FILLER_29_479 ();
 sg13g2_fill_2 FILLER_29_526 ();
 sg13g2_fill_1 FILLER_29_528 ();
 sg13g2_fill_2 FILLER_29_578 ();
 sg13g2_fill_1 FILLER_29_611 ();
 sg13g2_fill_2 FILLER_29_639 ();
 sg13g2_fill_2 FILLER_29_653 ();
 sg13g2_fill_1 FILLER_29_664 ();
 sg13g2_decap_8 FILLER_29_727 ();
 sg13g2_decap_8 FILLER_29_734 ();
 sg13g2_decap_8 FILLER_29_741 ();
 sg13g2_decap_8 FILLER_29_748 ();
 sg13g2_decap_8 FILLER_29_755 ();
 sg13g2_decap_8 FILLER_29_762 ();
 sg13g2_decap_8 FILLER_29_769 ();
 sg13g2_decap_8 FILLER_29_776 ();
 sg13g2_decap_8 FILLER_29_783 ();
 sg13g2_decap_8 FILLER_29_790 ();
 sg13g2_decap_8 FILLER_29_797 ();
 sg13g2_decap_8 FILLER_29_804 ();
 sg13g2_decap_8 FILLER_29_811 ();
 sg13g2_decap_8 FILLER_29_818 ();
 sg13g2_decap_8 FILLER_29_825 ();
 sg13g2_decap_8 FILLER_29_832 ();
 sg13g2_decap_8 FILLER_29_839 ();
 sg13g2_decap_8 FILLER_29_846 ();
 sg13g2_decap_8 FILLER_29_853 ();
 sg13g2_fill_2 FILLER_29_860 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_40 ();
 sg13g2_fill_2 FILLER_30_113 ();
 sg13g2_fill_1 FILLER_30_115 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_1 FILLER_30_225 ();
 sg13g2_fill_2 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_330 ();
 sg13g2_fill_2 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_396 ();
 sg13g2_fill_2 FILLER_30_410 ();
 sg13g2_fill_1 FILLER_30_421 ();
 sg13g2_fill_2 FILLER_30_440 ();
 sg13g2_fill_1 FILLER_30_442 ();
 sg13g2_decap_4 FILLER_30_448 ();
 sg13g2_fill_2 FILLER_30_452 ();
 sg13g2_fill_1 FILLER_30_517 ();
 sg13g2_fill_1 FILLER_30_549 ();
 sg13g2_fill_2 FILLER_30_600 ();
 sg13g2_fill_1 FILLER_30_602 ();
 sg13g2_fill_1 FILLER_30_661 ();
 sg13g2_fill_1 FILLER_30_683 ();
 sg13g2_fill_2 FILLER_30_699 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_fill_1 FILLER_30_861 ();
 sg13g2_fill_2 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_2 ();
 sg13g2_decap_4 FILLER_31_62 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_decap_4 FILLER_31_114 ();
 sg13g2_fill_2 FILLER_31_132 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_fill_2 FILLER_31_168 ();
 sg13g2_fill_1 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_decap_4 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_244 ();
 sg13g2_decap_4 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_fill_2 FILLER_31_393 ();
 sg13g2_fill_2 FILLER_31_417 ();
 sg13g2_fill_1 FILLER_31_462 ();
 sg13g2_decap_4 FILLER_31_489 ();
 sg13g2_fill_2 FILLER_31_537 ();
 sg13g2_fill_2 FILLER_31_567 ();
 sg13g2_fill_1 FILLER_31_590 ();
 sg13g2_fill_2 FILLER_31_623 ();
 sg13g2_fill_2 FILLER_31_670 ();
 sg13g2_fill_2 FILLER_31_690 ();
 sg13g2_fill_1 FILLER_31_692 ();
 sg13g2_decap_8 FILLER_31_729 ();
 sg13g2_decap_8 FILLER_31_736 ();
 sg13g2_decap_8 FILLER_31_743 ();
 sg13g2_decap_8 FILLER_31_750 ();
 sg13g2_decap_8 FILLER_31_757 ();
 sg13g2_decap_8 FILLER_31_764 ();
 sg13g2_decap_8 FILLER_31_771 ();
 sg13g2_decap_8 FILLER_31_778 ();
 sg13g2_decap_8 FILLER_31_785 ();
 sg13g2_decap_8 FILLER_31_792 ();
 sg13g2_decap_8 FILLER_31_799 ();
 sg13g2_decap_8 FILLER_31_806 ();
 sg13g2_decap_8 FILLER_31_813 ();
 sg13g2_decap_8 FILLER_31_820 ();
 sg13g2_decap_8 FILLER_31_827 ();
 sg13g2_decap_8 FILLER_31_834 ();
 sg13g2_decap_8 FILLER_31_841 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_8 FILLER_31_855 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_2 ();
 sg13g2_fill_2 FILLER_32_30 ();
 sg13g2_fill_1 FILLER_32_54 ();
 sg13g2_fill_1 FILLER_32_67 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_fill_1 FILLER_32_147 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_fill_2 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_302 ();
 sg13g2_decap_4 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_409 ();
 sg13g2_decap_4 FILLER_32_434 ();
 sg13g2_fill_2 FILLER_32_438 ();
 sg13g2_fill_2 FILLER_32_445 ();
 sg13g2_fill_1 FILLER_32_447 ();
 sg13g2_decap_8 FILLER_32_468 ();
 sg13g2_decap_4 FILLER_32_484 ();
 sg13g2_fill_2 FILLER_32_518 ();
 sg13g2_fill_2 FILLER_32_533 ();
 sg13g2_fill_2 FILLER_32_562 ();
 sg13g2_decap_8 FILLER_32_605 ();
 sg13g2_decap_4 FILLER_32_612 ();
 sg13g2_fill_2 FILLER_32_616 ();
 sg13g2_decap_4 FILLER_32_631 ();
 sg13g2_fill_2 FILLER_32_688 ();
 sg13g2_decap_8 FILLER_32_739 ();
 sg13g2_decap_8 FILLER_32_746 ();
 sg13g2_decap_8 FILLER_32_753 ();
 sg13g2_decap_8 FILLER_32_760 ();
 sg13g2_decap_8 FILLER_32_767 ();
 sg13g2_decap_8 FILLER_32_774 ();
 sg13g2_decap_8 FILLER_32_781 ();
 sg13g2_decap_8 FILLER_32_788 ();
 sg13g2_decap_8 FILLER_32_795 ();
 sg13g2_decap_8 FILLER_32_802 ();
 sg13g2_decap_8 FILLER_32_809 ();
 sg13g2_decap_8 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_823 ();
 sg13g2_decap_8 FILLER_32_830 ();
 sg13g2_decap_8 FILLER_32_837 ();
 sg13g2_decap_8 FILLER_32_844 ();
 sg13g2_decap_8 FILLER_32_851 ();
 sg13g2_decap_4 FILLER_32_858 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_4 ();
 sg13g2_decap_4 FILLER_33_45 ();
 sg13g2_decap_8 FILLER_33_66 ();
 sg13g2_decap_4 FILLER_33_73 ();
 sg13g2_fill_1 FILLER_33_77 ();
 sg13g2_fill_2 FILLER_33_87 ();
 sg13g2_decap_4 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_233 ();
 sg13g2_fill_1 FILLER_33_247 ();
 sg13g2_fill_2 FILLER_33_267 ();
 sg13g2_fill_2 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_344 ();
 sg13g2_fill_1 FILLER_33_346 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_decap_4 FILLER_33_414 ();
 sg13g2_fill_2 FILLER_33_418 ();
 sg13g2_decap_4 FILLER_33_458 ();
 sg13g2_decap_4 FILLER_33_490 ();
 sg13g2_fill_2 FILLER_33_494 ();
 sg13g2_decap_4 FILLER_33_514 ();
 sg13g2_fill_2 FILLER_33_518 ();
 sg13g2_decap_4 FILLER_33_533 ();
 sg13g2_fill_1 FILLER_33_537 ();
 sg13g2_fill_2 FILLER_33_547 ();
 sg13g2_fill_1 FILLER_33_549 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_fill_2 FILLER_33_631 ();
 sg13g2_fill_1 FILLER_33_688 ();
 sg13g2_fill_1 FILLER_33_699 ();
 sg13g2_decap_8 FILLER_33_736 ();
 sg13g2_decap_8 FILLER_33_743 ();
 sg13g2_decap_8 FILLER_33_750 ();
 sg13g2_decap_8 FILLER_33_757 ();
 sg13g2_decap_8 FILLER_33_764 ();
 sg13g2_decap_8 FILLER_33_771 ();
 sg13g2_decap_8 FILLER_33_778 ();
 sg13g2_decap_8 FILLER_33_785 ();
 sg13g2_decap_8 FILLER_33_792 ();
 sg13g2_decap_8 FILLER_33_799 ();
 sg13g2_decap_8 FILLER_33_806 ();
 sg13g2_decap_8 FILLER_33_813 ();
 sg13g2_decap_8 FILLER_33_820 ();
 sg13g2_decap_8 FILLER_33_827 ();
 sg13g2_decap_8 FILLER_33_834 ();
 sg13g2_decap_8 FILLER_33_841 ();
 sg13g2_decap_8 FILLER_33_848 ();
 sg13g2_decap_8 FILLER_33_855 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_18 ();
 sg13g2_fill_2 FILLER_34_28 ();
 sg13g2_decap_4 FILLER_34_62 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_fill_2 FILLER_34_152 ();
 sg13g2_decap_4 FILLER_34_181 ();
 sg13g2_fill_2 FILLER_34_185 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_204 ();
 sg13g2_fill_2 FILLER_34_231 ();
 sg13g2_fill_1 FILLER_34_298 ();
 sg13g2_fill_2 FILLER_34_304 ();
 sg13g2_fill_1 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_1 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_431 ();
 sg13g2_fill_2 FILLER_34_438 ();
 sg13g2_fill_2 FILLER_34_449 ();
 sg13g2_fill_1 FILLER_34_451 ();
 sg13g2_fill_1 FILLER_34_462 ();
 sg13g2_decap_4 FILLER_34_566 ();
 sg13g2_fill_1 FILLER_34_591 ();
 sg13g2_fill_1 FILLER_34_606 ();
 sg13g2_fill_1 FILLER_34_611 ();
 sg13g2_fill_2 FILLER_34_679 ();
 sg13g2_fill_1 FILLER_34_696 ();
 sg13g2_decap_8 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_740 ();
 sg13g2_decap_8 FILLER_34_747 ();
 sg13g2_decap_8 FILLER_34_754 ();
 sg13g2_decap_8 FILLER_34_761 ();
 sg13g2_decap_8 FILLER_34_768 ();
 sg13g2_decap_8 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_782 ();
 sg13g2_decap_8 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_796 ();
 sg13g2_decap_8 FILLER_34_803 ();
 sg13g2_decap_8 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_817 ();
 sg13g2_decap_8 FILLER_34_824 ();
 sg13g2_decap_8 FILLER_34_831 ();
 sg13g2_decap_8 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_fill_2 FILLER_34_859 ();
 sg13g2_fill_1 FILLER_34_861 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_30 ();
 sg13g2_fill_1 FILLER_35_32 ();
 sg13g2_decap_4 FILLER_35_42 ();
 sg13g2_fill_2 FILLER_35_46 ();
 sg13g2_decap_8 FILLER_35_58 ();
 sg13g2_fill_1 FILLER_35_65 ();
 sg13g2_fill_2 FILLER_35_103 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_fill_1 FILLER_35_130 ();
 sg13g2_fill_2 FILLER_35_140 ();
 sg13g2_fill_1 FILLER_35_197 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_1 FILLER_35_255 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_decap_4 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_fill_2 FILLER_35_350 ();
 sg13g2_fill_1 FILLER_35_352 ();
 sg13g2_fill_2 FILLER_35_358 ();
 sg13g2_fill_1 FILLER_35_360 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_1 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_fill_2 FILLER_35_436 ();
 sg13g2_fill_2 FILLER_35_460 ();
 sg13g2_fill_2 FILLER_35_494 ();
 sg13g2_fill_1 FILLER_35_496 ();
 sg13g2_fill_2 FILLER_35_511 ();
 sg13g2_fill_1 FILLER_35_513 ();
 sg13g2_fill_1 FILLER_35_523 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_4 FILLER_35_546 ();
 sg13g2_fill_1 FILLER_35_550 ();
 sg13g2_fill_2 FILLER_35_578 ();
 sg13g2_fill_2 FILLER_35_629 ();
 sg13g2_fill_2 FILLER_35_658 ();
 sg13g2_fill_1 FILLER_35_687 ();
 sg13g2_decap_4 FILLER_35_693 ();
 sg13g2_decap_4 FILLER_35_724 ();
 sg13g2_decap_8 FILLER_35_741 ();
 sg13g2_decap_8 FILLER_35_748 ();
 sg13g2_decap_8 FILLER_35_755 ();
 sg13g2_decap_8 FILLER_35_762 ();
 sg13g2_decap_8 FILLER_35_769 ();
 sg13g2_decap_8 FILLER_35_776 ();
 sg13g2_decap_8 FILLER_35_783 ();
 sg13g2_decap_8 FILLER_35_790 ();
 sg13g2_decap_8 FILLER_35_797 ();
 sg13g2_decap_8 FILLER_35_804 ();
 sg13g2_decap_8 FILLER_35_811 ();
 sg13g2_decap_8 FILLER_35_818 ();
 sg13g2_decap_8 FILLER_35_825 ();
 sg13g2_decap_8 FILLER_35_832 ();
 sg13g2_decap_8 FILLER_35_839 ();
 sg13g2_decap_8 FILLER_35_846 ();
 sg13g2_decap_8 FILLER_35_853 ();
 sg13g2_fill_2 FILLER_35_860 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_47 ();
 sg13g2_fill_1 FILLER_36_51 ();
 sg13g2_fill_2 FILLER_36_87 ();
 sg13g2_fill_2 FILLER_36_147 ();
 sg13g2_fill_1 FILLER_36_176 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_fill_1 FILLER_36_245 ();
 sg13g2_fill_2 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_296 ();
 sg13g2_fill_1 FILLER_36_298 ();
 sg13g2_decap_4 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_367 ();
 sg13g2_decap_4 FILLER_36_452 ();
 sg13g2_fill_2 FILLER_36_497 ();
 sg13g2_fill_1 FILLER_36_499 ();
 sg13g2_decap_4 FILLER_36_527 ();
 sg13g2_decap_8 FILLER_36_558 ();
 sg13g2_fill_1 FILLER_36_589 ();
 sg13g2_decap_4 FILLER_36_679 ();
 sg13g2_decap_8 FILLER_36_719 ();
 sg13g2_decap_8 FILLER_36_726 ();
 sg13g2_decap_8 FILLER_36_733 ();
 sg13g2_decap_8 FILLER_36_740 ();
 sg13g2_decap_8 FILLER_36_747 ();
 sg13g2_decap_8 FILLER_36_754 ();
 sg13g2_decap_8 FILLER_36_761 ();
 sg13g2_decap_8 FILLER_36_768 ();
 sg13g2_decap_8 FILLER_36_775 ();
 sg13g2_decap_8 FILLER_36_782 ();
 sg13g2_decap_8 FILLER_36_789 ();
 sg13g2_decap_8 FILLER_36_796 ();
 sg13g2_decap_8 FILLER_36_803 ();
 sg13g2_decap_8 FILLER_36_810 ();
 sg13g2_decap_8 FILLER_36_817 ();
 sg13g2_decap_8 FILLER_36_824 ();
 sg13g2_decap_8 FILLER_36_831 ();
 sg13g2_decap_8 FILLER_36_838 ();
 sg13g2_decap_8 FILLER_36_845 ();
 sg13g2_decap_8 FILLER_36_852 ();
 sg13g2_fill_2 FILLER_36_859 ();
 sg13g2_fill_1 FILLER_36_861 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_23 ();
 sg13g2_fill_1 FILLER_37_25 ();
 sg13g2_fill_2 FILLER_37_72 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_fill_2 FILLER_37_189 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_2 FILLER_37_301 ();
 sg13g2_fill_2 FILLER_37_331 ();
 sg13g2_decap_4 FILLER_37_343 ();
 sg13g2_fill_1 FILLER_37_347 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_fill_1 FILLER_37_363 ();
 sg13g2_decap_4 FILLER_37_377 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_8 FILLER_37_404 ();
 sg13g2_fill_2 FILLER_37_411 ();
 sg13g2_fill_2 FILLER_37_477 ();
 sg13g2_fill_1 FILLER_37_479 ();
 sg13g2_fill_2 FILLER_37_497 ();
 sg13g2_fill_1 FILLER_37_499 ();
 sg13g2_fill_2 FILLER_37_520 ();
 sg13g2_fill_1 FILLER_37_522 ();
 sg13g2_fill_1 FILLER_37_605 ();
 sg13g2_fill_1 FILLER_37_644 ();
 sg13g2_fill_2 FILLER_37_659 ();
 sg13g2_decap_8 FILLER_37_704 ();
 sg13g2_decap_8 FILLER_37_711 ();
 sg13g2_fill_1 FILLER_37_718 ();
 sg13g2_decap_8 FILLER_37_732 ();
 sg13g2_decap_8 FILLER_37_739 ();
 sg13g2_decap_8 FILLER_37_746 ();
 sg13g2_decap_8 FILLER_37_753 ();
 sg13g2_decap_8 FILLER_37_760 ();
 sg13g2_decap_8 FILLER_37_767 ();
 sg13g2_decap_8 FILLER_37_774 ();
 sg13g2_decap_8 FILLER_37_781 ();
 sg13g2_decap_8 FILLER_37_788 ();
 sg13g2_decap_8 FILLER_37_795 ();
 sg13g2_decap_8 FILLER_37_802 ();
 sg13g2_decap_8 FILLER_37_809 ();
 sg13g2_decap_8 FILLER_37_816 ();
 sg13g2_decap_8 FILLER_37_823 ();
 sg13g2_decap_8 FILLER_37_830 ();
 sg13g2_decap_8 FILLER_37_837 ();
 sg13g2_decap_8 FILLER_37_844 ();
 sg13g2_decap_8 FILLER_37_851 ();
 sg13g2_decap_4 FILLER_37_858 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_74 ();
 sg13g2_decap_8 FILLER_38_90 ();
 sg13g2_fill_1 FILLER_38_115 ();
 sg13g2_fill_2 FILLER_38_162 ();
 sg13g2_decap_4 FILLER_38_192 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_fill_2 FILLER_38_227 ();
 sg13g2_decap_4 FILLER_38_266 ();
 sg13g2_fill_1 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_fill_2 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_406 ();
 sg13g2_fill_2 FILLER_38_443 ();
 sg13g2_fill_2 FILLER_38_481 ();
 sg13g2_fill_1 FILLER_38_483 ();
 sg13g2_fill_2 FILLER_38_511 ();
 sg13g2_decap_4 FILLER_38_544 ();
 sg13g2_fill_2 FILLER_38_548 ();
 sg13g2_fill_1 FILLER_38_619 ();
 sg13g2_fill_2 FILLER_38_644 ();
 sg13g2_fill_1 FILLER_38_646 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_fill_1 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_46 ();
 sg13g2_fill_2 FILLER_39_50 ();
 sg13g2_fill_2 FILLER_39_79 ();
 sg13g2_fill_2 FILLER_39_136 ();
 sg13g2_decap_8 FILLER_39_174 ();
 sg13g2_fill_2 FILLER_39_181 ();
 sg13g2_fill_2 FILLER_39_202 ();
 sg13g2_decap_4 FILLER_39_246 ();
 sg13g2_decap_4 FILLER_39_296 ();
 sg13g2_fill_2 FILLER_39_310 ();
 sg13g2_decap_4 FILLER_39_325 ();
 sg13g2_fill_2 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_341 ();
 sg13g2_fill_2 FILLER_39_348 ();
 sg13g2_decap_4 FILLER_39_369 ();
 sg13g2_fill_1 FILLER_39_383 ();
 sg13g2_fill_1 FILLER_39_453 ();
 sg13g2_fill_1 FILLER_39_506 ();
 sg13g2_fill_2 FILLER_39_522 ();
 sg13g2_fill_1 FILLER_39_592 ();
 sg13g2_decap_8 FILLER_39_660 ();
 sg13g2_decap_8 FILLER_39_667 ();
 sg13g2_decap_8 FILLER_39_674 ();
 sg13g2_decap_8 FILLER_39_681 ();
 sg13g2_decap_8 FILLER_39_691 ();
 sg13g2_fill_1 FILLER_39_698 ();
 sg13g2_decap_8 FILLER_39_712 ();
 sg13g2_decap_8 FILLER_39_719 ();
 sg13g2_decap_8 FILLER_39_726 ();
 sg13g2_decap_8 FILLER_39_733 ();
 sg13g2_decap_8 FILLER_39_740 ();
 sg13g2_decap_8 FILLER_39_747 ();
 sg13g2_decap_8 FILLER_39_754 ();
 sg13g2_decap_8 FILLER_39_761 ();
 sg13g2_decap_8 FILLER_39_768 ();
 sg13g2_decap_8 FILLER_39_775 ();
 sg13g2_decap_8 FILLER_39_782 ();
 sg13g2_decap_8 FILLER_39_789 ();
 sg13g2_decap_8 FILLER_39_796 ();
 sg13g2_decap_8 FILLER_39_803 ();
 sg13g2_decap_8 FILLER_39_810 ();
 sg13g2_decap_8 FILLER_39_817 ();
 sg13g2_decap_8 FILLER_39_824 ();
 sg13g2_decap_8 FILLER_39_831 ();
 sg13g2_decap_8 FILLER_39_838 ();
 sg13g2_decap_8 FILLER_39_845 ();
 sg13g2_decap_8 FILLER_39_852 ();
 sg13g2_fill_2 FILLER_39_859 ();
 sg13g2_fill_1 FILLER_39_861 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_2 FILLER_40_4 ();
 sg13g2_decap_4 FILLER_40_45 ();
 sg13g2_decap_4 FILLER_40_59 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_fill_1 FILLER_40_168 ();
 sg13g2_fill_1 FILLER_40_208 ();
 sg13g2_decap_8 FILLER_40_222 ();
 sg13g2_fill_1 FILLER_40_243 ();
 sg13g2_decap_8 FILLER_40_257 ();
 sg13g2_decap_4 FILLER_40_264 ();
 sg13g2_decap_4 FILLER_40_306 ();
 sg13g2_fill_2 FILLER_40_366 ();
 sg13g2_decap_4 FILLER_40_373 ();
 sg13g2_fill_2 FILLER_40_377 ();
 sg13g2_decap_4 FILLER_40_388 ();
 sg13g2_fill_1 FILLER_40_392 ();
 sg13g2_fill_2 FILLER_40_452 ();
 sg13g2_fill_2 FILLER_40_473 ();
 sg13g2_fill_2 FILLER_40_484 ();
 sg13g2_fill_1 FILLER_40_514 ();
 sg13g2_fill_1 FILLER_40_546 ();
 sg13g2_decap_4 FILLER_40_585 ();
 sg13g2_fill_2 FILLER_40_589 ();
 sg13g2_decap_8 FILLER_40_617 ();
 sg13g2_decap_4 FILLER_40_647 ();
 sg13g2_fill_1 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_670 ();
 sg13g2_decap_8 FILLER_40_677 ();
 sg13g2_decap_8 FILLER_40_684 ();
 sg13g2_decap_8 FILLER_40_691 ();
 sg13g2_decap_8 FILLER_40_698 ();
 sg13g2_decap_8 FILLER_40_705 ();
 sg13g2_decap_8 FILLER_40_712 ();
 sg13g2_decap_8 FILLER_40_719 ();
 sg13g2_decap_8 FILLER_40_726 ();
 sg13g2_decap_8 FILLER_40_733 ();
 sg13g2_decap_8 FILLER_40_740 ();
 sg13g2_decap_8 FILLER_40_747 ();
 sg13g2_decap_8 FILLER_40_754 ();
 sg13g2_decap_8 FILLER_40_761 ();
 sg13g2_decap_8 FILLER_40_768 ();
 sg13g2_decap_8 FILLER_40_775 ();
 sg13g2_decap_8 FILLER_40_782 ();
 sg13g2_decap_8 FILLER_40_789 ();
 sg13g2_decap_8 FILLER_40_796 ();
 sg13g2_decap_8 FILLER_40_803 ();
 sg13g2_decap_8 FILLER_40_810 ();
 sg13g2_decap_8 FILLER_40_817 ();
 sg13g2_decap_8 FILLER_40_824 ();
 sg13g2_decap_8 FILLER_40_831 ();
 sg13g2_decap_8 FILLER_40_838 ();
 sg13g2_decap_8 FILLER_40_845 ();
 sg13g2_decap_8 FILLER_40_852 ();
 sg13g2_fill_2 FILLER_40_859 ();
 sg13g2_fill_1 FILLER_40_861 ();
 sg13g2_fill_1 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_29 ();
 sg13g2_fill_2 FILLER_41_111 ();
 sg13g2_decap_4 FILLER_41_130 ();
 sg13g2_fill_1 FILLER_41_134 ();
 sg13g2_decap_4 FILLER_41_174 ();
 sg13g2_fill_2 FILLER_41_192 ();
 sg13g2_decap_4 FILLER_41_222 ();
 sg13g2_decap_4 FILLER_41_244 ();
 sg13g2_fill_2 FILLER_41_248 ();
 sg13g2_fill_1 FILLER_41_259 ();
 sg13g2_fill_1 FILLER_41_275 ();
 sg13g2_fill_2 FILLER_41_285 ();
 sg13g2_decap_8 FILLER_41_296 ();
 sg13g2_fill_2 FILLER_41_303 ();
 sg13g2_fill_1 FILLER_41_305 ();
 sg13g2_fill_2 FILLER_41_317 ();
 sg13g2_fill_1 FILLER_41_319 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_fill_2 FILLER_41_343 ();
 sg13g2_fill_1 FILLER_41_345 ();
 sg13g2_fill_1 FILLER_41_483 ();
 sg13g2_fill_2 FILLER_41_520 ();
 sg13g2_fill_2 FILLER_41_544 ();
 sg13g2_fill_1 FILLER_41_564 ();
 sg13g2_fill_2 FILLER_41_579 ();
 sg13g2_fill_1 FILLER_41_635 ();
 sg13g2_decap_4 FILLER_41_646 ();
 sg13g2_decap_8 FILLER_41_677 ();
 sg13g2_fill_2 FILLER_41_684 ();
 sg13g2_fill_1 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_fill_1 FILLER_41_861 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_23 ();
 sg13g2_fill_2 FILLER_42_84 ();
 sg13g2_fill_2 FILLER_42_94 ();
 sg13g2_fill_1 FILLER_42_203 ();
 sg13g2_fill_1 FILLER_42_266 ();
 sg13g2_fill_1 FILLER_42_358 ();
 sg13g2_fill_2 FILLER_42_368 ();
 sg13g2_decap_8 FILLER_42_383 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_4 FILLER_42_397 ();
 sg13g2_fill_1 FILLER_42_401 ();
 sg13g2_fill_2 FILLER_42_419 ();
 sg13g2_fill_2 FILLER_42_434 ();
 sg13g2_fill_1 FILLER_42_436 ();
 sg13g2_fill_2 FILLER_42_446 ();
 sg13g2_fill_1 FILLER_42_470 ();
 sg13g2_fill_2 FILLER_42_483 ();
 sg13g2_fill_1 FILLER_42_485 ();
 sg13g2_fill_1 FILLER_42_495 ();
 sg13g2_fill_2 FILLER_42_532 ();
 sg13g2_fill_2 FILLER_42_598 ();
 sg13g2_fill_1 FILLER_42_600 ();
 sg13g2_fill_2 FILLER_42_615 ();
 sg13g2_decap_8 FILLER_42_627 ();
 sg13g2_fill_1 FILLER_42_634 ();
 sg13g2_decap_8 FILLER_42_692 ();
 sg13g2_decap_8 FILLER_42_699 ();
 sg13g2_decap_8 FILLER_42_706 ();
 sg13g2_decap_8 FILLER_42_713 ();
 sg13g2_decap_8 FILLER_42_720 ();
 sg13g2_decap_8 FILLER_42_727 ();
 sg13g2_decap_8 FILLER_42_734 ();
 sg13g2_decap_8 FILLER_42_741 ();
 sg13g2_decap_8 FILLER_42_748 ();
 sg13g2_decap_8 FILLER_42_755 ();
 sg13g2_decap_8 FILLER_42_762 ();
 sg13g2_decap_8 FILLER_42_769 ();
 sg13g2_decap_8 FILLER_42_776 ();
 sg13g2_decap_8 FILLER_42_783 ();
 sg13g2_decap_8 FILLER_42_790 ();
 sg13g2_decap_8 FILLER_42_797 ();
 sg13g2_decap_8 FILLER_42_804 ();
 sg13g2_decap_8 FILLER_42_811 ();
 sg13g2_decap_8 FILLER_42_818 ();
 sg13g2_decap_8 FILLER_42_825 ();
 sg13g2_decap_8 FILLER_42_832 ();
 sg13g2_decap_8 FILLER_42_839 ();
 sg13g2_decap_8 FILLER_42_846 ();
 sg13g2_decap_8 FILLER_42_853 ();
 sg13g2_fill_2 FILLER_42_860 ();
 sg13g2_fill_1 FILLER_43_40 ();
 sg13g2_fill_2 FILLER_43_54 ();
 sg13g2_fill_1 FILLER_43_56 ();
 sg13g2_fill_2 FILLER_43_84 ();
 sg13g2_fill_2 FILLER_43_91 ();
 sg13g2_fill_1 FILLER_43_147 ();
 sg13g2_fill_1 FILLER_43_157 ();
 sg13g2_fill_1 FILLER_43_167 ();
 sg13g2_decap_4 FILLER_43_182 ();
 sg13g2_decap_4 FILLER_43_195 ();
 sg13g2_fill_1 FILLER_43_199 ();
 sg13g2_fill_1 FILLER_43_245 ();
 sg13g2_decap_4 FILLER_43_253 ();
 sg13g2_fill_2 FILLER_43_257 ();
 sg13g2_decap_4 FILLER_43_281 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_fill_1 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_325 ();
 sg13g2_decap_4 FILLER_43_332 ();
 sg13g2_fill_2 FILLER_43_336 ();
 sg13g2_decap_4 FILLER_43_344 ();
 sg13g2_fill_1 FILLER_43_384 ();
 sg13g2_fill_1 FILLER_43_412 ();
 sg13g2_fill_2 FILLER_43_440 ();
 sg13g2_fill_2 FILLER_43_490 ();
 sg13g2_fill_1 FILLER_43_492 ();
 sg13g2_fill_1 FILLER_43_579 ();
 sg13g2_fill_2 FILLER_43_593 ();
 sg13g2_fill_1 FILLER_43_622 ();
 sg13g2_fill_2 FILLER_43_650 ();
 sg13g2_fill_1 FILLER_43_652 ();
 sg13g2_decap_8 FILLER_43_711 ();
 sg13g2_decap_8 FILLER_43_718 ();
 sg13g2_decap_8 FILLER_43_725 ();
 sg13g2_decap_8 FILLER_43_732 ();
 sg13g2_decap_8 FILLER_43_739 ();
 sg13g2_decap_8 FILLER_43_746 ();
 sg13g2_decap_8 FILLER_43_753 ();
 sg13g2_decap_8 FILLER_43_760 ();
 sg13g2_decap_8 FILLER_43_767 ();
 sg13g2_decap_8 FILLER_43_774 ();
 sg13g2_decap_8 FILLER_43_781 ();
 sg13g2_decap_8 FILLER_43_788 ();
 sg13g2_decap_8 FILLER_43_795 ();
 sg13g2_decap_8 FILLER_43_802 ();
 sg13g2_decap_8 FILLER_43_809 ();
 sg13g2_decap_8 FILLER_43_816 ();
 sg13g2_decap_8 FILLER_43_823 ();
 sg13g2_decap_8 FILLER_43_830 ();
 sg13g2_decap_8 FILLER_43_837 ();
 sg13g2_decap_8 FILLER_43_844 ();
 sg13g2_decap_8 FILLER_43_851 ();
 sg13g2_decap_4 FILLER_43_858 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_2 ();
 sg13g2_decap_4 FILLER_44_38 ();
 sg13g2_decap_8 FILLER_44_61 ();
 sg13g2_fill_1 FILLER_44_68 ();
 sg13g2_decap_4 FILLER_44_81 ();
 sg13g2_fill_1 FILLER_44_85 ();
 sg13g2_fill_1 FILLER_44_91 ();
 sg13g2_decap_8 FILLER_44_101 ();
 sg13g2_decap_8 FILLER_44_167 ();
 sg13g2_fill_2 FILLER_44_279 ();
 sg13g2_fill_1 FILLER_44_336 ();
 sg13g2_fill_2 FILLER_44_356 ();
 sg13g2_fill_1 FILLER_44_358 ();
 sg13g2_fill_2 FILLER_44_375 ();
 sg13g2_fill_2 FILLER_44_404 ();
 sg13g2_fill_1 FILLER_44_406 ();
 sg13g2_fill_1 FILLER_44_435 ();
 sg13g2_fill_1 FILLER_44_472 ();
 sg13g2_fill_1 FILLER_44_530 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_4 FILLER_44_638 ();
 sg13g2_fill_1 FILLER_44_642 ();
 sg13g2_fill_2 FILLER_44_678 ();
 sg13g2_fill_1 FILLER_44_680 ();
 sg13g2_decap_8 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_742 ();
 sg13g2_decap_8 FILLER_44_749 ();
 sg13g2_decap_8 FILLER_44_756 ();
 sg13g2_decap_8 FILLER_44_763 ();
 sg13g2_decap_8 FILLER_44_770 ();
 sg13g2_decap_8 FILLER_44_777 ();
 sg13g2_decap_8 FILLER_44_784 ();
 sg13g2_decap_8 FILLER_44_791 ();
 sg13g2_decap_8 FILLER_44_798 ();
 sg13g2_decap_8 FILLER_44_805 ();
 sg13g2_decap_8 FILLER_44_812 ();
 sg13g2_decap_8 FILLER_44_819 ();
 sg13g2_decap_8 FILLER_44_826 ();
 sg13g2_decap_8 FILLER_44_833 ();
 sg13g2_decap_8 FILLER_44_840 ();
 sg13g2_decap_8 FILLER_44_847 ();
 sg13g2_decap_8 FILLER_44_854 ();
 sg13g2_fill_1 FILLER_44_861 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_87 ();
 sg13g2_fill_1 FILLER_45_89 ();
 sg13g2_fill_2 FILLER_45_117 ();
 sg13g2_fill_1 FILLER_45_129 ();
 sg13g2_fill_2 FILLER_45_149 ();
 sg13g2_decap_4 FILLER_45_196 ();
 sg13g2_fill_1 FILLER_45_200 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_fill_1 FILLER_45_217 ();
 sg13g2_fill_2 FILLER_45_231 ();
 sg13g2_fill_2 FILLER_45_247 ();
 sg13g2_fill_1 FILLER_45_249 ();
 sg13g2_fill_2 FILLER_45_262 ();
 sg13g2_fill_1 FILLER_45_264 ();
 sg13g2_decap_8 FILLER_45_274 ();
 sg13g2_decap_8 FILLER_45_281 ();
 sg13g2_fill_2 FILLER_45_288 ();
 sg13g2_decap_8 FILLER_45_318 ();
 sg13g2_fill_2 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_4 FILLER_45_382 ();
 sg13g2_fill_1 FILLER_45_386 ();
 sg13g2_fill_1 FILLER_45_405 ();
 sg13g2_fill_2 FILLER_45_440 ();
 sg13g2_fill_1 FILLER_45_451 ();
 sg13g2_fill_2 FILLER_45_470 ();
 sg13g2_fill_2 FILLER_45_487 ();
 sg13g2_fill_1 FILLER_45_489 ();
 sg13g2_decap_4 FILLER_45_522 ();
 sg13g2_fill_2 FILLER_45_526 ();
 sg13g2_fill_1 FILLER_45_555 ();
 sg13g2_fill_2 FILLER_45_569 ();
 sg13g2_fill_1 FILLER_45_571 ();
 sg13g2_fill_2 FILLER_45_578 ();
 sg13g2_fill_1 FILLER_45_580 ();
 sg13g2_fill_2 FILLER_45_607 ();
 sg13g2_fill_2 FILLER_45_650 ();
 sg13g2_fill_1 FILLER_45_652 ();
 sg13g2_fill_1 FILLER_45_670 ();
 sg13g2_fill_2 FILLER_45_715 ();
 sg13g2_decap_8 FILLER_45_726 ();
 sg13g2_decap_8 FILLER_45_733 ();
 sg13g2_decap_8 FILLER_45_740 ();
 sg13g2_decap_8 FILLER_45_747 ();
 sg13g2_decap_8 FILLER_45_754 ();
 sg13g2_decap_8 FILLER_45_761 ();
 sg13g2_decap_8 FILLER_45_768 ();
 sg13g2_decap_8 FILLER_45_775 ();
 sg13g2_decap_8 FILLER_45_782 ();
 sg13g2_decap_8 FILLER_45_789 ();
 sg13g2_decap_8 FILLER_45_796 ();
 sg13g2_decap_8 FILLER_45_803 ();
 sg13g2_decap_8 FILLER_45_810 ();
 sg13g2_decap_8 FILLER_45_817 ();
 sg13g2_decap_8 FILLER_45_824 ();
 sg13g2_decap_8 FILLER_45_831 ();
 sg13g2_decap_8 FILLER_45_838 ();
 sg13g2_decap_8 FILLER_45_845 ();
 sg13g2_decap_8 FILLER_45_852 ();
 sg13g2_fill_2 FILLER_45_859 ();
 sg13g2_fill_1 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_fill_2 FILLER_46_11 ();
 sg13g2_decap_8 FILLER_46_32 ();
 sg13g2_decap_4 FILLER_46_52 ();
 sg13g2_decap_8 FILLER_46_66 ();
 sg13g2_fill_1 FILLER_46_73 ();
 sg13g2_decap_4 FILLER_46_106 ();
 sg13g2_fill_1 FILLER_46_110 ();
 sg13g2_fill_2 FILLER_46_152 ();
 sg13g2_decap_4 FILLER_46_185 ();
 sg13g2_fill_2 FILLER_46_189 ();
 sg13g2_decap_4 FILLER_46_219 ();
 sg13g2_fill_2 FILLER_46_238 ();
 sg13g2_fill_2 FILLER_46_264 ();
 sg13g2_decap_4 FILLER_46_279 ();
 sg13g2_decap_8 FILLER_46_352 ();
 sg13g2_decap_4 FILLER_46_359 ();
 sg13g2_fill_2 FILLER_46_363 ();
 sg13g2_decap_8 FILLER_46_380 ();
 sg13g2_fill_2 FILLER_46_387 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_fill_2 FILLER_46_412 ();
 sg13g2_fill_1 FILLER_46_414 ();
 sg13g2_fill_1 FILLER_46_421 ();
 sg13g2_fill_1 FILLER_46_434 ();
 sg13g2_decap_4 FILLER_46_508 ();
 sg13g2_fill_1 FILLER_46_512 ();
 sg13g2_fill_2 FILLER_46_540 ();
 sg13g2_fill_2 FILLER_46_565 ();
 sg13g2_fill_1 FILLER_46_567 ();
 sg13g2_fill_1 FILLER_46_590 ();
 sg13g2_fill_1 FILLER_46_622 ();
 sg13g2_fill_2 FILLER_46_678 ();
 sg13g2_fill_1 FILLER_46_680 ();
 sg13g2_fill_1 FILLER_46_694 ();
 sg13g2_decap_8 FILLER_46_732 ();
 sg13g2_decap_8 FILLER_46_739 ();
 sg13g2_decap_8 FILLER_46_746 ();
 sg13g2_decap_8 FILLER_46_753 ();
 sg13g2_decap_8 FILLER_46_760 ();
 sg13g2_decap_8 FILLER_46_767 ();
 sg13g2_decap_8 FILLER_46_774 ();
 sg13g2_decap_8 FILLER_46_781 ();
 sg13g2_decap_8 FILLER_46_788 ();
 sg13g2_decap_8 FILLER_46_795 ();
 sg13g2_decap_8 FILLER_46_802 ();
 sg13g2_decap_8 FILLER_46_809 ();
 sg13g2_decap_8 FILLER_46_816 ();
 sg13g2_decap_8 FILLER_46_823 ();
 sg13g2_decap_8 FILLER_46_830 ();
 sg13g2_decap_8 FILLER_46_837 ();
 sg13g2_decap_8 FILLER_46_844 ();
 sg13g2_decap_8 FILLER_46_851 ();
 sg13g2_decap_4 FILLER_46_858 ();
 sg13g2_fill_2 FILLER_47_27 ();
 sg13g2_fill_2 FILLER_47_56 ();
 sg13g2_fill_1 FILLER_47_58 ();
 sg13g2_fill_2 FILLER_47_86 ();
 sg13g2_fill_1 FILLER_47_88 ();
 sg13g2_fill_2 FILLER_47_119 ();
 sg13g2_decap_4 FILLER_47_193 ();
 sg13g2_fill_2 FILLER_47_197 ();
 sg13g2_fill_2 FILLER_47_259 ();
 sg13g2_fill_1 FILLER_47_261 ();
 sg13g2_fill_2 FILLER_47_286 ();
 sg13g2_decap_8 FILLER_47_298 ();
 sg13g2_decap_4 FILLER_47_324 ();
 sg13g2_fill_1 FILLER_47_328 ();
 sg13g2_decap_8 FILLER_47_366 ();
 sg13g2_fill_2 FILLER_47_397 ();
 sg13g2_fill_1 FILLER_47_399 ();
 sg13g2_fill_2 FILLER_47_410 ();
 sg13g2_fill_1 FILLER_47_418 ();
 sg13g2_fill_2 FILLER_47_425 ();
 sg13g2_fill_1 FILLER_47_462 ();
 sg13g2_fill_2 FILLER_47_508 ();
 sg13g2_fill_1 FILLER_47_556 ();
 sg13g2_fill_2 FILLER_47_590 ();
 sg13g2_decap_4 FILLER_47_603 ();
 sg13g2_fill_2 FILLER_47_616 ();
 sg13g2_fill_2 FILLER_47_632 ();
 sg13g2_fill_1 FILLER_47_677 ();
 sg13g2_fill_1 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_727 ();
 sg13g2_decap_8 FILLER_47_734 ();
 sg13g2_decap_8 FILLER_47_741 ();
 sg13g2_decap_8 FILLER_47_748 ();
 sg13g2_decap_8 FILLER_47_755 ();
 sg13g2_decap_8 FILLER_47_762 ();
 sg13g2_decap_8 FILLER_47_769 ();
 sg13g2_decap_8 FILLER_47_776 ();
 sg13g2_decap_8 FILLER_47_783 ();
 sg13g2_decap_8 FILLER_47_790 ();
 sg13g2_decap_8 FILLER_47_797 ();
 sg13g2_decap_8 FILLER_47_804 ();
 sg13g2_decap_8 FILLER_47_811 ();
 sg13g2_decap_8 FILLER_47_818 ();
 sg13g2_decap_8 FILLER_47_825 ();
 sg13g2_decap_8 FILLER_47_832 ();
 sg13g2_decap_8 FILLER_47_839 ();
 sg13g2_decap_8 FILLER_47_846 ();
 sg13g2_decap_8 FILLER_47_853 ();
 sg13g2_fill_2 FILLER_47_860 ();
 sg13g2_decap_4 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_4 ();
 sg13g2_decap_8 FILLER_48_32 ();
 sg13g2_fill_1 FILLER_48_39 ();
 sg13g2_fill_1 FILLER_48_69 ();
 sg13g2_fill_1 FILLER_48_98 ();
 sg13g2_fill_1 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_200 ();
 sg13g2_decap_4 FILLER_48_207 ();
 sg13g2_fill_2 FILLER_48_211 ();
 sg13g2_decap_4 FILLER_48_235 ();
 sg13g2_fill_1 FILLER_48_239 ();
 sg13g2_fill_2 FILLER_48_254 ();
 sg13g2_fill_1 FILLER_48_256 ();
 sg13g2_fill_1 FILLER_48_267 ();
 sg13g2_decap_8 FILLER_48_297 ();
 sg13g2_decap_4 FILLER_48_313 ();
 sg13g2_decap_8 FILLER_48_340 ();
 sg13g2_decap_4 FILLER_48_347 ();
 sg13g2_decap_8 FILLER_48_356 ();
 sg13g2_decap_8 FILLER_48_363 ();
 sg13g2_fill_1 FILLER_48_370 ();
 sg13g2_fill_2 FILLER_48_386 ();
 sg13g2_fill_1 FILLER_48_391 ();
 sg13g2_fill_1 FILLER_48_402 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_fill_1 FILLER_48_439 ();
 sg13g2_fill_1 FILLER_48_448 ();
 sg13g2_fill_2 FILLER_48_476 ();
 sg13g2_fill_2 FILLER_48_505 ();
 sg13g2_decap_8 FILLER_48_535 ();
 sg13g2_decap_8 FILLER_48_542 ();
 sg13g2_fill_2 FILLER_48_549 ();
 sg13g2_fill_1 FILLER_48_564 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_fill_2 FILLER_48_588 ();
 sg13g2_fill_2 FILLER_48_706 ();
 sg13g2_fill_1 FILLER_48_708 ();
 sg13g2_decap_8 FILLER_48_726 ();
 sg13g2_decap_8 FILLER_48_733 ();
 sg13g2_decap_8 FILLER_48_740 ();
 sg13g2_decap_8 FILLER_48_747 ();
 sg13g2_decap_8 FILLER_48_754 ();
 sg13g2_decap_8 FILLER_48_761 ();
 sg13g2_decap_8 FILLER_48_768 ();
 sg13g2_decap_8 FILLER_48_775 ();
 sg13g2_decap_8 FILLER_48_782 ();
 sg13g2_decap_8 FILLER_48_789 ();
 sg13g2_decap_8 FILLER_48_796 ();
 sg13g2_decap_8 FILLER_48_803 ();
 sg13g2_decap_8 FILLER_48_810 ();
 sg13g2_decap_8 FILLER_48_817 ();
 sg13g2_decap_8 FILLER_48_824 ();
 sg13g2_decap_8 FILLER_48_831 ();
 sg13g2_decap_8 FILLER_48_838 ();
 sg13g2_decap_8 FILLER_48_845 ();
 sg13g2_decap_8 FILLER_48_852 ();
 sg13g2_fill_2 FILLER_48_859 ();
 sg13g2_fill_1 FILLER_48_861 ();
 sg13g2_fill_2 FILLER_49_48 ();
 sg13g2_fill_1 FILLER_49_50 ();
 sg13g2_decap_4 FILLER_49_70 ();
 sg13g2_fill_2 FILLER_49_74 ();
 sg13g2_fill_1 FILLER_49_137 ();
 sg13g2_fill_2 FILLER_49_177 ();
 sg13g2_fill_1 FILLER_49_179 ();
 sg13g2_fill_2 FILLER_49_241 ();
 sg13g2_fill_1 FILLER_49_243 ();
 sg13g2_decap_4 FILLER_49_257 ();
 sg13g2_fill_1 FILLER_49_261 ();
 sg13g2_fill_2 FILLER_49_278 ();
 sg13g2_fill_1 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_390 ();
 sg13g2_fill_2 FILLER_49_397 ();
 sg13g2_fill_1 FILLER_49_399 ();
 sg13g2_decap_4 FILLER_49_409 ();
 sg13g2_fill_2 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_447 ();
 sg13g2_decap_8 FILLER_49_454 ();
 sg13g2_fill_2 FILLER_49_461 ();
 sg13g2_fill_1 FILLER_49_463 ();
 sg13g2_fill_2 FILLER_49_500 ();
 sg13g2_fill_1 FILLER_49_502 ();
 sg13g2_fill_2 FILLER_49_521 ();
 sg13g2_fill_1 FILLER_49_523 ();
 sg13g2_fill_1 FILLER_49_574 ();
 sg13g2_decap_4 FILLER_49_580 ();
 sg13g2_fill_1 FILLER_49_584 ();
 sg13g2_fill_1 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_642 ();
 sg13g2_fill_1 FILLER_49_649 ();
 sg13g2_fill_2 FILLER_49_672 ();
 sg13g2_fill_1 FILLER_49_674 ();
 sg13g2_fill_2 FILLER_49_706 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_fill_1 FILLER_49_861 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_29 ();
 sg13g2_fill_1 FILLER_50_36 ();
 sg13g2_decap_4 FILLER_50_64 ();
 sg13g2_fill_2 FILLER_50_95 ();
 sg13g2_fill_2 FILLER_50_110 ();
 sg13g2_fill_1 FILLER_50_121 ();
 sg13g2_fill_2 FILLER_50_135 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_2 FILLER_50_180 ();
 sg13g2_fill_1 FILLER_50_182 ();
 sg13g2_fill_1 FILLER_50_204 ();
 sg13g2_fill_1 FILLER_50_251 ();
 sg13g2_fill_2 FILLER_50_265 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_277 ();
 sg13g2_fill_2 FILLER_50_282 ();
 sg13g2_fill_1 FILLER_50_284 ();
 sg13g2_fill_2 FILLER_50_298 ();
 sg13g2_fill_1 FILLER_50_300 ();
 sg13g2_decap_4 FILLER_50_335 ();
 sg13g2_fill_2 FILLER_50_339 ();
 sg13g2_fill_2 FILLER_50_363 ();
 sg13g2_fill_1 FILLER_50_365 ();
 sg13g2_decap_4 FILLER_50_393 ();
 sg13g2_fill_1 FILLER_50_397 ();
 sg13g2_fill_2 FILLER_50_402 ();
 sg13g2_fill_1 FILLER_50_416 ();
 sg13g2_fill_1 FILLER_50_423 ();
 sg13g2_decap_8 FILLER_50_440 ();
 sg13g2_decap_4 FILLER_50_447 ();
 sg13g2_fill_2 FILLER_50_468 ();
 sg13g2_fill_1 FILLER_50_491 ();
 sg13g2_fill_2 FILLER_50_496 ();
 sg13g2_fill_1 FILLER_50_498 ();
 sg13g2_decap_8 FILLER_50_507 ();
 sg13g2_fill_1 FILLER_50_536 ();
 sg13g2_decap_8 FILLER_50_542 ();
 sg13g2_decap_4 FILLER_50_549 ();
 sg13g2_fill_2 FILLER_50_553 ();
 sg13g2_fill_1 FILLER_50_586 ();
 sg13g2_fill_1 FILLER_50_653 ();
 sg13g2_decap_8 FILLER_50_682 ();
 sg13g2_decap_4 FILLER_50_716 ();
 sg13g2_fill_1 FILLER_50_720 ();
 sg13g2_decap_8 FILLER_50_730 ();
 sg13g2_decap_8 FILLER_50_737 ();
 sg13g2_decap_8 FILLER_50_744 ();
 sg13g2_decap_8 FILLER_50_751 ();
 sg13g2_decap_8 FILLER_50_758 ();
 sg13g2_decap_8 FILLER_50_765 ();
 sg13g2_decap_8 FILLER_50_772 ();
 sg13g2_decap_8 FILLER_50_779 ();
 sg13g2_decap_8 FILLER_50_786 ();
 sg13g2_decap_8 FILLER_50_793 ();
 sg13g2_decap_8 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_807 ();
 sg13g2_decap_8 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_821 ();
 sg13g2_decap_8 FILLER_50_828 ();
 sg13g2_decap_8 FILLER_50_835 ();
 sg13g2_decap_8 FILLER_50_842 ();
 sg13g2_decap_8 FILLER_50_849 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_2 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_30 ();
 sg13g2_decap_8 FILLER_51_41 ();
 sg13g2_decap_8 FILLER_51_48 ();
 sg13g2_decap_4 FILLER_51_55 ();
 sg13g2_fill_1 FILLER_51_59 ();
 sg13g2_fill_1 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_105 ();
 sg13g2_fill_1 FILLER_51_107 ();
 sg13g2_fill_2 FILLER_51_189 ();
 sg13g2_fill_1 FILLER_51_191 ();
 sg13g2_decap_4 FILLER_51_235 ();
 sg13g2_decap_4 FILLER_51_248 ();
 sg13g2_decap_4 FILLER_51_269 ();
 sg13g2_fill_2 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_285 ();
 sg13g2_fill_2 FILLER_51_314 ();
 sg13g2_fill_1 FILLER_51_331 ();
 sg13g2_decap_8 FILLER_51_392 ();
 sg13g2_fill_2 FILLER_51_399 ();
 sg13g2_fill_1 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_412 ();
 sg13g2_decap_4 FILLER_51_438 ();
 sg13g2_fill_2 FILLER_51_442 ();
 sg13g2_decap_4 FILLER_51_448 ();
 sg13g2_fill_2 FILLER_51_452 ();
 sg13g2_decap_8 FILLER_51_476 ();
 sg13g2_decap_4 FILLER_51_532 ();
 sg13g2_fill_2 FILLER_51_554 ();
 sg13g2_decap_8 FILLER_51_561 ();
 sg13g2_decap_4 FILLER_51_568 ();
 sg13g2_decap_4 FILLER_51_577 ();
 sg13g2_fill_2 FILLER_51_586 ();
 sg13g2_fill_1 FILLER_51_611 ();
 sg13g2_decap_8 FILLER_51_636 ();
 sg13g2_fill_1 FILLER_51_706 ();
 sg13g2_decap_8 FILLER_51_734 ();
 sg13g2_decap_8 FILLER_51_741 ();
 sg13g2_decap_8 FILLER_51_748 ();
 sg13g2_decap_8 FILLER_51_755 ();
 sg13g2_decap_8 FILLER_51_762 ();
 sg13g2_decap_8 FILLER_51_769 ();
 sg13g2_decap_8 FILLER_51_776 ();
 sg13g2_decap_8 FILLER_51_783 ();
 sg13g2_decap_8 FILLER_51_790 ();
 sg13g2_decap_8 FILLER_51_797 ();
 sg13g2_decap_8 FILLER_51_804 ();
 sg13g2_decap_8 FILLER_51_811 ();
 sg13g2_decap_8 FILLER_51_818 ();
 sg13g2_decap_8 FILLER_51_825 ();
 sg13g2_decap_8 FILLER_51_832 ();
 sg13g2_decap_8 FILLER_51_839 ();
 sg13g2_decap_8 FILLER_51_846 ();
 sg13g2_decap_8 FILLER_51_853 ();
 sg13g2_fill_2 FILLER_51_860 ();
 sg13g2_decap_4 FILLER_52_36 ();
 sg13g2_fill_2 FILLER_52_40 ();
 sg13g2_fill_2 FILLER_52_52 ();
 sg13g2_fill_1 FILLER_52_97 ();
 sg13g2_fill_2 FILLER_52_117 ();
 sg13g2_fill_2 FILLER_52_218 ();
 sg13g2_fill_1 FILLER_52_253 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_fill_2 FILLER_52_266 ();
 sg13g2_fill_1 FILLER_52_268 ();
 sg13g2_fill_1 FILLER_52_288 ();
 sg13g2_fill_1 FILLER_52_311 ();
 sg13g2_fill_1 FILLER_52_320 ();
 sg13g2_fill_2 FILLER_52_330 ();
 sg13g2_fill_1 FILLER_52_332 ();
 sg13g2_fill_2 FILLER_52_346 ();
 sg13g2_fill_1 FILLER_52_348 ();
 sg13g2_decap_4 FILLER_52_380 ();
 sg13g2_fill_2 FILLER_52_412 ();
 sg13g2_fill_1 FILLER_52_414 ();
 sg13g2_fill_1 FILLER_52_421 ();
 sg13g2_decap_8 FILLER_52_431 ();
 sg13g2_fill_2 FILLER_52_438 ();
 sg13g2_decap_4 FILLER_52_478 ();
 sg13g2_fill_1 FILLER_52_482 ();
 sg13g2_decap_8 FILLER_52_503 ();
 sg13g2_decap_8 FILLER_52_510 ();
 sg13g2_fill_2 FILLER_52_517 ();
 sg13g2_fill_1 FILLER_52_542 ();
 sg13g2_fill_2 FILLER_52_552 ();
 sg13g2_fill_1 FILLER_52_572 ();
 sg13g2_fill_2 FILLER_52_587 ();
 sg13g2_fill_1 FILLER_52_589 ();
 sg13g2_fill_2 FILLER_52_616 ();
 sg13g2_fill_1 FILLER_52_618 ();
 sg13g2_fill_2 FILLER_52_625 ();
 sg13g2_decap_8 FILLER_52_632 ();
 sg13g2_decap_4 FILLER_52_649 ();
 sg13g2_fill_1 FILLER_52_653 ();
 sg13g2_decap_4 FILLER_52_663 ();
 sg13g2_fill_1 FILLER_52_667 ();
 sg13g2_decap_4 FILLER_52_714 ();
 sg13g2_fill_1 FILLER_52_718 ();
 sg13g2_decap_8 FILLER_52_728 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_decap_8 FILLER_52_742 ();
 sg13g2_decap_8 FILLER_52_749 ();
 sg13g2_decap_8 FILLER_52_756 ();
 sg13g2_decap_8 FILLER_52_763 ();
 sg13g2_decap_8 FILLER_52_770 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_decap_8 FILLER_52_791 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_fill_1 FILLER_52_861 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_47 ();
 sg13g2_fill_2 FILLER_53_58 ();
 sg13g2_fill_2 FILLER_53_96 ();
 sg13g2_fill_2 FILLER_53_103 ();
 sg13g2_fill_1 FILLER_53_142 ();
 sg13g2_fill_1 FILLER_53_186 ();
 sg13g2_fill_1 FILLER_53_205 ();
 sg13g2_decap_8 FILLER_53_215 ();
 sg13g2_decap_4 FILLER_53_222 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_8 FILLER_53_254 ();
 sg13g2_decap_4 FILLER_53_261 ();
 sg13g2_fill_2 FILLER_53_265 ();
 sg13g2_fill_2 FILLER_53_339 ();
 sg13g2_decap_4 FILLER_53_380 ();
 sg13g2_fill_2 FILLER_53_384 ();
 sg13g2_decap_4 FILLER_53_414 ();
 sg13g2_fill_1 FILLER_53_418 ();
 sg13g2_fill_2 FILLER_53_456 ();
 sg13g2_fill_2 FILLER_53_486 ();
 sg13g2_decap_4 FILLER_53_496 ();
 sg13g2_fill_1 FILLER_53_500 ();
 sg13g2_fill_2 FILLER_53_519 ();
 sg13g2_decap_8 FILLER_53_531 ();
 sg13g2_fill_2 FILLER_53_538 ();
 sg13g2_fill_1 FILLER_53_540 ();
 sg13g2_decap_8 FILLER_53_598 ();
 sg13g2_fill_1 FILLER_53_605 ();
 sg13g2_fill_2 FILLER_53_634 ();
 sg13g2_fill_2 FILLER_53_646 ();
 sg13g2_fill_1 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_728 ();
 sg13g2_decap_8 FILLER_53_735 ();
 sg13g2_decap_8 FILLER_53_742 ();
 sg13g2_decap_8 FILLER_53_749 ();
 sg13g2_decap_8 FILLER_53_756 ();
 sg13g2_decap_8 FILLER_53_763 ();
 sg13g2_decap_8 FILLER_53_770 ();
 sg13g2_decap_8 FILLER_53_777 ();
 sg13g2_decap_8 FILLER_53_784 ();
 sg13g2_decap_8 FILLER_53_791 ();
 sg13g2_decap_8 FILLER_53_798 ();
 sg13g2_decap_8 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_812 ();
 sg13g2_decap_8 FILLER_53_819 ();
 sg13g2_decap_8 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_833 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_53_847 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_fill_1 FILLER_53_861 ();
 sg13g2_fill_2 FILLER_54_66 ();
 sg13g2_fill_2 FILLER_54_103 ();
 sg13g2_fill_1 FILLER_54_105 ();
 sg13g2_fill_2 FILLER_54_143 ();
 sg13g2_fill_1 FILLER_54_145 ();
 sg13g2_fill_2 FILLER_54_224 ();
 sg13g2_fill_1 FILLER_54_267 ();
 sg13g2_decap_8 FILLER_54_282 ();
 sg13g2_fill_2 FILLER_54_289 ();
 sg13g2_fill_2 FILLER_54_311 ();
 sg13g2_fill_1 FILLER_54_313 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_decap_8 FILLER_54_403 ();
 sg13g2_decap_8 FILLER_54_410 ();
 sg13g2_fill_1 FILLER_54_432 ();
 sg13g2_decap_4 FILLER_54_437 ();
 sg13g2_decap_8 FILLER_54_459 ();
 sg13g2_decap_8 FILLER_54_466 ();
 sg13g2_decap_8 FILLER_54_473 ();
 sg13g2_fill_2 FILLER_54_480 ();
 sg13g2_decap_8 FILLER_54_487 ();
 sg13g2_decap_4 FILLER_54_494 ();
 sg13g2_fill_2 FILLER_54_498 ();
 sg13g2_decap_4 FILLER_54_513 ();
 sg13g2_fill_1 FILLER_54_517 ();
 sg13g2_decap_4 FILLER_54_541 ();
 sg13g2_fill_2 FILLER_54_545 ();
 sg13g2_decap_8 FILLER_54_555 ();
 sg13g2_decap_8 FILLER_54_570 ();
 sg13g2_fill_1 FILLER_54_577 ();
 sg13g2_decap_4 FILLER_54_587 ();
 sg13g2_fill_2 FILLER_54_591 ();
 sg13g2_decap_8 FILLER_54_613 ();
 sg13g2_fill_1 FILLER_54_626 ();
 sg13g2_decap_8 FILLER_54_632 ();
 sg13g2_fill_2 FILLER_54_680 ();
 sg13g2_fill_1 FILLER_54_682 ();
 sg13g2_fill_1 FILLER_54_714 ();
 sg13g2_decap_8 FILLER_54_732 ();
 sg13g2_decap_8 FILLER_54_739 ();
 sg13g2_decap_8 FILLER_54_746 ();
 sg13g2_decap_8 FILLER_54_753 ();
 sg13g2_decap_8 FILLER_54_760 ();
 sg13g2_decap_8 FILLER_54_767 ();
 sg13g2_decap_8 FILLER_54_774 ();
 sg13g2_decap_8 FILLER_54_781 ();
 sg13g2_decap_8 FILLER_54_788 ();
 sg13g2_decap_8 FILLER_54_795 ();
 sg13g2_decap_8 FILLER_54_802 ();
 sg13g2_decap_8 FILLER_54_809 ();
 sg13g2_decap_8 FILLER_54_816 ();
 sg13g2_decap_8 FILLER_54_823 ();
 sg13g2_decap_8 FILLER_54_830 ();
 sg13g2_decap_8 FILLER_54_837 ();
 sg13g2_decap_8 FILLER_54_844 ();
 sg13g2_decap_8 FILLER_54_851 ();
 sg13g2_decap_4 FILLER_54_858 ();
 sg13g2_fill_2 FILLER_55_34 ();
 sg13g2_fill_1 FILLER_55_62 ();
 sg13g2_fill_2 FILLER_55_184 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_fill_2 FILLER_55_238 ();
 sg13g2_fill_1 FILLER_55_240 ();
 sg13g2_fill_2 FILLER_55_270 ();
 sg13g2_fill_1 FILLER_55_322 ();
 sg13g2_fill_1 FILLER_55_332 ();
 sg13g2_fill_1 FILLER_55_344 ();
 sg13g2_decap_8 FILLER_55_358 ();
 sg13g2_decap_8 FILLER_55_365 ();
 sg13g2_fill_1 FILLER_55_372 ();
 sg13g2_decap_4 FILLER_55_401 ();
 sg13g2_fill_2 FILLER_55_462 ();
 sg13g2_fill_2 FILLER_55_528 ();
 sg13g2_decap_8 FILLER_55_542 ();
 sg13g2_fill_1 FILLER_55_549 ();
 sg13g2_fill_1 FILLER_55_560 ();
 sg13g2_decap_4 FILLER_55_566 ();
 sg13g2_fill_1 FILLER_55_579 ();
 sg13g2_fill_1 FILLER_55_597 ();
 sg13g2_fill_1 FILLER_55_691 ();
 sg13g2_decap_8 FILLER_55_723 ();
 sg13g2_decap_8 FILLER_55_730 ();
 sg13g2_decap_8 FILLER_55_737 ();
 sg13g2_decap_8 FILLER_55_744 ();
 sg13g2_decap_8 FILLER_55_751 ();
 sg13g2_decap_8 FILLER_55_758 ();
 sg13g2_decap_8 FILLER_55_765 ();
 sg13g2_decap_8 FILLER_55_772 ();
 sg13g2_decap_8 FILLER_55_779 ();
 sg13g2_decap_8 FILLER_55_786 ();
 sg13g2_decap_8 FILLER_55_793 ();
 sg13g2_decap_8 FILLER_55_800 ();
 sg13g2_decap_8 FILLER_55_807 ();
 sg13g2_decap_8 FILLER_55_814 ();
 sg13g2_decap_8 FILLER_55_821 ();
 sg13g2_decap_8 FILLER_55_828 ();
 sg13g2_decap_8 FILLER_55_835 ();
 sg13g2_decap_8 FILLER_55_842 ();
 sg13g2_decap_8 FILLER_55_849 ();
 sg13g2_decap_4 FILLER_55_856 ();
 sg13g2_fill_2 FILLER_55_860 ();
 sg13g2_fill_1 FILLER_56_18 ();
 sg13g2_fill_2 FILLER_56_45 ();
 sg13g2_fill_1 FILLER_56_78 ();
 sg13g2_fill_1 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_102 ();
 sg13g2_fill_1 FILLER_56_134 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_fill_1 FILLER_56_155 ();
 sg13g2_fill_1 FILLER_56_169 ();
 sg13g2_fill_1 FILLER_56_183 ();
 sg13g2_decap_4 FILLER_56_224 ();
 sg13g2_fill_1 FILLER_56_228 ();
 sg13g2_decap_8 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_377 ();
 sg13g2_fill_2 FILLER_56_423 ();
 sg13g2_fill_1 FILLER_56_425 ();
 sg13g2_decap_4 FILLER_56_452 ();
 sg13g2_fill_1 FILLER_56_495 ();
 sg13g2_fill_1 FILLER_56_509 ();
 sg13g2_fill_2 FILLER_56_553 ();
 sg13g2_fill_1 FILLER_56_555 ();
 sg13g2_decap_8 FILLER_56_590 ();
 sg13g2_decap_8 FILLER_56_597 ();
 sg13g2_decap_8 FILLER_56_604 ();
 sg13g2_fill_1 FILLER_56_611 ();
 sg13g2_decap_8 FILLER_56_627 ();
 sg13g2_decap_8 FILLER_56_634 ();
 sg13g2_decap_4 FILLER_56_641 ();
 sg13g2_fill_2 FILLER_56_645 ();
 sg13g2_fill_1 FILLER_56_701 ();
 sg13g2_decap_8 FILLER_56_723 ();
 sg13g2_decap_8 FILLER_56_730 ();
 sg13g2_decap_8 FILLER_56_737 ();
 sg13g2_decap_8 FILLER_56_744 ();
 sg13g2_decap_8 FILLER_56_751 ();
 sg13g2_decap_8 FILLER_56_758 ();
 sg13g2_decap_8 FILLER_56_765 ();
 sg13g2_decap_8 FILLER_56_772 ();
 sg13g2_decap_8 FILLER_56_779 ();
 sg13g2_decap_8 FILLER_56_786 ();
 sg13g2_decap_8 FILLER_56_793 ();
 sg13g2_decap_8 FILLER_56_800 ();
 sg13g2_decap_8 FILLER_56_807 ();
 sg13g2_decap_8 FILLER_56_814 ();
 sg13g2_decap_8 FILLER_56_821 ();
 sg13g2_decap_8 FILLER_56_828 ();
 sg13g2_decap_8 FILLER_56_835 ();
 sg13g2_decap_8 FILLER_56_842 ();
 sg13g2_decap_8 FILLER_56_849 ();
 sg13g2_decap_4 FILLER_56_856 ();
 sg13g2_fill_2 FILLER_56_860 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_49 ();
 sg13g2_fill_1 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_119 ();
 sg13g2_fill_2 FILLER_57_138 ();
 sg13g2_fill_2 FILLER_57_167 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_fill_1 FILLER_57_204 ();
 sg13g2_fill_1 FILLER_57_232 ();
 sg13g2_decap_4 FILLER_57_259 ();
 sg13g2_fill_1 FILLER_57_263 ();
 sg13g2_fill_1 FILLER_57_273 ();
 sg13g2_fill_2 FILLER_57_366 ();
 sg13g2_fill_1 FILLER_57_368 ();
 sg13g2_fill_1 FILLER_57_409 ();
 sg13g2_fill_1 FILLER_57_419 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_57_505 ();
 sg13g2_decap_8 FILLER_57_512 ();
 sg13g2_fill_2 FILLER_57_519 ();
 sg13g2_decap_8 FILLER_57_530 ();
 sg13g2_fill_2 FILLER_57_547 ();
 sg13g2_fill_1 FILLER_57_549 ();
 sg13g2_fill_1 FILLER_57_569 ();
 sg13g2_fill_2 FILLER_57_604 ();
 sg13g2_fill_2 FILLER_57_661 ();
 sg13g2_fill_1 FILLER_57_663 ();
 sg13g2_decap_8 FILLER_57_718 ();
 sg13g2_decap_8 FILLER_57_725 ();
 sg13g2_decap_8 FILLER_57_732 ();
 sg13g2_decap_8 FILLER_57_739 ();
 sg13g2_decap_8 FILLER_57_746 ();
 sg13g2_decap_8 FILLER_57_753 ();
 sg13g2_decap_8 FILLER_57_760 ();
 sg13g2_decap_8 FILLER_57_767 ();
 sg13g2_decap_8 FILLER_57_774 ();
 sg13g2_decap_8 FILLER_57_781 ();
 sg13g2_decap_8 FILLER_57_788 ();
 sg13g2_decap_8 FILLER_57_795 ();
 sg13g2_decap_8 FILLER_57_802 ();
 sg13g2_decap_8 FILLER_57_809 ();
 sg13g2_decap_8 FILLER_57_816 ();
 sg13g2_decap_8 FILLER_57_823 ();
 sg13g2_decap_8 FILLER_57_830 ();
 sg13g2_decap_8 FILLER_57_837 ();
 sg13g2_decap_8 FILLER_57_844 ();
 sg13g2_decap_8 FILLER_57_851 ();
 sg13g2_decap_4 FILLER_57_858 ();
 sg13g2_fill_2 FILLER_58_45 ();
 sg13g2_fill_2 FILLER_58_57 ();
 sg13g2_fill_2 FILLER_58_82 ();
 sg13g2_fill_1 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_126 ();
 sg13g2_fill_1 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_181 ();
 sg13g2_decap_8 FILLER_58_234 ();
 sg13g2_decap_4 FILLER_58_241 ();
 sg13g2_fill_1 FILLER_58_245 ();
 sg13g2_decap_4 FILLER_58_273 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_345 ();
 sg13g2_fill_1 FILLER_58_407 ();
 sg13g2_fill_1 FILLER_58_440 ();
 sg13g2_fill_1 FILLER_58_513 ();
 sg13g2_fill_1 FILLER_58_526 ();
 sg13g2_fill_2 FILLER_58_532 ();
 sg13g2_fill_1 FILLER_58_534 ();
 sg13g2_fill_1 FILLER_58_539 ();
 sg13g2_fill_2 FILLER_58_551 ();
 sg13g2_fill_1 FILLER_58_553 ();
 sg13g2_decap_8 FILLER_58_573 ();
 sg13g2_decap_8 FILLER_58_589 ();
 sg13g2_fill_2 FILLER_58_596 ();
 sg13g2_fill_1 FILLER_58_606 ();
 sg13g2_fill_1 FILLER_58_633 ();
 sg13g2_fill_1 FILLER_58_690 ();
 sg13g2_fill_2 FILLER_58_704 ();
 sg13g2_fill_1 FILLER_58_706 ();
 sg13g2_decap_8 FILLER_58_716 ();
 sg13g2_decap_8 FILLER_58_723 ();
 sg13g2_decap_8 FILLER_58_730 ();
 sg13g2_decap_8 FILLER_58_737 ();
 sg13g2_decap_8 FILLER_58_744 ();
 sg13g2_decap_8 FILLER_58_751 ();
 sg13g2_decap_8 FILLER_58_758 ();
 sg13g2_decap_8 FILLER_58_765 ();
 sg13g2_decap_8 FILLER_58_772 ();
 sg13g2_decap_8 FILLER_58_779 ();
 sg13g2_decap_8 FILLER_58_786 ();
 sg13g2_decap_8 FILLER_58_793 ();
 sg13g2_decap_8 FILLER_58_800 ();
 sg13g2_decap_8 FILLER_58_807 ();
 sg13g2_decap_8 FILLER_58_814 ();
 sg13g2_decap_8 FILLER_58_821 ();
 sg13g2_decap_8 FILLER_58_828 ();
 sg13g2_decap_8 FILLER_58_835 ();
 sg13g2_decap_8 FILLER_58_842 ();
 sg13g2_decap_8 FILLER_58_849 ();
 sg13g2_decap_4 FILLER_58_856 ();
 sg13g2_fill_2 FILLER_58_860 ();
 sg13g2_fill_1 FILLER_59_49 ();
 sg13g2_fill_2 FILLER_59_85 ();
 sg13g2_fill_2 FILLER_59_142 ();
 sg13g2_fill_1 FILLER_59_144 ();
 sg13g2_fill_2 FILLER_59_226 ();
 sg13g2_fill_1 FILLER_59_228 ();
 sg13g2_decap_8 FILLER_59_257 ();
 sg13g2_fill_2 FILLER_59_291 ();
 sg13g2_fill_1 FILLER_59_293 ();
 sg13g2_fill_1 FILLER_59_353 ();
 sg13g2_fill_2 FILLER_59_363 ();
 sg13g2_fill_1 FILLER_59_365 ();
 sg13g2_fill_1 FILLER_59_377 ();
 sg13g2_fill_2 FILLER_59_445 ();
 sg13g2_fill_2 FILLER_59_479 ();
 sg13g2_fill_2 FILLER_59_509 ();
 sg13g2_fill_1 FILLER_59_540 ();
 sg13g2_fill_1 FILLER_59_686 ();
 sg13g2_decap_8 FILLER_59_701 ();
 sg13g2_decap_8 FILLER_59_708 ();
 sg13g2_decap_8 FILLER_59_715 ();
 sg13g2_decap_8 FILLER_59_722 ();
 sg13g2_decap_8 FILLER_59_729 ();
 sg13g2_decap_8 FILLER_59_736 ();
 sg13g2_decap_8 FILLER_59_743 ();
 sg13g2_decap_8 FILLER_59_750 ();
 sg13g2_decap_8 FILLER_59_757 ();
 sg13g2_decap_8 FILLER_59_764 ();
 sg13g2_decap_8 FILLER_59_771 ();
 sg13g2_decap_8 FILLER_59_778 ();
 sg13g2_decap_8 FILLER_59_785 ();
 sg13g2_decap_8 FILLER_59_792 ();
 sg13g2_decap_8 FILLER_59_799 ();
 sg13g2_decap_8 FILLER_59_806 ();
 sg13g2_decap_8 FILLER_59_813 ();
 sg13g2_decap_8 FILLER_59_820 ();
 sg13g2_decap_8 FILLER_59_827 ();
 sg13g2_decap_8 FILLER_59_834 ();
 sg13g2_decap_8 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_fill_1 FILLER_60_40 ();
 sg13g2_fill_2 FILLER_60_85 ();
 sg13g2_fill_1 FILLER_60_87 ();
 sg13g2_fill_2 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_164 ();
 sg13g2_fill_1 FILLER_60_189 ();
 sg13g2_decap_8 FILLER_60_245 ();
 sg13g2_decap_4 FILLER_60_252 ();
 sg13g2_fill_1 FILLER_60_256 ();
 sg13g2_fill_2 FILLER_60_267 ();
 sg13g2_fill_1 FILLER_60_278 ();
 sg13g2_fill_1 FILLER_60_288 ();
 sg13g2_fill_1 FILLER_60_344 ();
 sg13g2_fill_2 FILLER_60_381 ();
 sg13g2_fill_2 FILLER_60_388 ();
 sg13g2_fill_2 FILLER_60_426 ();
 sg13g2_decap_4 FILLER_60_504 ();
 sg13g2_fill_1 FILLER_60_508 ();
 sg13g2_fill_1 FILLER_60_517 ();
 sg13g2_fill_1 FILLER_60_532 ();
 sg13g2_decap_4 FILLER_60_542 ();
 sg13g2_fill_2 FILLER_60_560 ();
 sg13g2_decap_8 FILLER_60_593 ();
 sg13g2_fill_1 FILLER_60_672 ();
 sg13g2_fill_1 FILLER_60_679 ();
 sg13g2_decap_8 FILLER_60_708 ();
 sg13g2_decap_8 FILLER_60_715 ();
 sg13g2_decap_8 FILLER_60_722 ();
 sg13g2_decap_8 FILLER_60_729 ();
 sg13g2_decap_8 FILLER_60_736 ();
 sg13g2_decap_8 FILLER_60_743 ();
 sg13g2_decap_8 FILLER_60_750 ();
 sg13g2_decap_8 FILLER_60_757 ();
 sg13g2_decap_8 FILLER_60_764 ();
 sg13g2_decap_8 FILLER_60_771 ();
 sg13g2_decap_8 FILLER_60_778 ();
 sg13g2_decap_8 FILLER_60_785 ();
 sg13g2_decap_8 FILLER_60_792 ();
 sg13g2_decap_8 FILLER_60_799 ();
 sg13g2_decap_8 FILLER_60_806 ();
 sg13g2_decap_8 FILLER_60_813 ();
 sg13g2_decap_8 FILLER_60_820 ();
 sg13g2_decap_8 FILLER_60_827 ();
 sg13g2_decap_8 FILLER_60_834 ();
 sg13g2_decap_8 FILLER_60_841 ();
 sg13g2_decap_8 FILLER_60_848 ();
 sg13g2_decap_8 FILLER_60_855 ();
 sg13g2_fill_1 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_141 ();
 sg13g2_fill_2 FILLER_61_198 ();
 sg13g2_fill_1 FILLER_61_200 ();
 sg13g2_fill_2 FILLER_61_319 ();
 sg13g2_fill_2 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_fill_1 FILLER_61_452 ();
 sg13g2_fill_2 FILLER_61_512 ();
 sg13g2_fill_1 FILLER_61_514 ();
 sg13g2_fill_2 FILLER_61_554 ();
 sg13g2_decap_4 FILLER_61_569 ();
 sg13g2_fill_1 FILLER_61_573 ();
 sg13g2_fill_1 FILLER_61_581 ();
 sg13g2_decap_8 FILLER_61_590 ();
 sg13g2_fill_1 FILLER_61_597 ();
 sg13g2_fill_2 FILLER_61_632 ();
 sg13g2_fill_1 FILLER_61_701 ();
 sg13g2_decap_8 FILLER_61_730 ();
 sg13g2_decap_8 FILLER_61_737 ();
 sg13g2_decap_8 FILLER_61_744 ();
 sg13g2_decap_8 FILLER_61_751 ();
 sg13g2_decap_8 FILLER_61_758 ();
 sg13g2_decap_8 FILLER_61_765 ();
 sg13g2_decap_8 FILLER_61_772 ();
 sg13g2_decap_8 FILLER_61_779 ();
 sg13g2_decap_8 FILLER_61_786 ();
 sg13g2_decap_8 FILLER_61_793 ();
 sg13g2_decap_8 FILLER_61_800 ();
 sg13g2_decap_8 FILLER_61_807 ();
 sg13g2_decap_8 FILLER_61_814 ();
 sg13g2_decap_8 FILLER_61_821 ();
 sg13g2_decap_8 FILLER_61_828 ();
 sg13g2_decap_8 FILLER_61_835 ();
 sg13g2_decap_8 FILLER_61_842 ();
 sg13g2_decap_8 FILLER_61_849 ();
 sg13g2_decap_4 FILLER_61_856 ();
 sg13g2_fill_2 FILLER_61_860 ();
 sg13g2_fill_1 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_161 ();
 sg13g2_fill_2 FILLER_62_191 ();
 sg13g2_fill_1 FILLER_62_193 ();
 sg13g2_fill_1 FILLER_62_228 ();
 sg13g2_fill_2 FILLER_62_242 ();
 sg13g2_fill_2 FILLER_62_253 ();
 sg13g2_fill_1 FILLER_62_255 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_fill_2 FILLER_62_278 ();
 sg13g2_fill_2 FILLER_62_288 ();
 sg13g2_fill_1 FILLER_62_290 ();
 sg13g2_fill_1 FILLER_62_295 ();
 sg13g2_fill_2 FILLER_62_467 ();
 sg13g2_fill_1 FILLER_62_469 ();
 sg13g2_fill_2 FILLER_62_483 ();
 sg13g2_fill_1 FILLER_62_518 ();
 sg13g2_decap_8 FILLER_62_529 ();
 sg13g2_decap_8 FILLER_62_536 ();
 sg13g2_decap_8 FILLER_62_543 ();
 sg13g2_decap_4 FILLER_62_550 ();
 sg13g2_fill_2 FILLER_62_554 ();
 sg13g2_decap_4 FILLER_62_559 ();
 sg13g2_fill_1 FILLER_62_563 ();
 sg13g2_fill_2 FILLER_62_605 ();
 sg13g2_fill_1 FILLER_62_638 ();
 sg13g2_fill_2 FILLER_62_663 ();
 sg13g2_fill_2 FILLER_62_681 ();
 sg13g2_fill_2 FILLER_62_696 ();
 sg13g2_fill_1 FILLER_62_698 ();
 sg13g2_decap_8 FILLER_62_723 ();
 sg13g2_decap_8 FILLER_62_730 ();
 sg13g2_decap_8 FILLER_62_737 ();
 sg13g2_decap_8 FILLER_62_744 ();
 sg13g2_decap_8 FILLER_62_751 ();
 sg13g2_decap_8 FILLER_62_758 ();
 sg13g2_decap_8 FILLER_62_765 ();
 sg13g2_decap_8 FILLER_62_772 ();
 sg13g2_decap_8 FILLER_62_779 ();
 sg13g2_decap_8 FILLER_62_786 ();
 sg13g2_decap_8 FILLER_62_793 ();
 sg13g2_decap_8 FILLER_62_800 ();
 sg13g2_decap_8 FILLER_62_807 ();
 sg13g2_decap_8 FILLER_62_814 ();
 sg13g2_decap_8 FILLER_62_821 ();
 sg13g2_decap_8 FILLER_62_828 ();
 sg13g2_decap_8 FILLER_62_835 ();
 sg13g2_decap_8 FILLER_62_842 ();
 sg13g2_decap_8 FILLER_62_849 ();
 sg13g2_decap_4 FILLER_62_856 ();
 sg13g2_fill_2 FILLER_62_860 ();
 sg13g2_fill_2 FILLER_63_83 ();
 sg13g2_fill_2 FILLER_63_210 ();
 sg13g2_fill_2 FILLER_63_221 ();
 sg13g2_decap_4 FILLER_63_269 ();
 sg13g2_fill_2 FILLER_63_273 ();
 sg13g2_fill_2 FILLER_63_280 ();
 sg13g2_fill_1 FILLER_63_282 ();
 sg13g2_decap_4 FILLER_63_288 ();
 sg13g2_fill_2 FILLER_63_292 ();
 sg13g2_fill_1 FILLER_63_322 ();
 sg13g2_fill_2 FILLER_63_332 ();
 sg13g2_fill_2 FILLER_63_340 ();
 sg13g2_fill_1 FILLER_63_342 ();
 sg13g2_fill_2 FILLER_63_370 ();
 sg13g2_fill_2 FILLER_63_386 ();
 sg13g2_fill_2 FILLER_63_433 ();
 sg13g2_decap_8 FILLER_63_509 ();
 sg13g2_fill_2 FILLER_63_516 ();
 sg13g2_fill_2 FILLER_63_557 ();
 sg13g2_decap_4 FILLER_63_567 ();
 sg13g2_fill_2 FILLER_63_639 ();
 sg13g2_fill_2 FILLER_63_659 ();
 sg13g2_fill_2 FILLER_63_676 ();
 sg13g2_fill_2 FILLER_63_688 ();
 sg13g2_decap_8 FILLER_63_726 ();
 sg13g2_decap_8 FILLER_63_733 ();
 sg13g2_decap_8 FILLER_63_740 ();
 sg13g2_decap_8 FILLER_63_747 ();
 sg13g2_decap_8 FILLER_63_754 ();
 sg13g2_decap_8 FILLER_63_761 ();
 sg13g2_decap_8 FILLER_63_768 ();
 sg13g2_decap_8 FILLER_63_775 ();
 sg13g2_decap_8 FILLER_63_782 ();
 sg13g2_decap_8 FILLER_63_789 ();
 sg13g2_decap_8 FILLER_63_796 ();
 sg13g2_decap_8 FILLER_63_803 ();
 sg13g2_decap_8 FILLER_63_810 ();
 sg13g2_decap_8 FILLER_63_817 ();
 sg13g2_decap_8 FILLER_63_824 ();
 sg13g2_decap_8 FILLER_63_831 ();
 sg13g2_decap_8 FILLER_63_838 ();
 sg13g2_decap_8 FILLER_63_845 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_fill_2 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_861 ();
 sg13g2_fill_2 FILLER_64_37 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_fill_2 FILLER_64_167 ();
 sg13g2_fill_2 FILLER_64_209 ();
 sg13g2_decap_4 FILLER_64_289 ();
 sg13g2_fill_2 FILLER_64_293 ();
 sg13g2_fill_2 FILLER_64_312 ();
 sg13g2_fill_2 FILLER_64_477 ();
 sg13g2_fill_2 FILLER_64_498 ();
 sg13g2_fill_1 FILLER_64_500 ();
 sg13g2_fill_2 FILLER_64_504 ();
 sg13g2_decap_8 FILLER_64_510 ();
 sg13g2_fill_2 FILLER_64_588 ();
 sg13g2_fill_2 FILLER_64_620 ();
 sg13g2_fill_1 FILLER_64_657 ();
 sg13g2_decap_8 FILLER_64_716 ();
 sg13g2_decap_8 FILLER_64_723 ();
 sg13g2_decap_8 FILLER_64_730 ();
 sg13g2_decap_8 FILLER_64_737 ();
 sg13g2_decap_8 FILLER_64_744 ();
 sg13g2_decap_8 FILLER_64_751 ();
 sg13g2_decap_8 FILLER_64_758 ();
 sg13g2_decap_8 FILLER_64_765 ();
 sg13g2_decap_8 FILLER_64_772 ();
 sg13g2_decap_8 FILLER_64_779 ();
 sg13g2_decap_8 FILLER_64_786 ();
 sg13g2_decap_8 FILLER_64_793 ();
 sg13g2_decap_8 FILLER_64_800 ();
 sg13g2_decap_8 FILLER_64_807 ();
 sg13g2_decap_8 FILLER_64_814 ();
 sg13g2_decap_8 FILLER_64_821 ();
 sg13g2_decap_8 FILLER_64_828 ();
 sg13g2_decap_8 FILLER_64_835 ();
 sg13g2_decap_8 FILLER_64_842 ();
 sg13g2_decap_8 FILLER_64_849 ();
 sg13g2_decap_4 FILLER_64_856 ();
 sg13g2_fill_2 FILLER_64_860 ();
 sg13g2_fill_2 FILLER_65_33 ();
 sg13g2_fill_2 FILLER_65_81 ();
 sg13g2_fill_2 FILLER_65_176 ();
 sg13g2_fill_1 FILLER_65_230 ();
 sg13g2_fill_1 FILLER_65_244 ();
 sg13g2_fill_1 FILLER_65_285 ();
 sg13g2_fill_1 FILLER_65_290 ();
 sg13g2_fill_2 FILLER_65_319 ();
 sg13g2_fill_1 FILLER_65_321 ();
 sg13g2_fill_2 FILLER_65_327 ();
 sg13g2_fill_1 FILLER_65_366 ();
 sg13g2_fill_2 FILLER_65_384 ();
 sg13g2_fill_1 FILLER_65_386 ();
 sg13g2_fill_2 FILLER_65_396 ();
 sg13g2_fill_1 FILLER_65_398 ();
 sg13g2_fill_1 FILLER_65_442 ();
 sg13g2_fill_2 FILLER_65_456 ();
 sg13g2_fill_1 FILLER_65_471 ();
 sg13g2_decap_8 FILLER_65_495 ();
 sg13g2_decap_8 FILLER_65_502 ();
 sg13g2_fill_1 FILLER_65_512 ();
 sg13g2_fill_2 FILLER_65_541 ();
 sg13g2_fill_1 FILLER_65_543 ();
 sg13g2_fill_2 FILLER_65_552 ();
 sg13g2_fill_1 FILLER_65_624 ();
 sg13g2_fill_2 FILLER_65_670 ();
 sg13g2_fill_2 FILLER_65_699 ();
 sg13g2_decap_8 FILLER_65_714 ();
 sg13g2_decap_8 FILLER_65_721 ();
 sg13g2_decap_8 FILLER_65_728 ();
 sg13g2_decap_8 FILLER_65_735 ();
 sg13g2_decap_8 FILLER_65_742 ();
 sg13g2_decap_8 FILLER_65_749 ();
 sg13g2_decap_8 FILLER_65_756 ();
 sg13g2_decap_8 FILLER_65_763 ();
 sg13g2_decap_8 FILLER_65_770 ();
 sg13g2_decap_8 FILLER_65_777 ();
 sg13g2_decap_8 FILLER_65_784 ();
 sg13g2_decap_8 FILLER_65_791 ();
 sg13g2_decap_8 FILLER_65_798 ();
 sg13g2_decap_8 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_decap_8 FILLER_65_819 ();
 sg13g2_decap_8 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_65_847 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_fill_1 FILLER_65_861 ();
 sg13g2_fill_1 FILLER_66_0 ();
 sg13g2_fill_2 FILLER_66_86 ();
 sg13g2_fill_2 FILLER_66_172 ();
 sg13g2_fill_1 FILLER_66_174 ();
 sg13g2_fill_2 FILLER_66_197 ();
 sg13g2_fill_2 FILLER_66_236 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_fill_2 FILLER_66_288 ();
 sg13g2_fill_1 FILLER_66_331 ();
 sg13g2_fill_2 FILLER_66_338 ();
 sg13g2_fill_1 FILLER_66_340 ();
 sg13g2_decap_8 FILLER_66_346 ();
 sg13g2_fill_2 FILLER_66_353 ();
 sg13g2_fill_1 FILLER_66_355 ();
 sg13g2_fill_2 FILLER_66_376 ();
 sg13g2_fill_1 FILLER_66_378 ();
 sg13g2_fill_2 FILLER_66_399 ();
 sg13g2_fill_1 FILLER_66_439 ();
 sg13g2_fill_1 FILLER_66_534 ();
 sg13g2_fill_2 FILLER_66_540 ();
 sg13g2_fill_2 FILLER_66_640 ();
 sg13g2_fill_1 FILLER_66_642 ();
 sg13g2_fill_1 FILLER_66_679 ();
 sg13g2_decap_8 FILLER_66_712 ();
 sg13g2_decap_8 FILLER_66_719 ();
 sg13g2_decap_8 FILLER_66_726 ();
 sg13g2_decap_8 FILLER_66_733 ();
 sg13g2_decap_8 FILLER_66_740 ();
 sg13g2_decap_8 FILLER_66_747 ();
 sg13g2_decap_8 FILLER_66_754 ();
 sg13g2_decap_8 FILLER_66_761 ();
 sg13g2_decap_8 FILLER_66_768 ();
 sg13g2_decap_8 FILLER_66_775 ();
 sg13g2_decap_8 FILLER_66_782 ();
 sg13g2_decap_8 FILLER_66_789 ();
 sg13g2_decap_8 FILLER_66_796 ();
 sg13g2_decap_8 FILLER_66_803 ();
 sg13g2_decap_8 FILLER_66_810 ();
 sg13g2_decap_8 FILLER_66_817 ();
 sg13g2_decap_8 FILLER_66_824 ();
 sg13g2_decap_8 FILLER_66_831 ();
 sg13g2_decap_8 FILLER_66_838 ();
 sg13g2_decap_8 FILLER_66_845 ();
 sg13g2_decap_8 FILLER_66_852 ();
 sg13g2_fill_2 FILLER_66_859 ();
 sg13g2_fill_1 FILLER_66_861 ();
 sg13g2_fill_1 FILLER_67_0 ();
 sg13g2_fill_1 FILLER_67_179 ();
 sg13g2_fill_2 FILLER_67_207 ();
 sg13g2_decap_4 FILLER_67_263 ();
 sg13g2_fill_2 FILLER_67_267 ();
 sg13g2_fill_2 FILLER_67_303 ();
 sg13g2_fill_1 FILLER_67_314 ();
 sg13g2_fill_2 FILLER_67_340 ();
 sg13g2_fill_1 FILLER_67_342 ();
 sg13g2_decap_4 FILLER_67_352 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_decap_4 FILLER_67_363 ();
 sg13g2_fill_2 FILLER_67_391 ();
 sg13g2_decap_4 FILLER_67_492 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_fill_2 FILLER_67_511 ();
 sg13g2_fill_1 FILLER_67_513 ();
 sg13g2_fill_2 FILLER_67_529 ();
 sg13g2_fill_1 FILLER_67_599 ();
 sg13g2_fill_2 FILLER_67_666 ();
 sg13g2_decap_8 FILLER_67_701 ();
 sg13g2_decap_8 FILLER_67_708 ();
 sg13g2_decap_8 FILLER_67_715 ();
 sg13g2_decap_8 FILLER_67_722 ();
 sg13g2_decap_8 FILLER_67_729 ();
 sg13g2_decap_8 FILLER_67_736 ();
 sg13g2_decap_8 FILLER_67_743 ();
 sg13g2_decap_8 FILLER_67_750 ();
 sg13g2_decap_8 FILLER_67_757 ();
 sg13g2_decap_8 FILLER_67_764 ();
 sg13g2_decap_8 FILLER_67_771 ();
 sg13g2_decap_8 FILLER_67_778 ();
 sg13g2_decap_8 FILLER_67_785 ();
 sg13g2_decap_8 FILLER_67_792 ();
 sg13g2_decap_8 FILLER_67_799 ();
 sg13g2_decap_8 FILLER_67_806 ();
 sg13g2_decap_8 FILLER_67_813 ();
 sg13g2_decap_8 FILLER_67_820 ();
 sg13g2_decap_8 FILLER_67_827 ();
 sg13g2_decap_8 FILLER_67_834 ();
 sg13g2_decap_8 FILLER_67_841 ();
 sg13g2_decap_8 FILLER_67_848 ();
 sg13g2_decap_8 FILLER_67_855 ();
 sg13g2_fill_1 FILLER_68_33 ();
 sg13g2_fill_2 FILLER_68_128 ();
 sg13g2_fill_1 FILLER_68_154 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_179 ();
 sg13g2_fill_2 FILLER_68_220 ();
 sg13g2_fill_1 FILLER_68_231 ();
 sg13g2_fill_2 FILLER_68_265 ();
 sg13g2_fill_2 FILLER_68_282 ();
 sg13g2_fill_2 FILLER_68_322 ();
 sg13g2_fill_1 FILLER_68_324 ();
 sg13g2_fill_2 FILLER_68_358 ();
 sg13g2_fill_1 FILLER_68_360 ();
 sg13g2_fill_1 FILLER_68_366 ();
 sg13g2_fill_1 FILLER_68_372 ();
 sg13g2_fill_2 FILLER_68_429 ();
 sg13g2_fill_2 FILLER_68_466 ();
 sg13g2_fill_1 FILLER_68_468 ();
 sg13g2_fill_2 FILLER_68_505 ();
 sg13g2_decap_8 FILLER_68_722 ();
 sg13g2_decap_8 FILLER_68_729 ();
 sg13g2_decap_8 FILLER_68_736 ();
 sg13g2_decap_8 FILLER_68_743 ();
 sg13g2_decap_8 FILLER_68_750 ();
 sg13g2_decap_8 FILLER_68_757 ();
 sg13g2_decap_8 FILLER_68_764 ();
 sg13g2_decap_8 FILLER_68_771 ();
 sg13g2_decap_8 FILLER_68_778 ();
 sg13g2_decap_8 FILLER_68_785 ();
 sg13g2_decap_8 FILLER_68_792 ();
 sg13g2_decap_8 FILLER_68_799 ();
 sg13g2_decap_8 FILLER_68_806 ();
 sg13g2_decap_8 FILLER_68_813 ();
 sg13g2_decap_8 FILLER_68_820 ();
 sg13g2_decap_8 FILLER_68_827 ();
 sg13g2_decap_8 FILLER_68_834 ();
 sg13g2_decap_8 FILLER_68_841 ();
 sg13g2_decap_8 FILLER_68_848 ();
 sg13g2_decap_8 FILLER_68_855 ();
 sg13g2_fill_2 FILLER_69_56 ();
 sg13g2_fill_2 FILLER_69_125 ();
 sg13g2_fill_1 FILLER_69_127 ();
 sg13g2_fill_2 FILLER_69_146 ();
 sg13g2_fill_2 FILLER_69_157 ();
 sg13g2_fill_1 FILLER_69_159 ();
 sg13g2_fill_1 FILLER_69_230 ();
 sg13g2_fill_2 FILLER_69_288 ();
 sg13g2_fill_1 FILLER_69_290 ();
 sg13g2_fill_1 FILLER_69_300 ();
 sg13g2_fill_2 FILLER_69_411 ();
 sg13g2_fill_1 FILLER_69_422 ();
 sg13g2_fill_2 FILLER_69_468 ();
 sg13g2_fill_2 FILLER_69_500 ();
 sg13g2_fill_1 FILLER_69_511 ();
 sg13g2_fill_2 FILLER_69_604 ();
 sg13g2_fill_1 FILLER_69_633 ();
 sg13g2_decap_4 FILLER_69_674 ();
 sg13g2_fill_2 FILLER_69_678 ();
 sg13g2_fill_1 FILLER_69_684 ();
 sg13g2_fill_1 FILLER_69_692 ();
 sg13g2_fill_1 FILLER_69_705 ();
 sg13g2_decap_8 FILLER_69_715 ();
 sg13g2_decap_8 FILLER_69_722 ();
 sg13g2_decap_8 FILLER_69_729 ();
 sg13g2_decap_8 FILLER_69_736 ();
 sg13g2_decap_8 FILLER_69_743 ();
 sg13g2_decap_8 FILLER_69_750 ();
 sg13g2_decap_8 FILLER_69_757 ();
 sg13g2_decap_8 FILLER_69_764 ();
 sg13g2_decap_8 FILLER_69_771 ();
 sg13g2_decap_8 FILLER_69_778 ();
 sg13g2_decap_8 FILLER_69_785 ();
 sg13g2_decap_8 FILLER_69_792 ();
 sg13g2_decap_8 FILLER_69_799 ();
 sg13g2_decap_8 FILLER_69_806 ();
 sg13g2_decap_8 FILLER_69_813 ();
 sg13g2_decap_8 FILLER_69_820 ();
 sg13g2_decap_8 FILLER_69_827 ();
 sg13g2_decap_8 FILLER_69_834 ();
 sg13g2_decap_8 FILLER_69_841 ();
 sg13g2_decap_8 FILLER_69_848 ();
 sg13g2_decap_8 FILLER_69_855 ();
 sg13g2_fill_1 FILLER_70_33 ();
 sg13g2_fill_2 FILLER_70_101 ();
 sg13g2_fill_2 FILLER_70_136 ();
 sg13g2_fill_1 FILLER_70_138 ();
 sg13g2_fill_1 FILLER_70_218 ();
 sg13g2_fill_1 FILLER_70_250 ();
 sg13g2_fill_1 FILLER_70_271 ();
 sg13g2_fill_2 FILLER_70_279 ();
 sg13g2_fill_2 FILLER_70_286 ();
 sg13g2_decap_8 FILLER_70_345 ();
 sg13g2_decap_4 FILLER_70_352 ();
 sg13g2_fill_1 FILLER_70_378 ();
 sg13g2_fill_2 FILLER_70_392 ();
 sg13g2_fill_1 FILLER_70_403 ();
 sg13g2_fill_2 FILLER_70_431 ();
 sg13g2_fill_1 FILLER_70_495 ();
 sg13g2_fill_1 FILLER_70_610 ();
 sg13g2_fill_2 FILLER_70_625 ();
 sg13g2_decap_8 FILLER_70_725 ();
 sg13g2_decap_8 FILLER_70_732 ();
 sg13g2_decap_8 FILLER_70_739 ();
 sg13g2_decap_8 FILLER_70_746 ();
 sg13g2_decap_8 FILLER_70_753 ();
 sg13g2_decap_8 FILLER_70_760 ();
 sg13g2_decap_8 FILLER_70_767 ();
 sg13g2_decap_8 FILLER_70_774 ();
 sg13g2_decap_8 FILLER_70_781 ();
 sg13g2_decap_8 FILLER_70_788 ();
 sg13g2_decap_8 FILLER_70_795 ();
 sg13g2_decap_8 FILLER_70_802 ();
 sg13g2_decap_8 FILLER_70_809 ();
 sg13g2_decap_8 FILLER_70_816 ();
 sg13g2_decap_8 FILLER_70_823 ();
 sg13g2_decap_8 FILLER_70_830 ();
 sg13g2_decap_8 FILLER_70_837 ();
 sg13g2_decap_8 FILLER_70_844 ();
 sg13g2_decap_8 FILLER_70_851 ();
 sg13g2_decap_4 FILLER_70_858 ();
 sg13g2_fill_2 FILLER_71_34 ();
 sg13g2_fill_1 FILLER_71_45 ();
 sg13g2_fill_2 FILLER_71_63 ();
 sg13g2_fill_2 FILLER_71_161 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_fill_2 FILLER_71_387 ();
 sg13g2_fill_2 FILLER_71_419 ();
 sg13g2_fill_1 FILLER_71_421 ();
 sg13g2_fill_1 FILLER_71_460 ();
 sg13g2_fill_1 FILLER_71_527 ();
 sg13g2_fill_1 FILLER_71_542 ();
 sg13g2_fill_1 FILLER_71_594 ();
 sg13g2_fill_2 FILLER_71_637 ();
 sg13g2_fill_1 FILLER_71_661 ();
 sg13g2_fill_2 FILLER_71_666 ();
 sg13g2_fill_2 FILLER_71_686 ();
 sg13g2_fill_1 FILLER_71_688 ();
 sg13g2_decap_8 FILLER_71_735 ();
 sg13g2_decap_8 FILLER_71_742 ();
 sg13g2_decap_8 FILLER_71_749 ();
 sg13g2_decap_8 FILLER_71_756 ();
 sg13g2_decap_8 FILLER_71_763 ();
 sg13g2_decap_8 FILLER_71_770 ();
 sg13g2_decap_8 FILLER_71_777 ();
 sg13g2_decap_8 FILLER_71_784 ();
 sg13g2_decap_8 FILLER_71_791 ();
 sg13g2_decap_8 FILLER_71_798 ();
 sg13g2_decap_8 FILLER_71_805 ();
 sg13g2_decap_8 FILLER_71_812 ();
 sg13g2_decap_8 FILLER_71_819 ();
 sg13g2_decap_8 FILLER_71_826 ();
 sg13g2_decap_8 FILLER_71_833 ();
 sg13g2_decap_8 FILLER_71_840 ();
 sg13g2_decap_8 FILLER_71_847 ();
 sg13g2_decap_8 FILLER_71_854 ();
 sg13g2_fill_1 FILLER_71_861 ();
 sg13g2_fill_1 FILLER_72_129 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_fill_1 FILLER_72_264 ();
 sg13g2_fill_1 FILLER_72_297 ();
 sg13g2_fill_2 FILLER_72_307 ();
 sg13g2_fill_2 FILLER_72_317 ();
 sg13g2_fill_1 FILLER_72_319 ();
 sg13g2_fill_2 FILLER_72_332 ();
 sg13g2_fill_2 FILLER_72_343 ();
 sg13g2_fill_2 FILLER_72_363 ();
 sg13g2_fill_1 FILLER_72_365 ();
 sg13g2_fill_2 FILLER_72_425 ();
 sg13g2_fill_1 FILLER_72_427 ();
 sg13g2_fill_2 FILLER_72_437 ();
 sg13g2_fill_2 FILLER_72_473 ();
 sg13g2_fill_1 FILLER_72_609 ();
 sg13g2_fill_2 FILLER_72_660 ();
 sg13g2_fill_2 FILLER_72_682 ();
 sg13g2_fill_1 FILLER_72_684 ();
 sg13g2_decap_8 FILLER_72_735 ();
 sg13g2_decap_8 FILLER_72_742 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_decap_8 FILLER_72_756 ();
 sg13g2_decap_8 FILLER_72_763 ();
 sg13g2_decap_8 FILLER_72_770 ();
 sg13g2_decap_8 FILLER_72_777 ();
 sg13g2_decap_8 FILLER_72_784 ();
 sg13g2_decap_8 FILLER_72_791 ();
 sg13g2_decap_8 FILLER_72_798 ();
 sg13g2_decap_8 FILLER_72_805 ();
 sg13g2_decap_8 FILLER_72_812 ();
 sg13g2_decap_8 FILLER_72_819 ();
 sg13g2_decap_8 FILLER_72_826 ();
 sg13g2_decap_8 FILLER_72_833 ();
 sg13g2_decap_8 FILLER_72_840 ();
 sg13g2_decap_8 FILLER_72_847 ();
 sg13g2_decap_8 FILLER_72_854 ();
 sg13g2_fill_1 FILLER_72_861 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_98 ();
 sg13g2_fill_1 FILLER_73_113 ();
 sg13g2_fill_1 FILLER_73_142 ();
 sg13g2_fill_1 FILLER_73_266 ();
 sg13g2_fill_2 FILLER_73_289 ();
 sg13g2_fill_2 FILLER_73_308 ();
 sg13g2_fill_2 FILLER_73_323 ();
 sg13g2_fill_1 FILLER_73_325 ();
 sg13g2_fill_2 FILLER_73_352 ();
 sg13g2_fill_1 FILLER_73_354 ();
 sg13g2_fill_1 FILLER_73_364 ();
 sg13g2_fill_1 FILLER_73_375 ();
 sg13g2_fill_2 FILLER_73_398 ();
 sg13g2_fill_2 FILLER_73_406 ();
 sg13g2_fill_1 FILLER_73_408 ();
 sg13g2_decap_8 FILLER_73_422 ();
 sg13g2_fill_2 FILLER_73_429 ();
 sg13g2_fill_2 FILLER_73_446 ();
 sg13g2_fill_2 FILLER_73_457 ();
 sg13g2_fill_1 FILLER_73_459 ();
 sg13g2_fill_2 FILLER_73_474 ();
 sg13g2_fill_1 FILLER_73_476 ();
 sg13g2_fill_2 FILLER_73_510 ();
 sg13g2_fill_2 FILLER_73_542 ();
 sg13g2_fill_2 FILLER_73_639 ();
 sg13g2_decap_8 FILLER_73_731 ();
 sg13g2_decap_8 FILLER_73_738 ();
 sg13g2_decap_8 FILLER_73_745 ();
 sg13g2_decap_8 FILLER_73_752 ();
 sg13g2_decap_8 FILLER_73_759 ();
 sg13g2_decap_8 FILLER_73_766 ();
 sg13g2_decap_8 FILLER_73_773 ();
 sg13g2_decap_8 FILLER_73_780 ();
 sg13g2_decap_8 FILLER_73_787 ();
 sg13g2_decap_8 FILLER_73_794 ();
 sg13g2_decap_8 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_808 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_decap_8 FILLER_73_822 ();
 sg13g2_decap_8 FILLER_73_829 ();
 sg13g2_decap_8 FILLER_73_836 ();
 sg13g2_decap_8 FILLER_73_843 ();
 sg13g2_decap_8 FILLER_73_850 ();
 sg13g2_decap_4 FILLER_73_857 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_fill_1 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_29 ();
 sg13g2_fill_1 FILLER_74_49 ();
 sg13g2_fill_2 FILLER_74_125 ();
 sg13g2_fill_2 FILLER_74_154 ();
 sg13g2_fill_1 FILLER_74_156 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_2 FILLER_74_225 ();
 sg13g2_fill_2 FILLER_74_232 ();
 sg13g2_fill_1 FILLER_74_243 ();
 sg13g2_fill_1 FILLER_74_258 ();
 sg13g2_fill_1 FILLER_74_264 ();
 sg13g2_fill_2 FILLER_74_278 ();
 sg13g2_fill_1 FILLER_74_305 ();
 sg13g2_fill_2 FILLER_74_337 ();
 sg13g2_fill_1 FILLER_74_339 ();
 sg13g2_fill_2 FILLER_74_368 ();
 sg13g2_fill_2 FILLER_74_375 ();
 sg13g2_decap_4 FILLER_74_437 ();
 sg13g2_fill_1 FILLER_74_445 ();
 sg13g2_fill_2 FILLER_74_449 ();
 sg13g2_decap_4 FILLER_74_504 ();
 sg13g2_fill_2 FILLER_74_508 ();
 sg13g2_fill_2 FILLER_74_518 ();
 sg13g2_fill_1 FILLER_74_520 ();
 sg13g2_fill_1 FILLER_74_569 ();
 sg13g2_fill_2 FILLER_74_624 ();
 sg13g2_decap_8 FILLER_74_629 ();
 sg13g2_fill_2 FILLER_74_636 ();
 sg13g2_fill_1 FILLER_74_638 ();
 sg13g2_decap_8 FILLER_74_643 ();
 sg13g2_decap_4 FILLER_74_650 ();
 sg13g2_fill_1 FILLER_74_654 ();
 sg13g2_decap_8 FILLER_74_659 ();
 sg13g2_decap_8 FILLER_74_666 ();
 sg13g2_decap_4 FILLER_74_673 ();
 sg13g2_fill_1 FILLER_74_677 ();
 sg13g2_decap_8 FILLER_74_682 ();
 sg13g2_fill_2 FILLER_74_695 ();
 sg13g2_fill_1 FILLER_74_711 ();
 sg13g2_decap_8 FILLER_74_721 ();
 sg13g2_decap_8 FILLER_74_728 ();
 sg13g2_decap_8 FILLER_74_735 ();
 sg13g2_decap_8 FILLER_74_742 ();
 sg13g2_decap_8 FILLER_74_749 ();
 sg13g2_decap_8 FILLER_74_756 ();
 sg13g2_decap_8 FILLER_74_763 ();
 sg13g2_decap_8 FILLER_74_770 ();
 sg13g2_decap_8 FILLER_74_777 ();
 sg13g2_decap_8 FILLER_74_784 ();
 sg13g2_decap_8 FILLER_74_791 ();
 sg13g2_decap_8 FILLER_74_798 ();
 sg13g2_decap_8 FILLER_74_805 ();
 sg13g2_decap_8 FILLER_74_812 ();
 sg13g2_decap_8 FILLER_74_819 ();
 sg13g2_decap_8 FILLER_74_826 ();
 sg13g2_decap_8 FILLER_74_833 ();
 sg13g2_decap_8 FILLER_74_840 ();
 sg13g2_decap_8 FILLER_74_847 ();
 sg13g2_decap_8 FILLER_74_854 ();
 sg13g2_fill_1 FILLER_74_861 ();
 sg13g2_fill_2 FILLER_75_83 ();
 sg13g2_fill_1 FILLER_75_85 ();
 sg13g2_fill_1 FILLER_75_100 ();
 sg13g2_fill_2 FILLER_75_141 ();
 sg13g2_fill_1 FILLER_75_143 ();
 sg13g2_fill_2 FILLER_75_180 ();
 sg13g2_fill_2 FILLER_75_302 ();
 sg13g2_fill_1 FILLER_75_304 ();
 sg13g2_fill_2 FILLER_75_309 ();
 sg13g2_fill_1 FILLER_75_311 ();
 sg13g2_fill_2 FILLER_75_329 ();
 sg13g2_fill_1 FILLER_75_331 ();
 sg13g2_fill_1 FILLER_75_381 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_fill_2 FILLER_75_400 ();
 sg13g2_decap_8 FILLER_75_421 ();
 sg13g2_decap_8 FILLER_75_428 ();
 sg13g2_fill_1 FILLER_75_435 ();
 sg13g2_fill_2 FILLER_75_440 ();
 sg13g2_fill_1 FILLER_75_442 ();
 sg13g2_fill_2 FILLER_75_456 ();
 sg13g2_fill_2 FILLER_75_497 ();
 sg13g2_fill_2 FILLER_75_517 ();
 sg13g2_fill_1 FILLER_75_524 ();
 sg13g2_decap_4 FILLER_75_547 ();
 sg13g2_decap_8 FILLER_75_559 ();
 sg13g2_decap_8 FILLER_75_566 ();
 sg13g2_fill_2 FILLER_75_573 ();
 sg13g2_fill_1 FILLER_75_575 ();
 sg13g2_fill_2 FILLER_75_591 ();
 sg13g2_decap_8 FILLER_75_614 ();
 sg13g2_decap_8 FILLER_75_621 ();
 sg13g2_decap_8 FILLER_75_628 ();
 sg13g2_decap_8 FILLER_75_635 ();
 sg13g2_decap_8 FILLER_75_642 ();
 sg13g2_decap_8 FILLER_75_649 ();
 sg13g2_decap_8 FILLER_75_656 ();
 sg13g2_decap_8 FILLER_75_663 ();
 sg13g2_decap_8 FILLER_75_670 ();
 sg13g2_decap_8 FILLER_75_677 ();
 sg13g2_decap_8 FILLER_75_684 ();
 sg13g2_decap_8 FILLER_75_691 ();
 sg13g2_decap_8 FILLER_75_698 ();
 sg13g2_decap_8 FILLER_75_705 ();
 sg13g2_decap_8 FILLER_75_712 ();
 sg13g2_decap_8 FILLER_75_719 ();
 sg13g2_decap_8 FILLER_75_726 ();
 sg13g2_decap_8 FILLER_75_733 ();
 sg13g2_decap_8 FILLER_75_740 ();
 sg13g2_decap_8 FILLER_75_747 ();
 sg13g2_decap_8 FILLER_75_754 ();
 sg13g2_decap_8 FILLER_75_761 ();
 sg13g2_decap_8 FILLER_75_768 ();
 sg13g2_decap_8 FILLER_75_775 ();
 sg13g2_decap_8 FILLER_75_782 ();
 sg13g2_decap_8 FILLER_75_789 ();
 sg13g2_decap_8 FILLER_75_796 ();
 sg13g2_decap_8 FILLER_75_803 ();
 sg13g2_decap_8 FILLER_75_810 ();
 sg13g2_decap_8 FILLER_75_817 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_8 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_859 ();
 sg13g2_fill_1 FILLER_75_861 ();
 sg13g2_fill_2 FILLER_76_27 ();
 sg13g2_fill_1 FILLER_76_55 ();
 sg13g2_fill_1 FILLER_76_95 ();
 sg13g2_fill_1 FILLER_76_200 ();
 sg13g2_fill_1 FILLER_76_292 ();
 sg13g2_fill_2 FILLER_76_298 ();
 sg13g2_fill_2 FILLER_76_335 ();
 sg13g2_decap_4 FILLER_76_388 ();
 sg13g2_fill_2 FILLER_76_392 ();
 sg13g2_fill_1 FILLER_76_400 ();
 sg13g2_fill_2 FILLER_76_414 ();
 sg13g2_decap_8 FILLER_76_420 ();
 sg13g2_decap_4 FILLER_76_427 ();
 sg13g2_fill_1 FILLER_76_472 ();
 sg13g2_fill_1 FILLER_76_494 ();
 sg13g2_decap_8 FILLER_76_536 ();
 sg13g2_decap_8 FILLER_76_543 ();
 sg13g2_decap_8 FILLER_76_550 ();
 sg13g2_decap_8 FILLER_76_557 ();
 sg13g2_decap_8 FILLER_76_564 ();
 sg13g2_decap_8 FILLER_76_571 ();
 sg13g2_decap_8 FILLER_76_578 ();
 sg13g2_decap_8 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_592 ();
 sg13g2_decap_8 FILLER_76_599 ();
 sg13g2_decap_8 FILLER_76_606 ();
 sg13g2_decap_8 FILLER_76_613 ();
 sg13g2_decap_8 FILLER_76_620 ();
 sg13g2_decap_8 FILLER_76_627 ();
 sg13g2_decap_8 FILLER_76_634 ();
 sg13g2_decap_8 FILLER_76_641 ();
 sg13g2_decap_8 FILLER_76_648 ();
 sg13g2_decap_8 FILLER_76_655 ();
 sg13g2_decap_8 FILLER_76_662 ();
 sg13g2_decap_8 FILLER_76_669 ();
 sg13g2_decap_8 FILLER_76_676 ();
 sg13g2_decap_8 FILLER_76_683 ();
 sg13g2_decap_8 FILLER_76_690 ();
 sg13g2_decap_8 FILLER_76_697 ();
 sg13g2_decap_8 FILLER_76_704 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_8 FILLER_76_718 ();
 sg13g2_decap_8 FILLER_76_725 ();
 sg13g2_decap_8 FILLER_76_732 ();
 sg13g2_decap_8 FILLER_76_739 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_767 ();
 sg13g2_decap_8 FILLER_76_774 ();
 sg13g2_decap_8 FILLER_76_781 ();
 sg13g2_decap_8 FILLER_76_788 ();
 sg13g2_decap_8 FILLER_76_795 ();
 sg13g2_decap_8 FILLER_76_802 ();
 sg13g2_decap_8 FILLER_76_809 ();
 sg13g2_decap_8 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_decap_8 FILLER_76_837 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_decap_8 FILLER_76_851 ();
 sg13g2_decap_4 FILLER_76_858 ();
 sg13g2_fill_1 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_41 ();
 sg13g2_fill_1 FILLER_77_55 ();
 sg13g2_fill_2 FILLER_77_128 ();
 sg13g2_fill_2 FILLER_77_173 ();
 sg13g2_fill_1 FILLER_77_237 ();
 sg13g2_fill_2 FILLER_77_291 ();
 sg13g2_fill_1 FILLER_77_293 ();
 sg13g2_fill_2 FILLER_77_299 ();
 sg13g2_fill_1 FILLER_77_301 ();
 sg13g2_fill_1 FILLER_77_317 ();
 sg13g2_fill_2 FILLER_77_373 ();
 sg13g2_fill_1 FILLER_77_375 ();
 sg13g2_fill_1 FILLER_77_393 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_fill_1 FILLER_77_409 ();
 sg13g2_fill_1 FILLER_77_465 ();
 sg13g2_fill_2 FILLER_77_507 ();
 sg13g2_decap_8 FILLER_77_544 ();
 sg13g2_decap_8 FILLER_77_551 ();
 sg13g2_decap_8 FILLER_77_558 ();
 sg13g2_decap_8 FILLER_77_565 ();
 sg13g2_decap_8 FILLER_77_572 ();
 sg13g2_decap_8 FILLER_77_579 ();
 sg13g2_decap_8 FILLER_77_586 ();
 sg13g2_decap_8 FILLER_77_593 ();
 sg13g2_decap_8 FILLER_77_600 ();
 sg13g2_decap_8 FILLER_77_607 ();
 sg13g2_decap_8 FILLER_77_614 ();
 sg13g2_decap_8 FILLER_77_621 ();
 sg13g2_decap_8 FILLER_77_628 ();
 sg13g2_decap_8 FILLER_77_635 ();
 sg13g2_decap_8 FILLER_77_642 ();
 sg13g2_decap_8 FILLER_77_649 ();
 sg13g2_decap_8 FILLER_77_656 ();
 sg13g2_decap_8 FILLER_77_663 ();
 sg13g2_decap_8 FILLER_77_670 ();
 sg13g2_decap_8 FILLER_77_677 ();
 sg13g2_decap_8 FILLER_77_684 ();
 sg13g2_decap_8 FILLER_77_691 ();
 sg13g2_decap_8 FILLER_77_698 ();
 sg13g2_decap_8 FILLER_77_705 ();
 sg13g2_decap_8 FILLER_77_712 ();
 sg13g2_decap_8 FILLER_77_719 ();
 sg13g2_decap_8 FILLER_77_726 ();
 sg13g2_decap_8 FILLER_77_733 ();
 sg13g2_decap_8 FILLER_77_740 ();
 sg13g2_decap_8 FILLER_77_747 ();
 sg13g2_decap_8 FILLER_77_754 ();
 sg13g2_decap_8 FILLER_77_761 ();
 sg13g2_decap_8 FILLER_77_768 ();
 sg13g2_decap_8 FILLER_77_775 ();
 sg13g2_decap_8 FILLER_77_782 ();
 sg13g2_decap_8 FILLER_77_789 ();
 sg13g2_decap_8 FILLER_77_796 ();
 sg13g2_decap_8 FILLER_77_803 ();
 sg13g2_decap_8 FILLER_77_810 ();
 sg13g2_decap_8 FILLER_77_817 ();
 sg13g2_decap_8 FILLER_77_824 ();
 sg13g2_decap_8 FILLER_77_831 ();
 sg13g2_decap_8 FILLER_77_838 ();
 sg13g2_decap_8 FILLER_77_845 ();
 sg13g2_decap_8 FILLER_77_852 ();
 sg13g2_fill_2 FILLER_77_859 ();
 sg13g2_fill_1 FILLER_77_861 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_31 ();
 sg13g2_fill_2 FILLER_78_46 ();
 sg13g2_fill_2 FILLER_78_75 ();
 sg13g2_fill_1 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_216 ();
 sg13g2_fill_1 FILLER_78_266 ();
 sg13g2_fill_2 FILLER_78_272 ();
 sg13g2_fill_2 FILLER_78_282 ();
 sg13g2_fill_2 FILLER_78_294 ();
 sg13g2_fill_1 FILLER_78_296 ();
 sg13g2_fill_1 FILLER_78_342 ();
 sg13g2_fill_2 FILLER_78_353 ();
 sg13g2_fill_2 FILLER_78_392 ();
 sg13g2_fill_1 FILLER_78_394 ();
 sg13g2_fill_1 FILLER_78_406 ();
 sg13g2_fill_2 FILLER_78_433 ();
 sg13g2_fill_1 FILLER_78_435 ();
 sg13g2_fill_2 FILLER_78_465 ();
 sg13g2_fill_1 FILLER_78_499 ();
 sg13g2_decap_8 FILLER_78_549 ();
 sg13g2_decap_8 FILLER_78_556 ();
 sg13g2_decap_8 FILLER_78_563 ();
 sg13g2_decap_8 FILLER_78_570 ();
 sg13g2_decap_8 FILLER_78_577 ();
 sg13g2_decap_8 FILLER_78_584 ();
 sg13g2_decap_8 FILLER_78_591 ();
 sg13g2_decap_8 FILLER_78_598 ();
 sg13g2_decap_8 FILLER_78_605 ();
 sg13g2_decap_8 FILLER_78_612 ();
 sg13g2_decap_8 FILLER_78_619 ();
 sg13g2_decap_8 FILLER_78_626 ();
 sg13g2_decap_8 FILLER_78_633 ();
 sg13g2_decap_8 FILLER_78_640 ();
 sg13g2_decap_8 FILLER_78_647 ();
 sg13g2_decap_8 FILLER_78_654 ();
 sg13g2_decap_8 FILLER_78_661 ();
 sg13g2_decap_8 FILLER_78_668 ();
 sg13g2_decap_8 FILLER_78_675 ();
 sg13g2_decap_8 FILLER_78_682 ();
 sg13g2_decap_8 FILLER_78_689 ();
 sg13g2_decap_8 FILLER_78_696 ();
 sg13g2_decap_8 FILLER_78_703 ();
 sg13g2_decap_8 FILLER_78_710 ();
 sg13g2_decap_8 FILLER_78_717 ();
 sg13g2_decap_8 FILLER_78_724 ();
 sg13g2_decap_8 FILLER_78_731 ();
 sg13g2_decap_8 FILLER_78_738 ();
 sg13g2_decap_8 FILLER_78_745 ();
 sg13g2_decap_8 FILLER_78_752 ();
 sg13g2_decap_8 FILLER_78_759 ();
 sg13g2_decap_8 FILLER_78_766 ();
 sg13g2_decap_8 FILLER_78_773 ();
 sg13g2_decap_8 FILLER_78_780 ();
 sg13g2_decap_8 FILLER_78_787 ();
 sg13g2_decap_8 FILLER_78_794 ();
 sg13g2_decap_8 FILLER_78_801 ();
 sg13g2_decap_8 FILLER_78_808 ();
 sg13g2_decap_8 FILLER_78_815 ();
 sg13g2_decap_8 FILLER_78_822 ();
 sg13g2_decap_8 FILLER_78_829 ();
 sg13g2_decap_8 FILLER_78_836 ();
 sg13g2_decap_8 FILLER_78_843 ();
 sg13g2_decap_8 FILLER_78_850 ();
 sg13g2_decap_4 FILLER_78_857 ();
 sg13g2_fill_1 FILLER_78_861 ();
 sg13g2_fill_1 FILLER_79_27 ();
 sg13g2_fill_1 FILLER_79_125 ();
 sg13g2_fill_1 FILLER_79_280 ();
 sg13g2_fill_2 FILLER_79_311 ();
 sg13g2_fill_1 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_428 ();
 sg13g2_decap_8 FILLER_79_489 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_536 ();
 sg13g2_decap_8 FILLER_79_543 ();
 sg13g2_decap_8 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_557 ();
 sg13g2_decap_8 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_decap_8 FILLER_79_578 ();
 sg13g2_decap_8 FILLER_79_585 ();
 sg13g2_decap_8 FILLER_79_592 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_620 ();
 sg13g2_decap_8 FILLER_79_627 ();
 sg13g2_decap_8 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_683 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_4 FILLER_79_858 ();
 sg13g2_fill_1 FILLER_80_0 ();
 sg13g2_fill_1 FILLER_80_45 ();
 sg13g2_fill_2 FILLER_80_72 ();
 sg13g2_fill_1 FILLER_80_164 ();
 sg13g2_fill_1 FILLER_80_216 ();
 sg13g2_fill_2 FILLER_80_342 ();
 sg13g2_fill_1 FILLER_80_344 ();
 sg13g2_fill_2 FILLER_80_382 ();
 sg13g2_fill_1 FILLER_80_384 ();
 sg13g2_decap_8 FILLER_80_429 ();
 sg13g2_decap_4 FILLER_80_436 ();
 sg13g2_decap_4 FILLER_80_444 ();
 sg13g2_fill_1 FILLER_80_448 ();
 sg13g2_decap_4 FILLER_80_453 ();
 sg13g2_fill_1 FILLER_80_457 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_fill_2 FILLER_80_469 ();
 sg13g2_fill_1 FILLER_80_471 ();
 sg13g2_decap_4 FILLER_80_495 ();
 sg13g2_fill_2 FILLER_80_511 ();
 sg13g2_fill_1 FILLER_80_513 ();
 sg13g2_decap_8 FILLER_80_523 ();
 sg13g2_decap_8 FILLER_80_530 ();
 sg13g2_decap_8 FILLER_80_537 ();
 sg13g2_decap_8 FILLER_80_544 ();
 sg13g2_decap_8 FILLER_80_551 ();
 sg13g2_decap_8 FILLER_80_558 ();
 sg13g2_decap_8 FILLER_80_565 ();
 sg13g2_decap_8 FILLER_80_572 ();
 sg13g2_decap_8 FILLER_80_579 ();
 sg13g2_decap_8 FILLER_80_586 ();
 sg13g2_decap_8 FILLER_80_593 ();
 sg13g2_decap_8 FILLER_80_600 ();
 sg13g2_decap_8 FILLER_80_607 ();
 sg13g2_decap_8 FILLER_80_614 ();
 sg13g2_decap_8 FILLER_80_621 ();
 sg13g2_decap_8 FILLER_80_628 ();
 sg13g2_decap_8 FILLER_80_635 ();
 sg13g2_decap_8 FILLER_80_642 ();
 sg13g2_decap_8 FILLER_80_649 ();
 sg13g2_decap_8 FILLER_80_656 ();
 sg13g2_decap_8 FILLER_80_663 ();
 sg13g2_decap_8 FILLER_80_670 ();
 sg13g2_decap_8 FILLER_80_677 ();
 sg13g2_decap_8 FILLER_80_684 ();
 sg13g2_decap_8 FILLER_80_691 ();
 sg13g2_decap_8 FILLER_80_698 ();
 sg13g2_decap_8 FILLER_80_705 ();
 sg13g2_decap_8 FILLER_80_712 ();
 sg13g2_decap_8 FILLER_80_719 ();
 sg13g2_decap_8 FILLER_80_726 ();
 sg13g2_decap_8 FILLER_80_733 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_decap_8 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_754 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_768 ();
 sg13g2_decap_8 FILLER_80_775 ();
 sg13g2_decap_8 FILLER_80_782 ();
 sg13g2_decap_8 FILLER_80_789 ();
 sg13g2_decap_8 FILLER_80_796 ();
 sg13g2_decap_8 FILLER_80_803 ();
 sg13g2_decap_8 FILLER_80_810 ();
 sg13g2_decap_8 FILLER_80_817 ();
 sg13g2_decap_8 FILLER_80_824 ();
 sg13g2_decap_8 FILLER_80_831 ();
 sg13g2_decap_8 FILLER_80_838 ();
 sg13g2_decap_8 FILLER_80_845 ();
 sg13g2_decap_8 FILLER_80_852 ();
 sg13g2_fill_2 FILLER_80_859 ();
 sg13g2_fill_1 FILLER_80_861 ();
 assign uio_oe[0] = net48;
 assign uio_oe[1] = net49;
 assign uio_oe[2] = net50;
 assign uio_oe[3] = net14;
 assign uio_oe[4] = net51;
 assign uio_oe[5] = net52;
 assign uio_oe[6] = net53;
 assign uio_oe[7] = net54;
 assign uio_out[3] = net15;
endmodule
