module tt_um_spi_aggregator (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire adc_cs_n;
 wire \adc_data0[0] ;
 wire \adc_data0[10] ;
 wire \adc_data0[11] ;
 wire \adc_data0[12] ;
 wire \adc_data0[13] ;
 wire \adc_data0[14] ;
 wire \adc_data0[15] ;
 wire \adc_data0[1] ;
 wire \adc_data0[2] ;
 wire \adc_data0[3] ;
 wire \adc_data0[4] ;
 wire \adc_data0[5] ;
 wire \adc_data0[6] ;
 wire \adc_data0[7] ;
 wire \adc_data0[8] ;
 wire \adc_data0[9] ;
 wire \adc_data1[0] ;
 wire \adc_data1[10] ;
 wire \adc_data1[11] ;
 wire \adc_data1[12] ;
 wire \adc_data1[13] ;
 wire \adc_data1[14] ;
 wire \adc_data1[15] ;
 wire \adc_data1[1] ;
 wire \adc_data1[2] ;
 wire \adc_data1[3] ;
 wire \adc_data1[4] ;
 wire \adc_data1[5] ;
 wire \adc_data1[6] ;
 wire \adc_data1[7] ;
 wire \adc_data1[8] ;
 wire \adc_data1[9] ;
 wire \adc_data2[0] ;
 wire \adc_data2[10] ;
 wire \adc_data2[11] ;
 wire \adc_data2[12] ;
 wire \adc_data2[13] ;
 wire \adc_data2[14] ;
 wire \adc_data2[15] ;
 wire \adc_data2[1] ;
 wire \adc_data2[2] ;
 wire \adc_data2[3] ;
 wire \adc_data2[4] ;
 wire \adc_data2[5] ;
 wire \adc_data2[6] ;
 wire \adc_data2[7] ;
 wire \adc_data2[8] ;
 wire \adc_data2[9] ;
 wire \adc_data3[0] ;
 wire \adc_data3[10] ;
 wire \adc_data3[11] ;
 wire \adc_data3[12] ;
 wire \adc_data3[13] ;
 wire \adc_data3[14] ;
 wire \adc_data3[15] ;
 wire \adc_data3[1] ;
 wire \adc_data3[2] ;
 wire \adc_data3[3] ;
 wire \adc_data3[4] ;
 wire \adc_data3[5] ;
 wire \adc_data3[6] ;
 wire \adc_data3[7] ;
 wire \adc_data3[8] ;
 wire \adc_data3[9] ;
 wire adc_sclk;
 wire \clk_div[0] ;
 wire \clk_div[1] ;
 wire \clk_div[2] ;
 wire \clk_div[3] ;
 wire \cycle[0] ;
 wire \cycle[1] ;
 wire \cycle[2] ;
 wire \cycle[3] ;
 wire \cycle[4] ;
 wire \cycle[5] ;
 wire tx_cs_n;
 wire \tx_cycle[0] ;
 wire \tx_cycle[1] ;
 wire \tx_cycle[2] ;
 wire \tx_cycle[3] ;
 wire \tx_cycle[4] ;
 wire \tx_cycle[5] ;
 wire \tx_cycle[6] ;
 wire tx_mosi;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net103;
 wire net104;
 wire clk_regs;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_4_0_0_clk_regs;
 wire clknet_4_1_0_clk_regs;
 wire clknet_4_2_0_clk_regs;
 wire clknet_4_3_0_clk_regs;
 wire clknet_4_4_0_clk_regs;
 wire clknet_4_5_0_clk_regs;
 wire clknet_4_6_0_clk_regs;
 wire clknet_4_7_0_clk_regs;
 wire clknet_4_8_0_clk_regs;
 wire clknet_4_9_0_clk_regs;
 wire clknet_4_10_0_clk_regs;
 wire clknet_4_11_0_clk_regs;
 wire clknet_4_12_0_clk_regs;
 wire clknet_4_13_0_clk_regs;
 wire clknet_4_14_0_clk_regs;
 wire clknet_4_15_0_clk_regs;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;

 sg13g2_inv_1 _0904_ (.Y(_0087_),
    .A(net117));
 sg13g2_inv_1 _0905_ (.Y(_0088_),
    .A(net172));
 sg13g2_inv_1 _0906_ (.Y(_0089_),
    .A(net180));
 sg13g2_inv_1 _0907_ (.Y(_0090_),
    .A(net198));
 sg13g2_inv_1 _0908_ (.Y(_0091_),
    .A(net174));
 sg13g2_inv_1 _0909_ (.Y(_0092_),
    .A(net152));
 sg13g2_inv_1 _0910_ (.Y(_0093_),
    .A(net202));
 sg13g2_inv_1 _0911_ (.Y(_0094_),
    .A(net196));
 sg13g2_inv_1 _0912_ (.Y(_0095_),
    .A(net205));
 sg13g2_inv_1 _0913_ (.Y(_0096_),
    .A(net177));
 sg13g2_inv_1 _0914_ (.Y(_0097_),
    .A(net137));
 sg13g2_inv_2 _0915_ (.Y(_0098_),
    .A(net131));
 sg13g2_inv_1 _0916_ (.Y(_0099_),
    .A(net181));
 sg13g2_inv_1 _0917_ (.Y(_0100_),
    .A(net178));
 sg13g2_inv_1 _0918_ (.Y(_0101_),
    .A(net179));
 sg13g2_inv_1 _0919_ (.Y(_0102_),
    .A(net146));
 sg13g2_inv_1 _0920_ (.Y(_0103_),
    .A(net142));
 sg13g2_inv_1 _0921_ (.Y(_0104_),
    .A(net132));
 sg13g2_inv_1 _0922_ (.Y(_0105_),
    .A(net149));
 sg13g2_inv_2 _0923_ (.Y(_0106_),
    .A(net108));
 sg13g2_inv_1 _0924_ (.Y(_0107_),
    .A(net136));
 sg13g2_inv_1 _0925_ (.Y(_0108_),
    .A(net113));
 sg13g2_inv_1 _0926_ (.Y(_0109_),
    .A(net212));
 sg13g2_inv_1 _0927_ (.Y(_0110_),
    .A(net170));
 sg13g2_inv_1 _0928_ (.Y(_0111_),
    .A(net210));
 sg13g2_inv_1 _0929_ (.Y(_0112_),
    .A(net183));
 sg13g2_inv_1 _0930_ (.Y(_0113_),
    .A(net204));
 sg13g2_inv_1 _0931_ (.Y(_0114_),
    .A(net186));
 sg13g2_inv_1 _0932_ (.Y(_0115_),
    .A(net197));
 sg13g2_inv_1 _0933_ (.Y(_0116_),
    .A(net193));
 sg13g2_inv_1 _0934_ (.Y(_0117_),
    .A(net166));
 sg13g2_inv_1 _0935_ (.Y(_0118_),
    .A(net138));
 sg13g2_inv_2 _0936_ (.Y(_0119_),
    .A(net123));
 sg13g2_inv_1 _0937_ (.Y(_0120_),
    .A(net182));
 sg13g2_inv_1 _0938_ (.Y(_0121_),
    .A(net195));
 sg13g2_inv_1 _0939_ (.Y(_0122_),
    .A(net185));
 sg13g2_inv_1 _0940_ (.Y(_0123_),
    .A(net203));
 sg13g2_inv_1 _0941_ (.Y(_0124_),
    .A(net150));
 sg13g2_inv_1 _0942_ (.Y(_0125_),
    .A(net190));
 sg13g2_inv_1 _0943_ (.Y(_0126_),
    .A(net206));
 sg13g2_inv_1 _0944_ (.Y(_0127_),
    .A(net171));
 sg13g2_inv_1 _0945_ (.Y(_0128_),
    .A(net141));
 sg13g2_inv_1 _0946_ (.Y(_0129_),
    .A(net115));
 sg13g2_inv_1 _0947_ (.Y(_0130_),
    .A(net192));
 sg13g2_inv_1 _0948_ (.Y(_0131_),
    .A(net299));
 sg13g2_inv_2 _0949_ (.Y(_0132_),
    .A(\tx_cycle[5] ));
 sg13g2_inv_2 _0950_ (.Y(_0133_),
    .A(net300));
 sg13g2_inv_1 _0951_ (.Y(_0134_),
    .A(net301));
 sg13g2_inv_2 _0952_ (.Y(_0135_),
    .A(net302));
 sg13g2_inv_1 _0953_ (.Y(_0136_),
    .A(net213));
 sg13g2_inv_1 _0954_ (.Y(_0137_),
    .A(net105));
 sg13g2_inv_2 _0955_ (.Y(_0138_),
    .A(\cycle[1] ));
 sg13g2_inv_1 _0956_ (.Y(_0139_),
    .A(\cycle[0] ));
 sg13g2_inv_4 _0957_ (.A(net328),
    .Y(_0140_));
 sg13g2_inv_1 _0958_ (.Y(_0141_),
    .A(net354));
 sg13g2_inv_1 _0959_ (.Y(_0142_),
    .A(net5));
 sg13g2_inv_1 _0960_ (.Y(_0143_),
    .A(net8));
 sg13g2_inv_1 _0961_ (.Y(_0144_),
    .A(net7));
 sg13g2_inv_1 _0962_ (.Y(_0145_),
    .A(net6));
 sg13g2_inv_1 _0963_ (.Y(_0146_),
    .A(net9));
 sg13g2_inv_1 _0964_ (.Y(_0147_),
    .A(net379));
 sg13g2_nand2_2 _0965_ (.Y(_0148_),
    .A(net359),
    .B(net375));
 sg13g2_and3_2 _0966_ (.X(_0149_),
    .A(net338),
    .B(net348),
    .C(net364));
 sg13g2_xnor2_1 _0967_ (.Y(_0150_),
    .A(net346),
    .B(_0148_));
 sg13g2_xor2_1 _0968_ (.B(_0148_),
    .A(net346),
    .X(_0151_));
 sg13g2_xor2_1 _0969_ (.B(net377),
    .A(net359),
    .X(_0152_));
 sg13g2_nand2_1 _0970_ (.Y(_0153_),
    .A(net3),
    .B(_0152_));
 sg13g2_nand2b_1 _0971_ (.Y(_0154_),
    .B(net2),
    .A_N(net377));
 sg13g2_xnor2_1 _0972_ (.Y(_0155_),
    .A(net3),
    .B(_0152_));
 sg13g2_o21ai_1 _0973_ (.B1(_0153_),
    .Y(_0156_),
    .A1(_0154_),
    .A2(_0155_));
 sg13g2_and3_1 _0974_ (.X(_0157_),
    .A(net335),
    .B(_0150_),
    .C(_0156_));
 sg13g2_nand3_1 _0975_ (.B(_0150_),
    .C(_0156_),
    .A(net335),
    .Y(_0158_));
 sg13g2_nand2_2 _0976_ (.Y(_0159_),
    .A(net331),
    .B(net338));
 sg13g2_nor2_2 _0977_ (.A(_0148_),
    .B(net311),
    .Y(_0160_));
 sg13g2_nand2_2 _0978_ (.Y(_0161_),
    .A(net335),
    .B(_0149_));
 sg13g2_or2_1 _0979_ (.X(_0162_),
    .B(_0149_),
    .A(net335));
 sg13g2_xnor2_1 _0980_ (.Y(_0163_),
    .A(net335),
    .B(_0149_));
 sg13g2_inv_1 _0981_ (.Y(_0164_),
    .A(net298));
 sg13g2_a21oi_1 _0982_ (.A1(_0150_),
    .A2(_0156_),
    .Y(_0165_),
    .B1(_0164_));
 sg13g2_o21ai_1 _0983_ (.B1(\cycle[3] ),
    .Y(_0166_),
    .A1(_0157_),
    .A2(_0165_));
 sg13g2_xnor2_1 _0984_ (.Y(_0167_),
    .A(_0150_),
    .B(_0156_));
 sg13g2_nand2_1 _0985_ (.Y(_0168_),
    .A(\cycle[2] ),
    .B(_0167_));
 sg13g2_nand2_1 _0986_ (.Y(_0169_),
    .A(\cycle[1] ),
    .B(_0155_));
 sg13g2_xor2_1 _0987_ (.B(_0155_),
    .A(_0154_),
    .X(_0170_));
 sg13g2_xor2_1 _0988_ (.B(net2),
    .A(net377),
    .X(_0171_));
 sg13g2_nor2_1 _0989_ (.A(\cycle[0] ),
    .B(_0171_),
    .Y(_0172_));
 sg13g2_a22oi_1 _0990_ (.Y(_0173_),
    .B1(_0172_),
    .B2(_0169_),
    .A2(_0170_),
    .A1(_0138_));
 sg13g2_o21ai_1 _0991_ (.B1(_0173_),
    .Y(_0174_),
    .A1(\cycle[2] ),
    .A2(_0167_));
 sg13g2_nand3_1 _0992_ (.B(_0168_),
    .C(_0174_),
    .A(_0166_),
    .Y(_0175_));
 sg13g2_nor3_1 _0993_ (.A(\cycle[3] ),
    .B(_0157_),
    .C(_0165_),
    .Y(_0176_));
 sg13g2_or3_1 _0994_ (.A(\cycle[3] ),
    .B(_0157_),
    .C(_0165_),
    .X(_0177_));
 sg13g2_and3_1 _0995_ (.X(_0178_),
    .A(\cycle[4] ),
    .B(_0158_),
    .C(_0161_));
 sg13g2_a21oi_1 _0996_ (.A1(_0158_),
    .A2(_0161_),
    .Y(_0179_),
    .B1(\cycle[4] ));
 sg13g2_or2_1 _0997_ (.X(_0180_),
    .B(_0179_),
    .A(_0178_));
 sg13g2_nor3_1 _0998_ (.A(_0176_),
    .B(_0178_),
    .C(_0179_),
    .Y(_0181_));
 sg13g2_or2_1 _0999_ (.X(_0182_),
    .B(_0178_),
    .A(\cycle[5] ));
 sg13g2_a21oi_2 _1000_ (.B1(_0182_),
    .Y(_0183_),
    .A2(_0181_),
    .A1(_0175_));
 sg13g2_inv_1 _1001_ (.Y(adc_cs_n),
    .A(net297));
 sg13g2_a21oi_1 _1002_ (.A1(\tx_cycle[5] ),
    .A2(_0161_),
    .Y(_0184_),
    .B1(\tx_cycle[6] ));
 sg13g2_nor2_1 _1003_ (.A(_0135_),
    .B(net375),
    .Y(_0185_));
 sg13g2_nor2_2 _1004_ (.A(net322),
    .B(net364),
    .Y(_0186_));
 sg13g2_nand2_1 _1005_ (.Y(_0187_),
    .A(net301),
    .B(net302));
 sg13g2_nor3_1 _1006_ (.A(\tx_cycle[3] ),
    .B(net359),
    .C(_0185_),
    .Y(_0188_));
 sg13g2_o21ai_1 _1007_ (.B1(_0187_),
    .Y(_0189_),
    .A1(_0186_),
    .A2(_0188_));
 sg13g2_o21ai_1 _1008_ (.B1(_0189_),
    .Y(_0190_),
    .A1(net300),
    .A2(_0151_));
 sg13g2_a221oi_1 _1009_ (.B2(\tx_cycle[5] ),
    .C1(\tx_cycle[6] ),
    .B1(net298),
    .A1(net300),
    .Y(_0191_),
    .A2(_0151_));
 sg13g2_a22oi_1 _1010_ (.Y(_0192_),
    .B1(_0190_),
    .B2(_0191_),
    .A2(_0184_),
    .A1(_0162_));
 sg13g2_nor2_2 _1011_ (.A(_0183_),
    .B(_0192_),
    .Y(_0193_));
 sg13g2_inv_2 _1012_ (.Y(tx_cs_n),
    .A(net295));
 sg13g2_nor2b_1 _1013_ (.A(net369),
    .B_N(net341),
    .Y(_0194_));
 sg13g2_xnor2_1 _1014_ (.Y(_0195_),
    .A(net341),
    .B(net369));
 sg13g2_xor2_1 _1015_ (.B(net375),
    .A(net346),
    .X(_0196_));
 sg13g2_nor2_2 _1016_ (.A(net303),
    .B(net375),
    .Y(_0197_));
 sg13g2_nor3_1 _1017_ (.A(net303),
    .B(\tx_cycle[0] ),
    .C(net375),
    .Y(_0198_));
 sg13g2_nand2_1 _1018_ (.Y(_0199_),
    .A(net303),
    .B(\tx_cycle[0] ));
 sg13g2_o21ai_1 _1019_ (.B1(net303),
    .Y(_0200_),
    .A1(\tx_cycle[0] ),
    .A2(net377));
 sg13g2_a21oi_1 _1020_ (.A1(net324),
    .A2(_0200_),
    .Y(_0201_),
    .B1(_0198_));
 sg13g2_a21oi_1 _1021_ (.A1(net302),
    .A2(_0195_),
    .Y(_0202_),
    .B1(_0201_));
 sg13g2_xor2_1 _1022_ (.B(net353),
    .A(net331),
    .X(_0203_));
 sg13g2_xnor2_1 _1023_ (.Y(_0204_),
    .A(_0194_),
    .B(_0203_));
 sg13g2_nand2_1 _1024_ (.Y(_0205_),
    .A(_0135_),
    .B(_0196_));
 sg13g2_o21ai_1 _1025_ (.B1(_0205_),
    .Y(_0206_),
    .A1(net301),
    .A2(_0204_));
 sg13g2_or2_1 _1026_ (.X(_0207_),
    .B(_0206_),
    .A(_0202_));
 sg13g2_o21ai_1 _1027_ (.B1(net341),
    .Y(_0208_),
    .A1(net353),
    .A2(net369));
 sg13g2_and2_1 _1028_ (.A(net326),
    .B(_0208_),
    .X(_0209_));
 sg13g2_o21ai_1 _1029_ (.B1(net331),
    .Y(_0210_),
    .A1(net341),
    .A2(net353));
 sg13g2_nor2_1 _1030_ (.A(_0149_),
    .B(_0210_),
    .Y(_0211_));
 sg13g2_nor2_1 _1031_ (.A(_0209_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_or2_1 _1032_ (.X(_0213_),
    .B(_0211_),
    .A(_0209_));
 sg13g2_a22oi_1 _1033_ (.Y(_0214_),
    .B1(_0213_),
    .B2(net300),
    .A2(_0204_),
    .A1(net301));
 sg13g2_nor2_1 _1034_ (.A(\tx_cycle[5] ),
    .B(_0210_),
    .Y(_0215_));
 sg13g2_a221oi_1 _1035_ (.B2(_0207_),
    .C1(_0215_),
    .B1(_0214_),
    .A1(_0133_),
    .Y(_0216_),
    .A2(_0212_));
 sg13g2_a21oi_1 _1036_ (.A1(\tx_cycle[5] ),
    .A2(_0210_),
    .Y(_0217_),
    .B1(\tx_cycle[6] ));
 sg13g2_nor2b_2 _1037_ (.A(_0216_),
    .B_N(_0217_),
    .Y(_0218_));
 sg13g2_inv_1 _1038_ (.Y(_0219_),
    .A(_0218_));
 sg13g2_nor2_1 _1039_ (.A(\adc_data3[15] ),
    .B(_0218_),
    .Y(_0220_));
 sg13g2_o21ai_1 _1040_ (.B1(_0135_),
    .Y(_0221_),
    .A1(_0152_),
    .A2(_0197_));
 sg13g2_a22oi_1 _1041_ (.Y(_0222_),
    .B1(_0197_),
    .B2(net359),
    .A2(_0150_),
    .A1(_0134_));
 sg13g2_and2_1 _1042_ (.A(net300),
    .B(_0163_),
    .X(_0223_));
 sg13g2_a221oi_1 _1043_ (.B2(_0222_),
    .C1(_0223_),
    .B1(_0221_),
    .A1(net301),
    .Y(_0224_),
    .A2(_0151_));
 sg13g2_nand2_1 _1044_ (.Y(_0225_),
    .A(_0132_),
    .B(_0160_));
 sg13g2_o21ai_1 _1045_ (.B1(_0225_),
    .Y(_0226_),
    .A1(net300),
    .A2(net298));
 sg13g2_o21ai_1 _1046_ (.B1(_0184_),
    .Y(_0227_),
    .A1(_0224_),
    .A2(_0226_));
 sg13g2_o21ai_1 _1047_ (.B1(_0227_),
    .Y(_0228_),
    .A1(\adc_data2[15] ),
    .A2(_0219_));
 sg13g2_o21ai_1 _1048_ (.B1(_0200_),
    .Y(_0229_),
    .A1(_0152_),
    .A2(_0198_));
 sg13g2_o21ai_1 _1049_ (.B1(_0229_),
    .Y(_0230_),
    .A1(net302),
    .A2(_0151_));
 sg13g2_a22oi_1 _1050_ (.Y(_0231_),
    .B1(net298),
    .B2(net301),
    .A2(_0151_),
    .A1(\tx_cycle[2] ));
 sg13g2_nor2_1 _1051_ (.A(\tx_cycle[3] ),
    .B(net298),
    .Y(_0232_));
 sg13g2_a221oi_1 _1052_ (.B2(_0231_),
    .C1(_0232_),
    .B1(_0230_),
    .A1(_0133_),
    .Y(_0233_),
    .A2(_0160_));
 sg13g2_o21ai_1 _1053_ (.B1(_0132_),
    .Y(_0234_),
    .A1(_0133_),
    .A2(_0160_));
 sg13g2_nor3_2 _1054_ (.A(\tx_cycle[6] ),
    .B(_0233_),
    .C(_0234_),
    .Y(_0235_));
 sg13g2_inv_1 _1055_ (.Y(_0236_),
    .A(_0235_));
 sg13g2_nor2_1 _1056_ (.A(_0227_),
    .B(_0235_),
    .Y(_0237_));
 sg13g2_or2_1 _1057_ (.X(_0238_),
    .B(_0235_),
    .A(_0227_));
 sg13g2_a22oi_1 _1058_ (.Y(_0239_),
    .B1(_0237_),
    .B2(\adc_data1[15] ),
    .A2(_0235_),
    .A1(\adc_data0[15] ));
 sg13g2_o21ai_1 _1059_ (.B1(_0239_),
    .Y(tx_mosi),
    .A1(_0220_),
    .A2(_0228_));
 sg13g2_a21oi_1 _1060_ (.A1(\clk_div[2] ),
    .A2(_0142_),
    .Y(_0240_),
    .B1(\clk_div[3] ));
 sg13g2_nand2b_1 _1061_ (.Y(_0241_),
    .B(net5),
    .A_N(\clk_div[2] ));
 sg13g2_xnor2_1 _1062_ (.Y(_0242_),
    .A(\clk_div[1] ),
    .B(net4));
 sg13g2_nand4_1 _1063_ (.B(_0240_),
    .C(_0241_),
    .A(net194),
    .Y(_0243_),
    .D(_0242_));
 sg13g2_and2_1 _1064_ (.A(net297),
    .B(_0243_),
    .X(_0244_));
 sg13g2_nand2_1 _1065_ (.Y(_0245_),
    .A(net297),
    .B(_0243_));
 sg13g2_nand2_1 _1066_ (.Y(_0246_),
    .A(net296),
    .B(_0192_));
 sg13g2_nor2_2 _1067_ (.A(net296),
    .B(_0243_),
    .Y(_0247_));
 sg13g2_or2_1 _1068_ (.X(_0248_),
    .B(_0243_),
    .A(net296));
 sg13g2_a22oi_1 _1069_ (.Y(_0249_),
    .B1(_0246_),
    .B2(_0248_),
    .A2(net297),
    .A1(_0131_));
 sg13g2_nand2_2 _1070_ (.Y(_0250_),
    .A(net379),
    .B(_0246_));
 sg13g2_xnor2_1 _1071_ (.Y(_0251_),
    .A(net211),
    .B(_0249_));
 sg13g2_nor2_1 _1072_ (.A(_0250_),
    .B(_0251_),
    .Y(_0000_));
 sg13g2_a21oi_1 _1073_ (.A1(\cycle[0] ),
    .A2(_0249_),
    .Y(_0252_),
    .B1(net128));
 sg13g2_nand3_1 _1074_ (.B(\cycle[0] ),
    .C(_0249_),
    .A(net128),
    .Y(_0253_));
 sg13g2_nand2b_1 _1075_ (.Y(_0254_),
    .B(_0253_),
    .A_N(_0250_));
 sg13g2_nor2_1 _1076_ (.A(net129),
    .B(_0254_),
    .Y(_0001_));
 sg13g2_nor2b_1 _1077_ (.A(net207),
    .B_N(_0253_),
    .Y(_0255_));
 sg13g2_and4_1 _1078_ (.A(net207),
    .B(net128),
    .C(\cycle[0] ),
    .D(_0249_),
    .X(_0256_));
 sg13g2_nor3_1 _1079_ (.A(_0250_),
    .B(net208),
    .C(_0256_),
    .Y(_0002_));
 sg13g2_xnor2_1 _1080_ (.Y(_0257_),
    .A(net200),
    .B(_0256_));
 sg13g2_nor2_1 _1081_ (.A(_0250_),
    .B(net201),
    .Y(_0003_));
 sg13g2_a21oi_1 _1082_ (.A1(\cycle[3] ),
    .A2(_0256_),
    .Y(_0258_),
    .B1(net110));
 sg13g2_nor2_1 _1083_ (.A(_0250_),
    .B(net111),
    .Y(_0004_));
 sg13g2_nor3_1 _1084_ (.A(_0137_),
    .B(net320),
    .C(_0249_),
    .Y(_0005_));
 sg13g2_nor2b_1 _1085_ (.A(_0170_),
    .B_N(_0171_),
    .Y(_0259_));
 sg13g2_nand2b_1 _1086_ (.Y(_0260_),
    .B(_0171_),
    .A_N(_0170_));
 sg13g2_nor2_1 _1087_ (.A(net311),
    .B(_0260_),
    .Y(_0261_));
 sg13g2_xnor2_1 _1088_ (.Y(_0262_),
    .A(_0180_),
    .B(_0261_));
 sg13g2_and2_1 _1089_ (.A(_0166_),
    .B(_0177_),
    .X(_0263_));
 sg13g2_nand2_1 _1090_ (.Y(_0264_),
    .A(_0167_),
    .B(_0259_));
 sg13g2_xnor2_1 _1091_ (.Y(_0265_),
    .A(_0263_),
    .B(_0264_));
 sg13g2_xor2_1 _1092_ (.B(_0167_),
    .A(\cycle[2] ),
    .X(_0266_));
 sg13g2_xnor2_1 _1093_ (.Y(_0267_),
    .A(\cycle[2] ),
    .B(_0167_));
 sg13g2_xnor2_1 _1094_ (.Y(_0268_),
    .A(_0138_),
    .B(_0170_));
 sg13g2_nand2_1 _1095_ (.Y(_0269_),
    .A(\cycle[0] ),
    .B(_0171_));
 sg13g2_o21ai_1 _1096_ (.B1(net299),
    .Y(_0270_),
    .A1(_0172_),
    .A2(_0268_));
 sg13g2_a21oi_1 _1097_ (.A1(_0259_),
    .A2(_0266_),
    .Y(_0271_),
    .B1(_0270_));
 sg13g2_a221oi_1 _1098_ (.B2(_0269_),
    .C1(\cycle[5] ),
    .B1(_0268_),
    .A1(_0260_),
    .Y(_0272_),
    .A2(_0267_));
 sg13g2_and2_1 _1099_ (.A(_0271_),
    .B(_0272_),
    .X(_0273_));
 sg13g2_and3_2 _1100_ (.X(_0274_),
    .A(_0262_),
    .B(_0265_),
    .C(_0273_));
 sg13g2_nand3_1 _1101_ (.B(_0265_),
    .C(_0273_),
    .A(_0262_),
    .Y(_0275_));
 sg13g2_o21ai_1 _1102_ (.B1(_0245_),
    .Y(_0276_),
    .A1(net296),
    .A2(net294));
 sg13g2_o21ai_1 _1103_ (.B1(net380),
    .Y(_0277_),
    .A1(_0136_),
    .A2(_0276_));
 sg13g2_a21oi_1 _1104_ (.A1(_0136_),
    .A2(tx_cs_n),
    .Y(_0006_),
    .B1(_0277_));
 sg13g2_xnor2_1 _1105_ (.Y(_0278_),
    .A(net303),
    .B(net213));
 sg13g2_inv_1 _1106_ (.Y(_0279_),
    .A(_0278_));
 sg13g2_a22oi_1 _1107_ (.Y(_0280_),
    .B1(_0279_),
    .B2(net295),
    .A2(_0276_),
    .A1(net303));
 sg13g2_nor2_1 _1108_ (.A(net321),
    .B(_0280_),
    .Y(_0007_));
 sg13g2_and3_2 _1109_ (.X(_0281_),
    .A(net302),
    .B(net303),
    .C(\tx_cycle[0] ));
 sg13g2_a21oi_1 _1110_ (.A1(\tx_cycle[1] ),
    .A2(\tx_cycle[0] ),
    .Y(_0282_),
    .B1(net302));
 sg13g2_nor2_2 _1111_ (.A(_0281_),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_a22oi_1 _1112_ (.Y(_0284_),
    .B1(_0283_),
    .B2(net295),
    .A2(_0276_),
    .A1(net302));
 sg13g2_nor2_1 _1113_ (.A(net317),
    .B(_0284_),
    .Y(_0008_));
 sg13g2_nand4_1 _1114_ (.B(net302),
    .C(net303),
    .A(net301),
    .Y(_0285_),
    .D(\tx_cycle[0] ));
 sg13g2_xnor2_1 _1115_ (.Y(_0286_),
    .A(_0134_),
    .B(_0281_));
 sg13g2_inv_1 _1116_ (.Y(_0287_),
    .A(_0286_));
 sg13g2_a22oi_1 _1117_ (.Y(_0288_),
    .B1(_0286_),
    .B2(net295),
    .A2(_0276_),
    .A1(net301));
 sg13g2_nor2_1 _1118_ (.A(net317),
    .B(_0288_),
    .Y(_0009_));
 sg13g2_or2_1 _1119_ (.X(_0289_),
    .B(_0285_),
    .A(_0133_));
 sg13g2_xnor2_1 _1120_ (.Y(_0290_),
    .A(net300),
    .B(_0285_));
 sg13g2_xnor2_1 _1121_ (.Y(_0291_),
    .A(_0133_),
    .B(_0285_));
 sg13g2_a22oi_1 _1122_ (.Y(_0292_),
    .B1(_0290_),
    .B2(net295),
    .A2(_0276_),
    .A1(net300));
 sg13g2_nor2_1 _1123_ (.A(net317),
    .B(_0292_),
    .Y(_0010_));
 sg13g2_nor2_1 _1124_ (.A(_0132_),
    .B(_0289_),
    .Y(_0293_));
 sg13g2_xnor2_1 _1125_ (.Y(_0294_),
    .A(\tx_cycle[5] ),
    .B(_0289_));
 sg13g2_xnor2_1 _1126_ (.Y(_0295_),
    .A(_0132_),
    .B(_0289_));
 sg13g2_a22oi_1 _1127_ (.Y(_0296_),
    .B1(_0294_),
    .B2(net295),
    .A2(_0276_),
    .A1(net217));
 sg13g2_nor2_1 _1128_ (.A(net317),
    .B(_0296_),
    .Y(_0011_));
 sg13g2_a22oi_1 _1129_ (.Y(_0297_),
    .B1(_0293_),
    .B2(net295),
    .A2(_0276_),
    .A1(net214));
 sg13g2_nor2_1 _1130_ (.A(net317),
    .B(net215),
    .Y(_0012_));
 sg13g2_nand3_1 _1131_ (.B(tx_cs_n),
    .C(_0245_),
    .A(net299),
    .Y(_0298_));
 sg13g2_o21ai_1 _1132_ (.B1(_0298_),
    .Y(_0299_),
    .A1(net299),
    .A2(_0247_));
 sg13g2_nor2_1 _1133_ (.A(net320),
    .B(net223),
    .Y(_0013_));
 sg13g2_xnor2_1 _1134_ (.Y(_0300_),
    .A(net194),
    .B(net297));
 sg13g2_nor2_1 _1135_ (.A(_0250_),
    .B(_0300_),
    .Y(_0014_));
 sg13g2_xor2_1 _1136_ (.B(net194),
    .A(net199),
    .X(_0301_));
 sg13g2_a22oi_1 _1137_ (.Y(_0302_),
    .B1(_0244_),
    .B2(_0301_),
    .A2(_0193_),
    .A1(net199));
 sg13g2_nor2_1 _1138_ (.A(net320),
    .B(_0302_),
    .Y(_0015_));
 sg13g2_nand3_1 _1139_ (.B(\clk_div[1] ),
    .C(\clk_div[0] ),
    .A(net175),
    .Y(_0303_));
 sg13g2_a21o_1 _1140_ (.A2(\clk_div[0] ),
    .A1(\clk_div[1] ),
    .B1(net175),
    .X(_0304_));
 sg13g2_and2_1 _1141_ (.A(_0303_),
    .B(_0304_),
    .X(_0305_));
 sg13g2_a22oi_1 _1142_ (.Y(_0306_),
    .B1(_0244_),
    .B2(_0305_),
    .A2(_0193_),
    .A1(net175));
 sg13g2_nor2_1 _1143_ (.A(net320),
    .B(net176),
    .Y(_0016_));
 sg13g2_xnor2_1 _1144_ (.Y(_0307_),
    .A(net188),
    .B(_0303_));
 sg13g2_a22oi_1 _1145_ (.Y(_0308_),
    .B1(_0244_),
    .B2(_0307_),
    .A2(net295),
    .A1(net188));
 sg13g2_nor2_1 _1146_ (.A(net320),
    .B(net189),
    .Y(_0017_));
 sg13g2_nand2b_1 _1147_ (.Y(_0309_),
    .B(_0295_),
    .A_N(_0210_));
 sg13g2_o21ai_1 _1148_ (.B1(net324),
    .Y(_0310_),
    .A1(_0197_),
    .A2(_0278_));
 sg13g2_or2_1 _1149_ (.X(_0311_),
    .B(_0199_),
    .A(net375));
 sg13g2_o21ai_1 _1150_ (.B1(_0196_),
    .Y(_0312_),
    .A1(_0281_),
    .A2(_0282_));
 sg13g2_nand3_1 _1151_ (.B(_0311_),
    .C(_0312_),
    .A(_0310_),
    .Y(_0313_));
 sg13g2_a22oi_1 _1152_ (.Y(_0314_),
    .B1(_0286_),
    .B2(_0204_),
    .A2(_0283_),
    .A1(_0195_));
 sg13g2_nor2_1 _1153_ (.A(_0204_),
    .B(_0286_),
    .Y(_0315_));
 sg13g2_a221oi_1 _1154_ (.B2(_0314_),
    .C1(_0315_),
    .B1(_0313_),
    .A1(_0212_),
    .Y(_0316_),
    .A2(_0291_));
 sg13g2_a22oi_1 _1155_ (.Y(_0317_),
    .B1(_0294_),
    .B2(_0210_),
    .A2(_0290_),
    .A1(_0213_));
 sg13g2_nand2b_1 _1156_ (.Y(_0318_),
    .B(_0317_),
    .A_N(_0316_));
 sg13g2_o21ai_1 _1157_ (.B1(_0152_),
    .Y(_0319_),
    .A1(_0281_),
    .A2(_0282_));
 sg13g2_o21ai_1 _1158_ (.B1(_0319_),
    .Y(_0320_),
    .A1(net375),
    .A2(_0279_));
 sg13g2_a22oi_1 _1159_ (.Y(_0321_),
    .B1(_0286_),
    .B2(_0151_),
    .A2(_0283_),
    .A1(net324));
 sg13g2_nor2_1 _1160_ (.A(net298),
    .B(_0290_),
    .Y(_0322_));
 sg13g2_a221oi_1 _1161_ (.B2(_0321_),
    .C1(_0322_),
    .B1(_0320_),
    .A1(_0150_),
    .Y(_0323_),
    .A2(_0287_));
 sg13g2_a221oi_1 _1162_ (.B2(_0161_),
    .C1(_0323_),
    .B1(_0294_),
    .A1(net298),
    .Y(_0324_),
    .A2(_0290_));
 sg13g2_a221oi_1 _1163_ (.B2(_0318_),
    .C1(_0324_),
    .B1(_0309_),
    .A1(_0160_),
    .Y(_0325_),
    .A2(_0295_));
 sg13g2_nor3_1 _1164_ (.A(_0161_),
    .B(_0290_),
    .C(_0294_),
    .Y(_0326_));
 sg13g2_nand2_1 _1165_ (.Y(_0327_),
    .A(_0164_),
    .B(_0287_));
 sg13g2_o21ai_1 _1166_ (.B1(_0152_),
    .Y(_0328_),
    .A1(_0197_),
    .A2(_0278_));
 sg13g2_nor2_1 _1167_ (.A(_0151_),
    .B(_0283_),
    .Y(_0329_));
 sg13g2_nand2_1 _1168_ (.Y(_0330_),
    .A(_0311_),
    .B(_0328_));
 sg13g2_a22oi_1 _1169_ (.Y(_0331_),
    .B1(_0286_),
    .B2(net298),
    .A2(_0283_),
    .A1(_0151_));
 sg13g2_o21ai_1 _1170_ (.B1(_0331_),
    .Y(_0332_),
    .A1(_0329_),
    .A2(_0330_));
 sg13g2_a221oi_1 _1171_ (.B2(_0332_),
    .C1(_0294_),
    .B1(_0327_),
    .A1(_0161_),
    .Y(_0333_),
    .A2(_0290_));
 sg13g2_or2_1 _1172_ (.X(_0334_),
    .B(_0333_),
    .A(_0326_));
 sg13g2_xnor2_1 _1173_ (.Y(_0335_),
    .A(\tx_cycle[6] ),
    .B(_0293_));
 sg13g2_o21ai_1 _1174_ (.B1(_0335_),
    .Y(_0336_),
    .A1(_0325_),
    .A2(_0334_));
 sg13g2_nand2_1 _1175_ (.Y(_0337_),
    .A(_0218_),
    .B(_0238_));
 sg13g2_xor2_1 _1176_ (.B(_0337_),
    .A(_0336_),
    .X(_0338_));
 sg13g2_nand2_1 _1177_ (.Y(_0339_),
    .A(\tx_cycle[5] ),
    .B(_0140_));
 sg13g2_xor2_1 _1178_ (.B(net359),
    .A(\tx_cycle[3] ),
    .X(_0340_));
 sg13g2_a22oi_1 _1179_ (.Y(_0341_),
    .B1(net375),
    .B2(_0135_),
    .A2(net335),
    .A1(_0132_));
 sg13g2_xnor2_1 _1180_ (.Y(_0342_),
    .A(\tx_cycle[4] ),
    .B(net346));
 sg13g2_nand3_1 _1181_ (.B(_0341_),
    .C(_0342_),
    .A(_0339_),
    .Y(_0343_));
 sg13g2_nor4_1 _1182_ (.A(_0185_),
    .B(_0199_),
    .C(_0340_),
    .D(_0343_),
    .Y(_0344_));
 sg13g2_or3_1 _1183_ (.A(tx_cs_n),
    .B(_0338_),
    .C(_0344_),
    .X(_0345_));
 sg13g2_mux2_1 _1184_ (.A0(_0235_),
    .A1(_0247_),
    .S(_0345_),
    .X(_0346_));
 sg13g2_mux2_1 _1185_ (.A0(_0236_),
    .A1(_0248_),
    .S(_0345_),
    .X(_0347_));
 sg13g2_a22oi_1 _1186_ (.Y(_0348_),
    .B1(net2),
    .B2(_0139_),
    .A2(net3),
    .A1(_0138_));
 sg13g2_nor4_1 _1187_ (.A(\cycle[5] ),
    .B(\cycle[4] ),
    .C(\cycle[3] ),
    .D(\cycle[2] ),
    .Y(_0349_));
 sg13g2_o21ai_1 _1188_ (.B1(_0349_),
    .Y(_0350_),
    .A1(_0138_),
    .A2(net3));
 sg13g2_nor2_2 _1189_ (.A(_0348_),
    .B(_0350_),
    .Y(_0351_));
 sg13g2_inv_1 _1190_ (.Y(_0352_),
    .A(_0351_));
 sg13g2_nor3_2 _1191_ (.A(net224),
    .B(net296),
    .C(_0351_),
    .Y(_0353_));
 sg13g2_a21oi_1 _1192_ (.A1(net270),
    .A2(net281),
    .Y(_0354_),
    .B1(net126));
 sg13g2_o21ai_1 _1193_ (.B1(net297),
    .Y(_0355_),
    .A1(_0160_),
    .A2(net287));
 sg13g2_a21oi_1 _1194_ (.A1(_0145_),
    .A2(net281),
    .Y(_0356_),
    .B1(_0355_));
 sg13g2_o21ai_1 _1195_ (.B1(net380),
    .Y(_0357_),
    .A1(_0347_),
    .A2(_0356_));
 sg13g2_nor2_1 _1196_ (.A(net127),
    .B(_0357_),
    .Y(_0018_));
 sg13g2_a21oi_1 _1197_ (.A1(_0131_),
    .A2(_0352_),
    .Y(_0358_),
    .B1(net296));
 sg13g2_o21ai_1 _1198_ (.B1(net297),
    .Y(_0359_),
    .A1(adc_sclk),
    .A2(_0351_));
 sg13g2_nor2_2 _1199_ (.A(net288),
    .B(net282),
    .Y(_0360_));
 sg13g2_nand2_2 _1200_ (.Y(_0361_),
    .A(net286),
    .B(net275));
 sg13g2_nand2_2 _1201_ (.Y(_0362_),
    .A(net270),
    .B(_0361_));
 sg13g2_nor2_1 _1202_ (.A(\adc_data0[0] ),
    .B(net367),
    .Y(_0363_));
 sg13g2_a21oi_1 _1203_ (.A1(_0130_),
    .A2(net367),
    .Y(_0364_),
    .B1(_0363_));
 sg13g2_and2_1 _1204_ (.A(net350),
    .B(_0364_),
    .X(_0365_));
 sg13g2_nand3_1 _1205_ (.B(net340),
    .C(_0365_),
    .A(net329),
    .Y(_0366_));
 sg13g2_nand2_1 _1206_ (.Y(_0367_),
    .A(net290),
    .B(_0366_));
 sg13g2_o21ai_1 _1207_ (.B1(_0367_),
    .Y(_0368_),
    .A1(net126),
    .A2(net277));
 sg13g2_a221oi_1 _1208_ (.B2(net269),
    .C1(net316),
    .B1(_0368_),
    .A1(_0130_),
    .Y(_0019_),
    .A2(_0362_));
 sg13g2_and2_1 _1209_ (.A(\adc_data0[0] ),
    .B(net367),
    .X(_0369_));
 sg13g2_mux2_1 _1210_ (.A0(_0130_),
    .A1(_0129_),
    .S(net367),
    .X(_0370_));
 sg13g2_nor2_1 _1211_ (.A(net351),
    .B(_0369_),
    .Y(_0371_));
 sg13g2_a21oi_1 _1212_ (.A1(net351),
    .A2(_0370_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_and2_1 _1213_ (.A(net340),
    .B(_0372_),
    .X(_0373_));
 sg13g2_nor2_2 _1214_ (.A(net326),
    .B(net286),
    .Y(_0374_));
 sg13g2_a22oi_1 _1215_ (.Y(_0375_),
    .B1(_0373_),
    .B2(_0374_),
    .A2(net283),
    .A1(\adc_data0[1] ));
 sg13g2_nand2b_1 _1216_ (.Y(_0376_),
    .B(net270),
    .A_N(_0375_));
 sg13g2_o21ai_1 _1217_ (.B1(net115),
    .Y(_0377_),
    .A1(_0347_),
    .A2(net272));
 sg13g2_a21oi_1 _1218_ (.A1(_0376_),
    .A2(_0377_),
    .Y(_0020_),
    .B1(net316));
 sg13g2_mux2_1 _1219_ (.A0(_0129_),
    .A1(_0128_),
    .S(net366),
    .X(_0378_));
 sg13g2_nand2_1 _1220_ (.Y(_0379_),
    .A(net322),
    .B(_0364_));
 sg13g2_o21ai_1 _1221_ (.B1(_0379_),
    .Y(_0380_),
    .A1(net325),
    .A2(_0378_));
 sg13g2_and2_1 _1222_ (.A(net339),
    .B(_0380_),
    .X(_0381_));
 sg13g2_a21oi_1 _1223_ (.A1(net329),
    .A2(_0381_),
    .Y(_0382_),
    .B1(net286));
 sg13g2_a21oi_1 _1224_ (.A1(_0129_),
    .A2(net283),
    .Y(_0383_),
    .B1(_0382_));
 sg13g2_o21ai_1 _1225_ (.B1(net380),
    .Y(_0384_),
    .A1(_0347_),
    .A2(_0383_));
 sg13g2_a21oi_1 _1226_ (.A1(_0128_),
    .A2(net260),
    .Y(_0021_),
    .B1(_0384_));
 sg13g2_nor2_1 _1227_ (.A(\adc_data0[3] ),
    .B(net366),
    .Y(_0385_));
 sg13g2_a21oi_1 _1228_ (.A1(_0127_),
    .A2(net366),
    .Y(_0386_),
    .B1(_0385_));
 sg13g2_nand2_1 _1229_ (.Y(_0387_),
    .A(net350),
    .B(_0386_));
 sg13g2_o21ai_1 _1230_ (.B1(_0387_),
    .Y(_0388_),
    .A1(net350),
    .A2(_0370_));
 sg13g2_nor2_2 _1231_ (.A(net338),
    .B(net322),
    .Y(_0389_));
 sg13g2_a22oi_1 _1232_ (.Y(_0390_),
    .B1(_0389_),
    .B2(_0369_),
    .A2(_0388_),
    .A1(net340));
 sg13g2_o21ai_1 _1233_ (.B1(net290),
    .Y(_0391_),
    .A1(net326),
    .A2(_0390_));
 sg13g2_o21ai_1 _1234_ (.B1(_0391_),
    .Y(_0392_),
    .A1(net141),
    .A2(net276));
 sg13g2_a221oi_1 _1235_ (.B2(net269),
    .C1(net315),
    .B1(_0392_),
    .A1(_0127_),
    .Y(_0022_),
    .A2(net260));
 sg13g2_nor2_1 _1236_ (.A(\adc_data0[4] ),
    .B(net366),
    .Y(_0393_));
 sg13g2_a21oi_1 _1237_ (.A1(_0126_),
    .A2(net366),
    .Y(_0394_),
    .B1(_0393_));
 sg13g2_nand2_1 _1238_ (.Y(_0395_),
    .A(net350),
    .B(_0394_));
 sg13g2_o21ai_1 _1239_ (.B1(_0395_),
    .Y(_0396_),
    .A1(net351),
    .A2(_0378_));
 sg13g2_mux2_1 _1240_ (.A0(_0365_),
    .A1(_0396_),
    .S(net339),
    .X(_0397_));
 sg13g2_a21o_1 _1241_ (.A2(_0397_),
    .A1(net329),
    .B1(net286),
    .X(_0398_));
 sg13g2_o21ai_1 _1242_ (.B1(_0398_),
    .Y(_0399_),
    .A1(net171),
    .A2(net276));
 sg13g2_a221oi_1 _1243_ (.B2(net269),
    .C1(net316),
    .B1(_0399_),
    .A1(_0126_),
    .Y(_0023_),
    .A2(net260));
 sg13g2_a22oi_1 _1244_ (.Y(_0400_),
    .B1(net277),
    .B2(\adc_data0[6] ),
    .A2(net281),
    .A1(\adc_data0[5] ));
 sg13g2_or2_1 _1245_ (.X(_0401_),
    .B(_0400_),
    .A(net291));
 sg13g2_nand2b_1 _1246_ (.Y(_0402_),
    .B(net367),
    .A_N(\adc_data0[6] ));
 sg13g2_o21ai_1 _1247_ (.B1(_0402_),
    .Y(_0403_),
    .A1(\adc_data0[5] ),
    .A2(net367));
 sg13g2_nor2_1 _1248_ (.A(net351),
    .B(_0386_),
    .Y(_0404_));
 sg13g2_a21oi_1 _1249_ (.A1(net350),
    .A2(_0403_),
    .Y(_0405_),
    .B1(_0404_));
 sg13g2_mux2_1 _1250_ (.A0(_0372_),
    .A1(_0405_),
    .S(net340),
    .X(_0406_));
 sg13g2_nand3_1 _1251_ (.B(_0374_),
    .C(_0406_),
    .A(net297),
    .Y(_0407_));
 sg13g2_nand2_1 _1252_ (.Y(_0408_),
    .A(net206),
    .B(net296));
 sg13g2_nand4_1 _1253_ (.B(_0401_),
    .C(_0407_),
    .A(net270),
    .Y(_0409_),
    .D(_0408_));
 sg13g2_o21ai_1 _1254_ (.B1(net380),
    .Y(_0410_),
    .A1(net216),
    .A2(net271));
 sg13g2_nor2b_1 _1255_ (.A(_0410_),
    .B_N(_0409_),
    .Y(_0024_));
 sg13g2_nor2_1 _1256_ (.A(\adc_data0[6] ),
    .B(net366),
    .Y(_0411_));
 sg13g2_a21oi_1 _1257_ (.A1(_0125_),
    .A2(net366),
    .Y(_0412_),
    .B1(_0411_));
 sg13g2_mux2_1 _1258_ (.A0(_0394_),
    .A1(_0412_),
    .S(net350),
    .X(_0413_));
 sg13g2_mux2_1 _1259_ (.A0(_0380_),
    .A1(_0413_),
    .S(net339),
    .X(_0414_));
 sg13g2_a21o_1 _1260_ (.A2(_0414_),
    .A1(net329),
    .B1(net287),
    .X(_0415_));
 sg13g2_o21ai_1 _1261_ (.B1(_0415_),
    .Y(_0416_),
    .A1(\adc_data0[6] ),
    .A2(net276));
 sg13g2_a221oi_1 _1262_ (.B2(net270),
    .C1(net316),
    .B1(_0416_),
    .A1(_0125_),
    .Y(_0025_),
    .A2(net260));
 sg13g2_mux4_1 _1263_ (.S0(net366),
    .A0(\adc_data0[5] ),
    .A1(\adc_data0[6] ),
    .A2(\adc_data0[7] ),
    .A3(\adc_data0[8] ),
    .S1(net350),
    .X(_0417_));
 sg13g2_nor2_1 _1264_ (.A(net308),
    .B(_0417_),
    .Y(_0418_));
 sg13g2_a21o_1 _1265_ (.A2(_0149_),
    .A1(\adc_data0[0] ),
    .B1(net329),
    .X(_0419_));
 sg13g2_o21ai_1 _1266_ (.B1(_0419_),
    .Y(_0420_),
    .A1(net339),
    .A2(_0388_));
 sg13g2_o21ai_1 _1267_ (.B1(net290),
    .Y(_0421_),
    .A1(_0418_),
    .A2(_0420_));
 sg13g2_o21ai_1 _1268_ (.B1(_0421_),
    .Y(_0422_),
    .A1(\adc_data0[7] ),
    .A2(net276));
 sg13g2_a221oi_1 _1269_ (.B2(net270),
    .C1(net315),
    .B1(_0422_),
    .A1(_0124_),
    .Y(_0026_),
    .A2(net260));
 sg13g2_nor2_1 _1270_ (.A(\adc_data0[8] ),
    .B(net365),
    .Y(_0423_));
 sg13g2_a21oi_1 _1271_ (.A1(_0123_),
    .A2(net365),
    .Y(_0424_),
    .B1(_0423_));
 sg13g2_mux2_1 _1272_ (.A0(_0412_),
    .A1(_0424_),
    .S(net350),
    .X(_0425_));
 sg13g2_nor2_1 _1273_ (.A(net308),
    .B(_0425_),
    .Y(_0426_));
 sg13g2_or2_1 _1274_ (.X(_0427_),
    .B(_0396_),
    .A(net339));
 sg13g2_a22oi_1 _1275_ (.Y(_0428_),
    .B1(_0427_),
    .B2(net329),
    .A2(_0365_),
    .A1(net339));
 sg13g2_nand2b_1 _1276_ (.Y(_0429_),
    .B(net328),
    .A_N(net338));
 sg13g2_o21ai_1 _1277_ (.B1(net291),
    .Y(_0430_),
    .A1(_0426_),
    .A2(_0428_));
 sg13g2_o21ai_1 _1278_ (.B1(_0430_),
    .Y(_0431_),
    .A1(net150),
    .A2(net277));
 sg13g2_a221oi_1 _1279_ (.B2(net269),
    .C1(net315),
    .B1(_0431_),
    .A1(_0123_),
    .Y(_0027_),
    .A2(net260));
 sg13g2_o21ai_1 _1280_ (.B1(net156),
    .Y(_0432_),
    .A1(_0347_),
    .A2(net272));
 sg13g2_nor2_1 _1281_ (.A(_0123_),
    .B(net276),
    .Y(_0433_));
 sg13g2_a21oi_1 _1282_ (.A1(net340),
    .A2(_0372_),
    .Y(_0434_),
    .B1(net329));
 sg13g2_mux4_1 _1283_ (.S0(net365),
    .A0(\adc_data0[7] ),
    .A1(\adc_data0[8] ),
    .A2(\adc_data0[9] ),
    .A3(\adc_data0[10] ),
    .S1(net352),
    .X(_0435_));
 sg13g2_nor2_1 _1284_ (.A(net308),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_nor2_1 _1285_ (.A(net339),
    .B(_0405_),
    .Y(_0437_));
 sg13g2_nor4_1 _1286_ (.A(net287),
    .B(_0434_),
    .C(_0436_),
    .D(_0437_),
    .Y(_0438_));
 sg13g2_o21ai_1 _1287_ (.B1(net269),
    .Y(_0439_),
    .A1(_0433_),
    .A2(_0438_));
 sg13g2_a21oi_1 _1288_ (.A1(_0432_),
    .A2(_0439_),
    .Y(_0028_),
    .B1(net315));
 sg13g2_nor2_1 _1289_ (.A(net329),
    .B(_0381_),
    .Y(_0440_));
 sg13g2_nor2_1 _1290_ (.A(\adc_data0[10] ),
    .B(net365),
    .Y(_0441_));
 sg13g2_a21oi_1 _1291_ (.A1(_0122_),
    .A2(net365),
    .Y(_0442_),
    .B1(_0441_));
 sg13g2_mux2_1 _1292_ (.A0(_0424_),
    .A1(_0442_),
    .S(net352),
    .X(_0443_));
 sg13g2_or2_1 _1293_ (.X(_0444_),
    .B(_0443_),
    .A(net308));
 sg13g2_o21ai_1 _1294_ (.B1(_0444_),
    .Y(_0445_),
    .A1(net339),
    .A2(_0413_));
 sg13g2_o21ai_1 _1295_ (.B1(net290),
    .Y(_0446_),
    .A1(_0440_),
    .A2(_0445_));
 sg13g2_o21ai_1 _1296_ (.B1(_0446_),
    .Y(_0447_),
    .A1(net156),
    .A2(net276));
 sg13g2_a221oi_1 _1297_ (.B2(net269),
    .C1(net315),
    .B1(_0447_),
    .A1(_0122_),
    .Y(_0029_),
    .A2(net260));
 sg13g2_mux4_1 _1298_ (.S0(net365),
    .A0(\adc_data0[9] ),
    .A1(\adc_data0[10] ),
    .A2(\adc_data0[11] ),
    .A3(\adc_data0[12] ),
    .S1(net352),
    .X(_0448_));
 sg13g2_nor2_1 _1299_ (.A(net308),
    .B(_0448_),
    .Y(_0449_));
 sg13g2_a21oi_1 _1300_ (.A1(net326),
    .A2(_0390_),
    .Y(_0450_),
    .B1(_0449_));
 sg13g2_o21ai_1 _1301_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_0417_),
    .A2(net304));
 sg13g2_nand2_1 _1302_ (.Y(_0452_),
    .A(net290),
    .B(_0451_));
 sg13g2_o21ai_1 _1303_ (.B1(_0452_),
    .Y(_0453_),
    .A1(net185),
    .A2(net276));
 sg13g2_a221oi_1 _1304_ (.B2(net269),
    .C1(net315),
    .B1(_0453_),
    .A1(_0121_),
    .Y(_0030_),
    .A2(net260));
 sg13g2_o21ai_1 _1305_ (.B1(net134),
    .Y(_0454_),
    .A1(_0347_),
    .A2(net272));
 sg13g2_or2_1 _1306_ (.X(_0455_),
    .B(net304),
    .A(_0425_));
 sg13g2_nand2_1 _1307_ (.Y(_0456_),
    .A(net325),
    .B(_0442_));
 sg13g2_nand2_1 _1308_ (.Y(_0457_),
    .A(\adc_data0[13] ),
    .B(net365));
 sg13g2_o21ai_1 _1309_ (.B1(_0457_),
    .Y(_0458_),
    .A1(_0121_),
    .A2(net365));
 sg13g2_a21oi_1 _1310_ (.A1(net352),
    .A2(_0458_),
    .Y(_0459_),
    .B1(net308));
 sg13g2_o21ai_1 _1311_ (.B1(_0455_),
    .Y(_0460_),
    .A1(net330),
    .A2(_0397_));
 sg13g2_a21oi_1 _1312_ (.A1(_0456_),
    .A2(_0459_),
    .Y(_0461_),
    .B1(_0460_));
 sg13g2_a22oi_1 _1313_ (.Y(_0462_),
    .B1(_0461_),
    .B2(net290),
    .A2(net283),
    .A1(\adc_data0[12] ));
 sg13g2_nand2b_1 _1314_ (.Y(_0463_),
    .B(net269),
    .A_N(_0462_));
 sg13g2_a21oi_1 _1315_ (.A1(_0454_),
    .A2(_0463_),
    .Y(_0031_),
    .B1(net315));
 sg13g2_nor2_1 _1316_ (.A(net330),
    .B(_0406_),
    .Y(_0464_));
 sg13g2_mux4_1 _1317_ (.S0(net368),
    .A0(\adc_data0[11] ),
    .A1(\adc_data0[12] ),
    .A2(\adc_data0[13] ),
    .A3(\adc_data0[14] ),
    .S1(net352),
    .X(_0465_));
 sg13g2_or2_1 _1318_ (.X(_0466_),
    .B(_0465_),
    .A(net308));
 sg13g2_o21ai_1 _1319_ (.B1(_0466_),
    .Y(_0467_),
    .A1(net306),
    .A2(_0435_));
 sg13g2_o21ai_1 _1320_ (.B1(net290),
    .Y(_0468_),
    .A1(_0464_),
    .A2(_0467_));
 sg13g2_o21ai_1 _1321_ (.B1(_0468_),
    .Y(_0469_),
    .A1(net134),
    .A2(net276));
 sg13g2_a221oi_1 _1322_ (.B2(net271),
    .C1(net315),
    .B1(_0469_),
    .A1(_0120_),
    .Y(_0032_),
    .A2(_0362_));
 sg13g2_a21oi_1 _1323_ (.A1(net271),
    .A2(net281),
    .Y(_0470_),
    .B1(net121));
 sg13g2_mux2_1 _1324_ (.A0(_0237_),
    .A1(_0247_),
    .S(_0345_),
    .X(_0471_));
 sg13g2_mux2_1 _1325_ (.A0(_0238_),
    .A1(_0248_),
    .S(_0345_),
    .X(_0472_));
 sg13g2_a21oi_1 _1326_ (.A1(_0144_),
    .A2(net281),
    .Y(_0473_),
    .B1(_0355_));
 sg13g2_o21ai_1 _1327_ (.B1(net379),
    .Y(_0474_),
    .A1(_0472_),
    .A2(_0473_));
 sg13g2_nor2_1 _1328_ (.A(net122),
    .B(_0474_),
    .Y(_0033_));
 sg13g2_nand2_2 _1329_ (.Y(_0475_),
    .A(_0361_),
    .B(net268));
 sg13g2_nor2_1 _1330_ (.A(\adc_data1[0] ),
    .B(net371),
    .Y(_0476_));
 sg13g2_a21oi_1 _1331_ (.A1(_0119_),
    .A2(net371),
    .Y(_0477_),
    .B1(_0476_));
 sg13g2_and2_1 _1332_ (.A(net355),
    .B(_0477_),
    .X(_0478_));
 sg13g2_nand3_1 _1333_ (.B(net343),
    .C(_0478_),
    .A(net332),
    .Y(_0479_));
 sg13g2_nand2_1 _1334_ (.Y(_0480_),
    .A(net292),
    .B(_0479_));
 sg13g2_o21ai_1 _1335_ (.B1(_0480_),
    .Y(_0481_),
    .A1(net121),
    .A2(net278));
 sg13g2_a221oi_1 _1336_ (.B2(net267),
    .C1(net319),
    .B1(_0481_),
    .A1(_0119_),
    .Y(_0034_),
    .A2(net259));
 sg13g2_and2_1 _1337_ (.A(\adc_data1[0] ),
    .B(net371),
    .X(_0482_));
 sg13g2_mux2_1 _1338_ (.A0(_0119_),
    .A1(_0118_),
    .S(net371),
    .X(_0483_));
 sg13g2_nor2_1 _1339_ (.A(net357),
    .B(_0482_),
    .Y(_0484_));
 sg13g2_a21oi_1 _1340_ (.A1(net357),
    .A2(_0483_),
    .Y(_0485_),
    .B1(_0484_));
 sg13g2_nand3_1 _1341_ (.B(net342),
    .C(_0485_),
    .A(net332),
    .Y(_0486_));
 sg13g2_a22oi_1 _1342_ (.Y(_0487_),
    .B1(_0486_),
    .B2(net293),
    .A2(net284),
    .A1(_0119_));
 sg13g2_o21ai_1 _1343_ (.B1(net380),
    .Y(_0488_),
    .A1(_0472_),
    .A2(_0487_));
 sg13g2_a21oi_1 _1344_ (.A1(_0118_),
    .A2(net259),
    .Y(_0035_),
    .B1(_0488_));
 sg13g2_nand2b_1 _1345_ (.Y(_0489_),
    .B(net363),
    .A_N(\adc_data1[3] ));
 sg13g2_o21ai_1 _1346_ (.B1(_0489_),
    .Y(_0490_),
    .A1(\adc_data1[2] ),
    .A2(net363));
 sg13g2_nand2_1 _1347_ (.Y(_0491_),
    .A(net323),
    .B(_0477_));
 sg13g2_o21ai_1 _1348_ (.B1(_0491_),
    .Y(_0492_),
    .A1(net323),
    .A2(_0490_));
 sg13g2_and2_1 _1349_ (.A(net342),
    .B(_0492_),
    .X(_0493_));
 sg13g2_a22oi_1 _1350_ (.Y(_0494_),
    .B1(_0374_),
    .B2(_0493_),
    .A2(net282),
    .A1(net138));
 sg13g2_nand2b_1 _1351_ (.Y(_0495_),
    .B(net267),
    .A_N(_0494_));
 sg13g2_o21ai_1 _1352_ (.B1(net168),
    .Y(_0496_),
    .A1(net272),
    .A2(_0472_));
 sg13g2_a21oi_1 _1353_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0036_),
    .B1(net313));
 sg13g2_nor2_1 _1354_ (.A(\adc_data1[3] ),
    .B(net363),
    .Y(_0497_));
 sg13g2_a21oi_1 _1355_ (.A1(_0117_),
    .A2(net364),
    .Y(_0498_),
    .B1(_0497_));
 sg13g2_nand2_1 _1356_ (.Y(_0499_),
    .A(net349),
    .B(_0498_));
 sg13g2_o21ai_1 _1357_ (.B1(_0499_),
    .Y(_0500_),
    .A1(net355),
    .A2(_0483_));
 sg13g2_a22oi_1 _1358_ (.Y(_0501_),
    .B1(_0500_),
    .B2(net342),
    .A2(_0482_),
    .A1(_0389_));
 sg13g2_o21ai_1 _1359_ (.B1(net289),
    .Y(_0502_),
    .A1(net326),
    .A2(_0501_));
 sg13g2_o21ai_1 _1360_ (.B1(_0502_),
    .Y(_0503_),
    .A1(\adc_data1[3] ),
    .A2(net278));
 sg13g2_a221oi_1 _1361_ (.B2(net267),
    .C1(net313),
    .B1(_0503_),
    .A1(_0117_),
    .Y(_0037_),
    .A2(net259));
 sg13g2_nor2_1 _1362_ (.A(\adc_data1[4] ),
    .B(net363),
    .Y(_0504_));
 sg13g2_a21oi_1 _1363_ (.A1(_0116_),
    .A2(net364),
    .Y(_0505_),
    .B1(_0504_));
 sg13g2_nand2_1 _1364_ (.Y(_0506_),
    .A(net349),
    .B(_0505_));
 sg13g2_o21ai_1 _1365_ (.B1(_0506_),
    .Y(_0507_),
    .A1(net349),
    .A2(_0490_));
 sg13g2_mux2_1 _1366_ (.A0(_0478_),
    .A1(_0507_),
    .S(net342),
    .X(_0508_));
 sg13g2_a21o_1 _1367_ (.A2(_0508_),
    .A1(net332),
    .B1(net287),
    .X(_0509_));
 sg13g2_o21ai_1 _1368_ (.B1(_0509_),
    .Y(_0510_),
    .A1(net166),
    .A2(net275));
 sg13g2_a221oi_1 _1369_ (.B2(net267),
    .C1(net313),
    .B1(_0510_),
    .A1(_0116_),
    .Y(_0038_),
    .A2(net259));
 sg13g2_nand2_1 _1370_ (.Y(_0511_),
    .A(_0115_),
    .B(net363));
 sg13g2_o21ai_1 _1371_ (.B1(_0511_),
    .Y(_0512_),
    .A1(\adc_data1[5] ),
    .A2(net370));
 sg13g2_nor2_1 _1372_ (.A(net349),
    .B(_0498_),
    .Y(_0513_));
 sg13g2_a21oi_1 _1373_ (.A1(net349),
    .A2(_0512_),
    .Y(_0514_),
    .B1(_0513_));
 sg13g2_mux2_1 _1374_ (.A0(_0485_),
    .A1(_0514_),
    .S(net342),
    .X(_0515_));
 sg13g2_a21o_1 _1375_ (.A2(_0515_),
    .A1(net332),
    .B1(net287),
    .X(_0516_));
 sg13g2_o21ai_1 _1376_ (.B1(_0516_),
    .Y(_0517_),
    .A1(net193),
    .A2(net278));
 sg13g2_a221oi_1 _1377_ (.B2(net267),
    .C1(net314),
    .B1(_0517_),
    .A1(_0115_),
    .Y(_0039_),
    .A2(net259));
 sg13g2_nor2_1 _1378_ (.A(\adc_data1[6] ),
    .B(net370),
    .Y(_0518_));
 sg13g2_a21oi_1 _1379_ (.A1(_0114_),
    .A2(net370),
    .Y(_0519_),
    .B1(_0518_));
 sg13g2_mux2_1 _1380_ (.A0(_0505_),
    .A1(_0519_),
    .S(net354),
    .X(_0520_));
 sg13g2_mux2_1 _1381_ (.A0(_0492_),
    .A1(_0520_),
    .S(net342),
    .X(_0521_));
 sg13g2_a21o_1 _1382_ (.A2(_0521_),
    .A1(net332),
    .B1(_0275_),
    .X(_0522_));
 sg13g2_o21ai_1 _1383_ (.B1(_0522_),
    .Y(_0523_),
    .A1(\adc_data1[6] ),
    .A2(net278));
 sg13g2_a221oi_1 _1384_ (.B2(net267),
    .C1(net318),
    .B1(_0523_),
    .A1(_0114_),
    .Y(_0040_),
    .A2(net259));
 sg13g2_nor2_1 _1385_ (.A(net343),
    .B(_0500_),
    .Y(_0524_));
 sg13g2_mux4_1 _1386_ (.S0(net370),
    .A0(\adc_data1[5] ),
    .A1(\adc_data1[6] ),
    .A2(\adc_data1[7] ),
    .A3(\adc_data1[8] ),
    .S1(net355),
    .X(_0525_));
 sg13g2_nor2_1 _1387_ (.A(net310),
    .B(_0525_),
    .Y(_0526_));
 sg13g2_a21oi_1 _1388_ (.A1(net121),
    .A2(_0149_),
    .Y(_0527_),
    .B1(net333));
 sg13g2_nor3_1 _1389_ (.A(_0524_),
    .B(_0526_),
    .C(_0527_),
    .Y(_0528_));
 sg13g2_a22oi_1 _1390_ (.Y(_0529_),
    .B1(_0528_),
    .B2(net292),
    .A2(net284),
    .A1(\adc_data1[7] ));
 sg13g2_nand2b_1 _1391_ (.Y(_0530_),
    .B(net267),
    .A_N(_0529_));
 sg13g2_o21ai_1 _1392_ (.B1(net162),
    .Y(_0531_),
    .A1(net273),
    .A2(_0472_));
 sg13g2_a21oi_1 _1393_ (.A1(_0530_),
    .A2(_0531_),
    .Y(_0041_),
    .B1(net318));
 sg13g2_nor2_1 _1394_ (.A(\adc_data1[8] ),
    .B(net370),
    .Y(_0532_));
 sg13g2_a21oi_1 _1395_ (.A1(_0113_),
    .A2(net371),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_mux2_1 _1396_ (.A0(_0519_),
    .A1(_0533_),
    .S(net355),
    .X(_0534_));
 sg13g2_or2_1 _1397_ (.X(_0535_),
    .B(_0534_),
    .A(net310));
 sg13g2_a21oi_1 _1398_ (.A1(net342),
    .A2(_0478_),
    .Y(_0536_),
    .B1(net332));
 sg13g2_o21ai_1 _1399_ (.B1(_0535_),
    .Y(_0537_),
    .A1(net305),
    .A2(_0507_));
 sg13g2_o21ai_1 _1400_ (.B1(net292),
    .Y(_0538_),
    .A1(_0536_),
    .A2(_0537_));
 sg13g2_o21ai_1 _1401_ (.B1(_0538_),
    .Y(_0539_),
    .A1(net162),
    .A2(net278));
 sg13g2_a221oi_1 _1402_ (.B2(net268),
    .C1(net318),
    .B1(_0539_),
    .A1(_0113_),
    .Y(_0042_),
    .A2(net259));
 sg13g2_a21oi_1 _1403_ (.A1(net343),
    .A2(_0485_),
    .Y(_0540_),
    .B1(net333));
 sg13g2_mux4_1 _1404_ (.S0(net370),
    .A0(\adc_data1[7] ),
    .A1(\adc_data1[8] ),
    .A2(\adc_data1[9] ),
    .A3(\adc_data1[10] ),
    .S1(net355),
    .X(_0541_));
 sg13g2_or2_1 _1405_ (.X(_0542_),
    .B(_0541_),
    .A(net310));
 sg13g2_o21ai_1 _1406_ (.B1(_0542_),
    .Y(_0543_),
    .A1(net343),
    .A2(_0514_));
 sg13g2_o21ai_1 _1407_ (.B1(net292),
    .Y(_0544_),
    .A1(_0540_),
    .A2(_0543_));
 sg13g2_o21ai_1 _1408_ (.B1(_0544_),
    .Y(_0545_),
    .A1(\adc_data1[9] ),
    .A2(net278));
 sg13g2_a221oi_1 _1409_ (.B2(net268),
    .C1(net318),
    .B1(_0545_),
    .A1(_0112_),
    .Y(_0043_),
    .A2(_0475_));
 sg13g2_nor2_1 _1410_ (.A(net332),
    .B(_0493_),
    .Y(_0546_));
 sg13g2_or2_1 _1411_ (.X(_0547_),
    .B(_0520_),
    .A(net342));
 sg13g2_mux2_1 _1412_ (.A0(_0112_),
    .A1(_0111_),
    .S(net370),
    .X(_0548_));
 sg13g2_nand2_1 _1413_ (.Y(_0549_),
    .A(net323),
    .B(_0533_));
 sg13g2_o21ai_1 _1414_ (.B1(_0549_),
    .Y(_0550_),
    .A1(net323),
    .A2(_0548_));
 sg13g2_o21ai_1 _1415_ (.B1(_0547_),
    .Y(_0551_),
    .A1(net310),
    .A2(_0550_));
 sg13g2_o21ai_1 _1416_ (.B1(net292),
    .Y(_0552_),
    .A1(_0546_),
    .A2(_0551_));
 sg13g2_o21ai_1 _1417_ (.B1(_0552_),
    .Y(_0553_),
    .A1(net183),
    .A2(net279));
 sg13g2_a221oi_1 _1418_ (.B2(net268),
    .C1(net318),
    .B1(_0553_),
    .A1(_0111_),
    .Y(_0044_),
    .A2(_0475_));
 sg13g2_o21ai_1 _1419_ (.B1(net147),
    .Y(_0554_),
    .A1(net273),
    .A2(_0472_));
 sg13g2_nor2_1 _1420_ (.A(_0111_),
    .B(net279),
    .Y(_0555_));
 sg13g2_nor2_1 _1421_ (.A(net305),
    .B(_0525_),
    .Y(_0556_));
 sg13g2_mux4_1 _1422_ (.S0(net370),
    .A0(\adc_data1[9] ),
    .A1(\adc_data1[10] ),
    .A2(\adc_data1[11] ),
    .A3(\adc_data1[12] ),
    .S1(net355),
    .X(_0557_));
 sg13g2_a21oi_1 _1423_ (.A1(net326),
    .A2(_0501_),
    .Y(_0558_),
    .B1(_0556_));
 sg13g2_o21ai_1 _1424_ (.B1(_0558_),
    .Y(_0559_),
    .A1(net309),
    .A2(_0557_));
 sg13g2_nor2_1 _1425_ (.A(net287),
    .B(_0559_),
    .Y(_0560_));
 sg13g2_o21ai_1 _1426_ (.B1(net268),
    .Y(_0561_),
    .A1(_0555_),
    .A2(_0560_));
 sg13g2_a21oi_1 _1427_ (.A1(_0554_),
    .A2(_0561_),
    .Y(_0045_),
    .B1(net320));
 sg13g2_nor2_1 _1428_ (.A(net305),
    .B(_0534_),
    .Y(_0562_));
 sg13g2_nor2_1 _1429_ (.A(\adc_data1[12] ),
    .B(net374),
    .Y(_0563_));
 sg13g2_a21oi_1 _1430_ (.A1(_0110_),
    .A2(net374),
    .Y(_0564_),
    .B1(_0563_));
 sg13g2_a21oi_1 _1431_ (.A1(net355),
    .A2(_0564_),
    .Y(_0565_),
    .B1(net310));
 sg13g2_o21ai_1 _1432_ (.B1(_0565_),
    .Y(_0566_),
    .A1(net355),
    .A2(_0548_));
 sg13g2_o21ai_1 _1433_ (.B1(_0566_),
    .Y(_0567_),
    .A1(net333),
    .A2(_0508_));
 sg13g2_o21ai_1 _1434_ (.B1(net292),
    .Y(_0568_),
    .A1(_0562_),
    .A2(_0567_));
 sg13g2_o21ai_1 _1435_ (.B1(_0568_),
    .Y(_0569_),
    .A1(net147),
    .A2(net278));
 sg13g2_a221oi_1 _1436_ (.B2(net268),
    .C1(net320),
    .B1(_0569_),
    .A1(_0110_),
    .Y(_0046_),
    .A2(_0475_));
 sg13g2_nor2_1 _1437_ (.A(net333),
    .B(_0515_),
    .Y(_0570_));
 sg13g2_mux4_1 _1438_ (.S0(net374),
    .A0(\adc_data1[11] ),
    .A1(\adc_data1[12] ),
    .A2(\adc_data1[13] ),
    .A3(\adc_data1[14] ),
    .S1(net356),
    .X(_0571_));
 sg13g2_or2_1 _1439_ (.X(_0572_),
    .B(_0571_),
    .A(net309));
 sg13g2_o21ai_1 _1440_ (.B1(_0572_),
    .Y(_0573_),
    .A1(net306),
    .A2(_0541_));
 sg13g2_o21ai_1 _1441_ (.B1(net292),
    .Y(_0574_),
    .A1(_0570_),
    .A2(_0573_));
 sg13g2_o21ai_1 _1442_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net170),
    .A2(net279));
 sg13g2_a221oi_1 _1443_ (.B2(net268),
    .C1(net318),
    .B1(_0575_),
    .A1(_0109_),
    .Y(_0047_),
    .A2(net259));
 sg13g2_a21oi_1 _1444_ (.A1(net271),
    .A2(net281),
    .Y(_0576_),
    .B1(net113));
 sg13g2_and2_1 _1445_ (.A(_0218_),
    .B(_0227_),
    .X(_0577_));
 sg13g2_nor4_1 _1446_ (.A(tx_cs_n),
    .B(_0338_),
    .C(_0344_),
    .D(_0577_),
    .Y(_0578_));
 sg13g2_a21oi_2 _1447_ (.B1(_0578_),
    .Y(_0579_),
    .A2(_0345_),
    .A1(_0248_));
 sg13g2_a21o_1 _1448_ (.A2(_0345_),
    .A1(_0248_),
    .B1(_0578_),
    .X(_0580_));
 sg13g2_a21oi_1 _1449_ (.A1(_0143_),
    .A2(net281),
    .Y(_0581_),
    .B1(_0355_));
 sg13g2_o21ai_1 _1450_ (.B1(net379),
    .Y(_0582_),
    .A1(net264),
    .A2(_0581_));
 sg13g2_nor2_1 _1451_ (.A(net114),
    .B(_0582_),
    .Y(_0048_));
 sg13g2_nand2_2 _1452_ (.Y(_0583_),
    .A(_0361_),
    .B(net265));
 sg13g2_nand2_1 _1453_ (.Y(_0584_),
    .A(\adc_data2[1] ),
    .B(net376));
 sg13g2_o21ai_1 _1454_ (.B1(_0584_),
    .Y(_0585_),
    .A1(_0108_),
    .A2(net376));
 sg13g2_and2_1 _1455_ (.A(net358),
    .B(_0585_),
    .X(_0586_));
 sg13g2_nand3_1 _1456_ (.B(net346),
    .C(_0586_),
    .A(net335),
    .Y(_0587_));
 sg13g2_a22oi_1 _1457_ (.Y(_0588_),
    .B1(_0587_),
    .B2(net294),
    .A2(net285),
    .A1(_0108_));
 sg13g2_o21ai_1 _1458_ (.B1(net379),
    .Y(_0589_),
    .A1(net264),
    .A2(_0588_));
 sg13g2_a21oi_1 _1459_ (.A1(_0107_),
    .A2(_0583_),
    .Y(_0049_),
    .B1(_0589_));
 sg13g2_and2_1 _1460_ (.A(\adc_data2[0] ),
    .B(net376),
    .X(_0590_));
 sg13g2_mux2_1 _1461_ (.A0(_0107_),
    .A1(_0106_),
    .S(net376),
    .X(_0591_));
 sg13g2_nor2_1 _1462_ (.A(net358),
    .B(_0590_),
    .Y(_0592_));
 sg13g2_a21oi_1 _1463_ (.A1(net358),
    .A2(_0591_),
    .Y(_0593_),
    .B1(_0592_));
 sg13g2_nand3_1 _1464_ (.B(net346),
    .C(_0593_),
    .A(net335),
    .Y(_0594_));
 sg13g2_a22oi_1 _1465_ (.Y(_0595_),
    .B1(_0594_),
    .B2(net294),
    .A2(net285),
    .A1(_0107_));
 sg13g2_o21ai_1 _1466_ (.B1(net379),
    .Y(_0596_),
    .A1(net264),
    .A2(_0595_));
 sg13g2_a21oi_1 _1467_ (.A1(_0106_),
    .A2(_0583_),
    .Y(_0050_),
    .B1(_0596_));
 sg13g2_mux2_1 _1468_ (.A0(_0106_),
    .A1(_0105_),
    .S(net376),
    .X(_0597_));
 sg13g2_nand2_1 _1469_ (.Y(_0598_),
    .A(net324),
    .B(_0585_));
 sg13g2_o21ai_1 _1470_ (.B1(_0598_),
    .Y(_0599_),
    .A1(net324),
    .A2(_0597_));
 sg13g2_and2_1 _1471_ (.A(net344),
    .B(_0599_),
    .X(_0600_));
 sg13g2_nand2_1 _1472_ (.Y(_0601_),
    .A(net336),
    .B(_0600_));
 sg13g2_a22oi_1 _1473_ (.Y(_0602_),
    .B1(_0601_),
    .B2(net294),
    .A2(net285),
    .A1(_0106_));
 sg13g2_o21ai_1 _1474_ (.B1(net379),
    .Y(_0603_),
    .A1(net263),
    .A2(_0602_));
 sg13g2_a21oi_1 _1475_ (.A1(_0105_),
    .A2(_0583_),
    .Y(_0051_),
    .B1(_0603_));
 sg13g2_o21ai_1 _1476_ (.B1(net139),
    .Y(_0604_),
    .A1(net273),
    .A2(net264));
 sg13g2_nand2_1 _1477_ (.Y(_0605_),
    .A(\adc_data2[4] ),
    .B(net376));
 sg13g2_o21ai_1 _1478_ (.B1(_0605_),
    .Y(_0606_),
    .A1(_0105_),
    .A2(net376));
 sg13g2_nand2_1 _1479_ (.Y(_0607_),
    .A(net358),
    .B(_0606_));
 sg13g2_o21ai_1 _1480_ (.B1(_0607_),
    .Y(_0608_),
    .A1(net358),
    .A2(_0591_));
 sg13g2_a22oi_1 _1481_ (.Y(_0609_),
    .B1(_0608_),
    .B2(net344),
    .A2(_0590_),
    .A1(_0389_));
 sg13g2_inv_1 _1482_ (.Y(_0610_),
    .A(_0609_));
 sg13g2_a22oi_1 _1483_ (.Y(_0611_),
    .B1(_0374_),
    .B2(_0610_),
    .A2(net285),
    .A1(\adc_data2[3] ));
 sg13g2_nand2b_1 _1484_ (.Y(_0612_),
    .B(net265),
    .A_N(_0611_));
 sg13g2_a21oi_1 _1485_ (.A1(_0604_),
    .A2(_0612_),
    .Y(_0052_),
    .B1(net321));
 sg13g2_o21ai_1 _1486_ (.B1(net145),
    .Y(_0613_),
    .A1(net273),
    .A2(net263));
 sg13g2_mux2_1 _1487_ (.A0(\adc_data2[4] ),
    .A1(\adc_data2[5] ),
    .S(net376),
    .X(_0614_));
 sg13g2_nand2_1 _1488_ (.Y(_0615_),
    .A(net358),
    .B(_0614_));
 sg13g2_o21ai_1 _1489_ (.B1(_0615_),
    .Y(_0616_),
    .A1(net358),
    .A2(_0597_));
 sg13g2_mux2_1 _1490_ (.A0(_0586_),
    .A1(_0616_),
    .S(net344),
    .X(_0617_));
 sg13g2_a22oi_1 _1491_ (.Y(_0618_),
    .B1(_0374_),
    .B2(_0617_),
    .A2(net285),
    .A1(net139));
 sg13g2_nand2b_1 _1492_ (.Y(_0619_),
    .B(net265),
    .A_N(_0618_));
 sg13g2_a21oi_1 _1493_ (.A1(_0613_),
    .A2(_0619_),
    .Y(_0053_),
    .B1(net321));
 sg13g2_o21ai_1 _1494_ (.B1(net143),
    .Y(_0620_),
    .A1(net273),
    .A2(net263));
 sg13g2_nor2b_1 _1495_ (.A(net372),
    .B_N(\adc_data2[5] ),
    .Y(_0621_));
 sg13g2_a21oi_1 _1496_ (.A1(\adc_data2[6] ),
    .A2(net372),
    .Y(_0622_),
    .B1(_0621_));
 sg13g2_nor2_1 _1497_ (.A(net358),
    .B(_0606_),
    .Y(_0623_));
 sg13g2_a21oi_1 _1498_ (.A1(net359),
    .A2(_0622_),
    .Y(_0624_),
    .B1(_0623_));
 sg13g2_mux2_1 _1499_ (.A0(_0593_),
    .A1(_0624_),
    .S(net344),
    .X(_0625_));
 sg13g2_a22oi_1 _1500_ (.Y(_0626_),
    .B1(_0374_),
    .B2(_0625_),
    .A2(net284),
    .A1(\adc_data2[5] ));
 sg13g2_nand2b_1 _1501_ (.Y(_0627_),
    .B(net265),
    .A_N(_0626_));
 sg13g2_a21oi_1 _1502_ (.A1(_0620_),
    .A2(_0627_),
    .Y(_0054_),
    .B1(net319));
 sg13g2_o21ai_1 _1503_ (.B1(net132),
    .Y(_0628_),
    .A1(net273),
    .A2(net263));
 sg13g2_nor2_1 _1504_ (.A(\adc_data2[6] ),
    .B(net373),
    .Y(_0629_));
 sg13g2_a21oi_1 _1505_ (.A1(_0104_),
    .A2(net372),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_mux2_1 _1506_ (.A0(_0614_),
    .A1(_0630_),
    .S(net356),
    .X(_0631_));
 sg13g2_mux2_1 _1507_ (.A0(_0599_),
    .A1(_0631_),
    .S(net344),
    .X(_0632_));
 sg13g2_a22oi_1 _1508_ (.Y(_0633_),
    .B1(_0374_),
    .B2(_0632_),
    .A2(net284),
    .A1(\adc_data2[6] ));
 sg13g2_nand2b_1 _1509_ (.Y(_0634_),
    .B(net265),
    .A_N(_0633_));
 sg13g2_a21oi_1 _1510_ (.A1(_0628_),
    .A2(_0634_),
    .Y(_0055_),
    .B1(net319));
 sg13g2_mux4_1 _1511_ (.S0(net373),
    .A0(\adc_data2[5] ),
    .A1(\adc_data2[6] ),
    .A2(\adc_data2[7] ),
    .A3(\adc_data2[8] ),
    .S1(net356),
    .X(_0635_));
 sg13g2_nor2_1 _1512_ (.A(net309),
    .B(_0635_),
    .Y(_0636_));
 sg13g2_a21oi_1 _1513_ (.A1(\adc_data2[0] ),
    .A2(_0149_),
    .Y(_0637_),
    .B1(net334));
 sg13g2_nor2_1 _1514_ (.A(_0636_),
    .B(_0637_),
    .Y(_0638_));
 sg13g2_o21ai_1 _1515_ (.B1(_0638_),
    .Y(_0639_),
    .A1(net344),
    .A2(_0608_));
 sg13g2_a22oi_1 _1516_ (.Y(_0640_),
    .B1(_0639_),
    .B2(net294),
    .A2(net284),
    .A1(_0104_));
 sg13g2_o21ai_1 _1517_ (.B1(net379),
    .Y(_0641_),
    .A1(net263),
    .A2(_0640_));
 sg13g2_a21oi_1 _1518_ (.A1(_0103_),
    .A2(_0583_),
    .Y(_0056_),
    .B1(_0641_));
 sg13g2_nor2_1 _1519_ (.A(\adc_data2[8] ),
    .B(net372),
    .Y(_0642_));
 sg13g2_a21oi_1 _1520_ (.A1(_0102_),
    .A2(net372),
    .Y(_0643_),
    .B1(_0642_));
 sg13g2_mux2_1 _1521_ (.A0(_0630_),
    .A1(_0643_),
    .S(net356),
    .X(_0644_));
 sg13g2_nor2_1 _1522_ (.A(net309),
    .B(_0644_),
    .Y(_0645_));
 sg13g2_a21oi_1 _1523_ (.A1(net344),
    .A2(_0586_),
    .Y(_0646_),
    .B1(net336));
 sg13g2_nor2_1 _1524_ (.A(_0645_),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_o21ai_1 _1525_ (.B1(_0647_),
    .Y(_0648_),
    .A1(net344),
    .A2(_0616_));
 sg13g2_a22oi_1 _1526_ (.Y(_0649_),
    .B1(_0648_),
    .B2(net294),
    .A2(net285),
    .A1(_0103_));
 sg13g2_o21ai_1 _1527_ (.B1(net1),
    .Y(_0650_),
    .A1(net263),
    .A2(_0649_));
 sg13g2_a21oi_1 _1528_ (.A1(_0102_),
    .A2(_0583_),
    .Y(_0057_),
    .B1(_0650_));
 sg13g2_a21oi_1 _1529_ (.A1(net345),
    .A2(_0593_),
    .Y(_0651_),
    .B1(net334));
 sg13g2_mux4_1 _1530_ (.S0(net372),
    .A0(\adc_data2[7] ),
    .A1(\adc_data2[8] ),
    .A2(\adc_data2[9] ),
    .A3(\adc_data2[10] ),
    .S1(net356),
    .X(_0652_));
 sg13g2_or2_1 _1531_ (.X(_0653_),
    .B(_0652_),
    .A(net309));
 sg13g2_o21ai_1 _1532_ (.B1(_0653_),
    .Y(_0654_),
    .A1(net345),
    .A2(_0624_));
 sg13g2_o21ai_1 _1533_ (.B1(net293),
    .Y(_0655_),
    .A1(_0651_),
    .A2(_0654_));
 sg13g2_o21ai_1 _1534_ (.B1(_0655_),
    .Y(_0656_),
    .A1(net146),
    .A2(net278));
 sg13g2_a221oi_1 _1535_ (.B2(net266),
    .C1(net319),
    .B1(_0656_),
    .A1(_0101_),
    .Y(_0058_),
    .A2(_0583_));
 sg13g2_o21ai_1 _1536_ (.B1(net160),
    .Y(_0657_),
    .A1(net273),
    .A2(net263));
 sg13g2_nor2_1 _1537_ (.A(net334),
    .B(_0600_),
    .Y(_0658_));
 sg13g2_nor2_1 _1538_ (.A(_0101_),
    .B(net372),
    .Y(_0659_));
 sg13g2_a21oi_1 _1539_ (.A1(\adc_data2[11] ),
    .A2(net372),
    .Y(_0660_),
    .B1(_0659_));
 sg13g2_nand2_1 _1540_ (.Y(_0661_),
    .A(net323),
    .B(_0643_));
 sg13g2_o21ai_1 _1541_ (.B1(_0661_),
    .Y(_0662_),
    .A1(net323),
    .A2(_0660_));
 sg13g2_nor2_1 _1542_ (.A(net309),
    .B(_0662_),
    .Y(_0663_));
 sg13g2_nor2_1 _1543_ (.A(net345),
    .B(_0631_),
    .Y(_0664_));
 sg13g2_nor3_1 _1544_ (.A(_0658_),
    .B(_0663_),
    .C(_0664_),
    .Y(_0665_));
 sg13g2_a22oi_1 _1545_ (.Y(_0666_),
    .B1(_0665_),
    .B2(net293),
    .A2(net284),
    .A1(\adc_data2[10] ));
 sg13g2_nand2b_1 _1546_ (.Y(_0667_),
    .B(net266),
    .A_N(_0666_));
 sg13g2_a21oi_1 _1547_ (.A1(_0657_),
    .A2(_0667_),
    .Y(_0059_),
    .B1(net319));
 sg13g2_o21ai_1 _1548_ (.B1(net169),
    .Y(_0668_),
    .A1(net273),
    .A2(net263));
 sg13g2_mux4_1 _1549_ (.S0(net374),
    .A0(\adc_data2[9] ),
    .A1(\adc_data2[10] ),
    .A2(\adc_data2[11] ),
    .A3(\adc_data2[12] ),
    .S1(net356),
    .X(_0669_));
 sg13g2_or2_1 _1550_ (.X(_0670_),
    .B(_0669_),
    .A(net309));
 sg13g2_o21ai_1 _1551_ (.B1(_0670_),
    .Y(_0671_),
    .A1(net305),
    .A2(_0635_));
 sg13g2_a21oi_1 _1552_ (.A1(_0140_),
    .A2(_0609_),
    .Y(_0672_),
    .B1(_0671_));
 sg13g2_a22oi_1 _1553_ (.Y(_0673_),
    .B1(_0672_),
    .B2(net293),
    .A2(net284),
    .A1(net160));
 sg13g2_nand2b_1 _1554_ (.Y(_0674_),
    .B(net266),
    .A_N(_0673_));
 sg13g2_a21oi_1 _1555_ (.A1(_0668_),
    .A2(_0674_),
    .Y(_0060_),
    .B1(net319));
 sg13g2_nor2_1 _1556_ (.A(net334),
    .B(_0617_),
    .Y(_0675_));
 sg13g2_nor2_1 _1557_ (.A(\adc_data2[12] ),
    .B(net373),
    .Y(_0676_));
 sg13g2_a21oi_1 _1558_ (.A1(_0100_),
    .A2(net373),
    .Y(_0677_),
    .B1(_0676_));
 sg13g2_a21oi_1 _1559_ (.A1(net356),
    .A2(_0677_),
    .Y(_0678_),
    .B1(net309));
 sg13g2_o21ai_1 _1560_ (.B1(_0678_),
    .Y(_0679_),
    .A1(net357),
    .A2(_0660_));
 sg13g2_o21ai_1 _1561_ (.B1(_0679_),
    .Y(_0680_),
    .A1(net305),
    .A2(_0644_));
 sg13g2_o21ai_1 _1562_ (.B1(net293),
    .Y(_0681_),
    .A1(_0675_),
    .A2(_0680_));
 sg13g2_o21ai_1 _1563_ (.B1(_0681_),
    .Y(_0682_),
    .A1(net169),
    .A2(net279));
 sg13g2_a221oi_1 _1564_ (.B2(net266),
    .C1(net319),
    .B1(_0682_),
    .A1(_0100_),
    .Y(_0061_),
    .A2(_0583_));
 sg13g2_nor2_1 _1565_ (.A(net305),
    .B(_0652_),
    .Y(_0683_));
 sg13g2_mux4_1 _1566_ (.S0(net373),
    .A0(\adc_data2[11] ),
    .A1(\adc_data2[12] ),
    .A2(\adc_data2[13] ),
    .A3(\adc_data2[14] ),
    .S1(net356),
    .X(_0684_));
 sg13g2_or2_1 _1567_ (.X(_0685_),
    .B(_0684_),
    .A(net311));
 sg13g2_o21ai_1 _1568_ (.B1(_0685_),
    .Y(_0686_),
    .A1(net334),
    .A2(_0625_));
 sg13g2_o21ai_1 _1569_ (.B1(net293),
    .Y(_0687_),
    .A1(_0683_),
    .A2(_0686_));
 sg13g2_o21ai_1 _1570_ (.B1(_0687_),
    .Y(_0688_),
    .A1(net178),
    .A2(net279));
 sg13g2_a221oi_1 _1571_ (.B2(net265),
    .C1(net318),
    .B1(_0688_),
    .A1(_0099_),
    .Y(_0062_),
    .A2(_0583_));
 sg13g2_a21oi_1 _1572_ (.A1(net270),
    .A2(net281),
    .Y(_0689_),
    .B1(net124));
 sg13g2_mux2_1 _1573_ (.A0(_0219_),
    .A1(_0247_),
    .S(_0345_),
    .X(_0690_));
 sg13g2_mux2_1 _1574_ (.A0(_0218_),
    .A1(_0248_),
    .S(_0345_),
    .X(_0691_));
 sg13g2_a21oi_1 _1575_ (.A1(_0146_),
    .A2(_0353_),
    .Y(_0692_),
    .B1(_0355_));
 sg13g2_o21ai_1 _1576_ (.B1(net380),
    .Y(_0693_),
    .A1(_0691_),
    .A2(_0692_));
 sg13g2_nor2_1 _1577_ (.A(net125),
    .B(_0693_),
    .Y(_0063_));
 sg13g2_nand2_1 _1578_ (.Y(_0694_),
    .A(_0361_),
    .B(net262));
 sg13g2_nor2_1 _1579_ (.A(\adc_data3[0] ),
    .B(net362),
    .Y(_0695_));
 sg13g2_a21oi_1 _1580_ (.A1(_0098_),
    .A2(net362),
    .Y(_0696_),
    .B1(_0695_));
 sg13g2_and2_1 _1581_ (.A(net348),
    .B(_0696_),
    .X(_0697_));
 sg13g2_nand3_1 _1582_ (.B(net338),
    .C(_0697_),
    .A(net328),
    .Y(_0698_));
 sg13g2_nand2_1 _1583_ (.Y(_0699_),
    .A(net289),
    .B(_0698_));
 sg13g2_o21ai_1 _1584_ (.B1(_0699_),
    .Y(_0700_),
    .A1(net124),
    .A2(net275));
 sg13g2_a221oi_1 _1585_ (.B2(net261),
    .C1(net313),
    .B1(_0700_),
    .A1(_0098_),
    .Y(_0064_),
    .A2(net257));
 sg13g2_and2_1 _1586_ (.A(\adc_data3[0] ),
    .B(net362),
    .X(_0701_));
 sg13g2_mux2_1 _1587_ (.A0(_0098_),
    .A1(_0097_),
    .S(net362),
    .X(_0702_));
 sg13g2_nor2_1 _1588_ (.A(net348),
    .B(_0701_),
    .Y(_0703_));
 sg13g2_a21oi_1 _1589_ (.A1(net348),
    .A2(_0702_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_nand3_1 _1590_ (.B(net338),
    .C(_0704_),
    .A(net328),
    .Y(_0705_));
 sg13g2_a22oi_1 _1591_ (.Y(_0706_),
    .B1(_0705_),
    .B2(net289),
    .A2(net282),
    .A1(_0098_));
 sg13g2_o21ai_1 _1592_ (.B1(net380),
    .Y(_0707_),
    .A1(_0691_),
    .A2(_0706_));
 sg13g2_a21oi_1 _1593_ (.A1(_0097_),
    .A2(net257),
    .Y(_0065_),
    .B1(_0707_));
 sg13g2_mux2_1 _1594_ (.A0(_0097_),
    .A1(_0096_),
    .S(net362),
    .X(_0708_));
 sg13g2_nand2_1 _1595_ (.Y(_0709_),
    .A(net322),
    .B(_0696_));
 sg13g2_o21ai_1 _1596_ (.B1(_0709_),
    .Y(_0710_),
    .A1(net322),
    .A2(_0708_));
 sg13g2_and2_1 _1597_ (.A(net337),
    .B(_0710_),
    .X(_0711_));
 sg13g2_a21o_1 _1598_ (.A2(_0711_),
    .A1(net328),
    .B1(net286),
    .X(_0712_));
 sg13g2_o21ai_1 _1599_ (.B1(_0712_),
    .Y(_0713_),
    .A1(net137),
    .A2(net275));
 sg13g2_a221oi_1 _1600_ (.B2(net262),
    .C1(net313),
    .B1(_0713_),
    .A1(_0096_),
    .Y(_0066_),
    .A2(net257));
 sg13g2_nor2_1 _1601_ (.A(\adc_data3[3] ),
    .B(net362),
    .Y(_0714_));
 sg13g2_a21oi_1 _1602_ (.A1(_0095_),
    .A2(net362),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nand2_1 _1603_ (.Y(_0716_),
    .A(net348),
    .B(_0715_));
 sg13g2_o21ai_1 _1604_ (.B1(_0716_),
    .Y(_0717_),
    .A1(net348),
    .A2(_0702_));
 sg13g2_a22oi_1 _1605_ (.Y(_0718_),
    .B1(_0717_),
    .B2(net337),
    .A2(_0701_),
    .A1(_0389_));
 sg13g2_o21ai_1 _1606_ (.B1(net288),
    .Y(_0719_),
    .A1(net326),
    .A2(_0718_));
 sg13g2_o21ai_1 _1607_ (.B1(_0719_),
    .Y(_0720_),
    .A1(net177),
    .A2(net274));
 sg13g2_a221oi_1 _1608_ (.B2(net262),
    .C1(net313),
    .B1(_0720_),
    .A1(_0095_),
    .Y(_0067_),
    .A2(net258));
 sg13g2_o21ai_1 _1609_ (.B1(net154),
    .Y(_0721_),
    .A1(net272),
    .A2(_0691_));
 sg13g2_nand2_1 _1610_ (.Y(_0722_),
    .A(\adc_data3[5] ),
    .B(net361));
 sg13g2_o21ai_1 _1611_ (.B1(_0722_),
    .Y(_0723_),
    .A1(_0095_),
    .A2(net360));
 sg13g2_nand2_1 _1612_ (.Y(_0724_),
    .A(net349),
    .B(_0723_));
 sg13g2_o21ai_1 _1613_ (.B1(_0724_),
    .Y(_0725_),
    .A1(net349),
    .A2(_0708_));
 sg13g2_mux2_1 _1614_ (.A0(_0697_),
    .A1(_0725_),
    .S(net337),
    .X(_0726_));
 sg13g2_a22oi_1 _1615_ (.Y(_0727_),
    .B1(_0374_),
    .B2(_0726_),
    .A2(net282),
    .A1(\adc_data3[4] ));
 sg13g2_nand2b_1 _1616_ (.Y(_0728_),
    .B(net261),
    .A_N(_0727_));
 sg13g2_a21oi_1 _1617_ (.A1(_0721_),
    .A2(_0728_),
    .Y(_0068_),
    .B1(net312));
 sg13g2_nand2_1 _1618_ (.Y(_0729_),
    .A(_0094_),
    .B(net361));
 sg13g2_o21ai_1 _1619_ (.B1(_0729_),
    .Y(_0730_),
    .A1(\adc_data3[5] ),
    .A2(net360));
 sg13g2_nor2_1 _1620_ (.A(net347),
    .B(_0715_),
    .Y(_0731_));
 sg13g2_a21oi_1 _1621_ (.A1(net347),
    .A2(_0730_),
    .Y(_0732_),
    .B1(_0731_));
 sg13g2_mux2_1 _1622_ (.A0(_0704_),
    .A1(_0732_),
    .S(net337),
    .X(_0733_));
 sg13g2_a21o_1 _1623_ (.A2(_0733_),
    .A1(net327),
    .B1(net286),
    .X(_0734_));
 sg13g2_o21ai_1 _1624_ (.B1(_0734_),
    .Y(_0735_),
    .A1(net154),
    .A2(net274));
 sg13g2_a221oi_1 _1625_ (.B2(net261),
    .C1(net312),
    .B1(_0735_),
    .A1(_0094_),
    .Y(_0069_),
    .A2(net257));
 sg13g2_nor2_1 _1626_ (.A(\adc_data3[6] ),
    .B(net360),
    .Y(_0736_));
 sg13g2_a21oi_1 _1627_ (.A1(_0093_),
    .A2(net360),
    .Y(_0737_),
    .B1(_0736_));
 sg13g2_mux2_1 _1628_ (.A0(_0723_),
    .A1(_0737_),
    .S(net347),
    .X(_0738_));
 sg13g2_mux2_1 _1629_ (.A0(_0710_),
    .A1(_0738_),
    .S(net337),
    .X(_0739_));
 sg13g2_a21o_1 _1630_ (.A2(_0739_),
    .A1(net327),
    .B1(net286),
    .X(_0740_));
 sg13g2_o21ai_1 _1631_ (.B1(_0740_),
    .Y(_0741_),
    .A1(net196),
    .A2(net274));
 sg13g2_a221oi_1 _1632_ (.B2(net261),
    .C1(net312),
    .B1(_0741_),
    .A1(_0093_),
    .Y(_0070_),
    .A2(net257));
 sg13g2_a21oi_1 _1633_ (.A1(net124),
    .A2(_0149_),
    .Y(_0742_),
    .B1(net328));
 sg13g2_mux4_1 _1634_ (.S0(net360),
    .A0(\adc_data3[5] ),
    .A1(\adc_data3[6] ),
    .A2(\adc_data3[7] ),
    .A3(\adc_data3[8] ),
    .S1(net347),
    .X(_0743_));
 sg13g2_or2_1 _1635_ (.X(_0744_),
    .B(_0743_),
    .A(net307));
 sg13g2_o21ai_1 _1636_ (.B1(_0744_),
    .Y(_0745_),
    .A1(net304),
    .A2(_0717_));
 sg13g2_o21ai_1 _1637_ (.B1(net288),
    .Y(_0746_),
    .A1(_0742_),
    .A2(_0745_));
 sg13g2_o21ai_1 _1638_ (.B1(_0746_),
    .Y(_0747_),
    .A1(\adc_data3[7] ),
    .A2(net274));
 sg13g2_a221oi_1 _1639_ (.B2(net261),
    .C1(net312),
    .B1(_0747_),
    .A1(_0092_),
    .Y(_0071_),
    .A2(net257));
 sg13g2_a21oi_1 _1640_ (.A1(net337),
    .A2(_0697_),
    .Y(_0748_),
    .B1(net327));
 sg13g2_nor2_1 _1641_ (.A(\adc_data3[8] ),
    .B(net360),
    .Y(_0749_));
 sg13g2_a21oi_1 _1642_ (.A1(_0091_),
    .A2(net360),
    .Y(_0750_),
    .B1(_0749_));
 sg13g2_mux2_1 _1643_ (.A0(_0737_),
    .A1(_0750_),
    .S(net347),
    .X(_0751_));
 sg13g2_or2_1 _1644_ (.X(_0752_),
    .B(_0751_),
    .A(net307));
 sg13g2_o21ai_1 _1645_ (.B1(_0752_),
    .Y(_0753_),
    .A1(net304),
    .A2(_0725_));
 sg13g2_o21ai_1 _1646_ (.B1(net288),
    .Y(_0754_),
    .A1(_0748_),
    .A2(_0753_));
 sg13g2_o21ai_1 _1647_ (.B1(_0754_),
    .Y(_0755_),
    .A1(net152),
    .A2(net274));
 sg13g2_a221oi_1 _1648_ (.B2(net261),
    .C1(net312),
    .B1(_0755_),
    .A1(_0091_),
    .Y(_0072_),
    .A2(net257));
 sg13g2_a21oi_1 _1649_ (.A1(net337),
    .A2(_0704_),
    .Y(_0756_),
    .B1(net327));
 sg13g2_mux4_1 _1650_ (.S0(net360),
    .A0(\adc_data3[7] ),
    .A1(\adc_data3[8] ),
    .A2(\adc_data3[9] ),
    .A3(\adc_data3[10] ),
    .S1(net347),
    .X(_0757_));
 sg13g2_or2_1 _1651_ (.X(_0758_),
    .B(_0757_),
    .A(net307));
 sg13g2_o21ai_1 _1652_ (.B1(_0758_),
    .Y(_0759_),
    .A1(net337),
    .A2(_0732_));
 sg13g2_o21ai_1 _1653_ (.B1(net288),
    .Y(_0760_),
    .A1(_0756_),
    .A2(_0759_));
 sg13g2_o21ai_1 _1654_ (.B1(_0760_),
    .Y(_0761_),
    .A1(net174),
    .A2(net274));
 sg13g2_a221oi_1 _1655_ (.B2(net261),
    .C1(net312),
    .B1(_0761_),
    .A1(_0090_),
    .Y(_0073_),
    .A2(net257));
 sg13g2_o21ai_1 _1656_ (.B1(net164),
    .Y(_0762_),
    .A1(net272),
    .A2(_0691_));
 sg13g2_nor2_1 _1657_ (.A(_0090_),
    .B(net274),
    .Y(_0763_));
 sg13g2_nor2_1 _1658_ (.A(net327),
    .B(_0711_),
    .Y(_0764_));
 sg13g2_nor2_1 _1659_ (.A(_0090_),
    .B(net361),
    .Y(_0765_));
 sg13g2_a21oi_1 _1660_ (.A1(\adc_data3[11] ),
    .A2(net361),
    .Y(_0766_),
    .B1(_0765_));
 sg13g2_nand2_1 _1661_ (.Y(_0767_),
    .A(net322),
    .B(_0750_));
 sg13g2_o21ai_1 _1662_ (.B1(_0767_),
    .Y(_0768_),
    .A1(net322),
    .A2(_0766_));
 sg13g2_nor2_1 _1663_ (.A(net307),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_nor2_1 _1664_ (.A(net338),
    .B(_0738_),
    .Y(_0770_));
 sg13g2_nor4_1 _1665_ (.A(net286),
    .B(_0764_),
    .C(_0769_),
    .D(_0770_),
    .Y(_0771_));
 sg13g2_o21ai_1 _1666_ (.B1(net261),
    .Y(_0772_),
    .A1(_0763_),
    .A2(_0771_));
 sg13g2_a21oi_1 _1667_ (.A1(_0762_),
    .A2(_0772_),
    .Y(_0074_),
    .B1(net312));
 sg13g2_o21ai_1 _1668_ (.B1(net158),
    .Y(_0773_),
    .A1(net272),
    .A2(_0691_));
 sg13g2_mux4_1 _1669_ (.S0(net361),
    .A0(\adc_data3[9] ),
    .A1(\adc_data3[10] ),
    .A2(\adc_data3[11] ),
    .A3(\adc_data3[12] ),
    .S1(net347),
    .X(_0774_));
 sg13g2_or2_1 _1670_ (.X(_0775_),
    .B(_0774_),
    .A(net307));
 sg13g2_o21ai_1 _1671_ (.B1(_0775_),
    .Y(_0776_),
    .A1(net304),
    .A2(_0743_));
 sg13g2_a21oi_1 _1672_ (.A1(net326),
    .A2(_0718_),
    .Y(_0777_),
    .B1(_0776_));
 sg13g2_a22oi_1 _1673_ (.Y(_0778_),
    .B1(_0777_),
    .B2(net288),
    .A2(net282),
    .A1(\adc_data3[11] ));
 sg13g2_nand2b_1 _1674_ (.Y(_0779_),
    .B(net262),
    .A_N(_0778_));
 sg13g2_a21oi_1 _1675_ (.A1(_0773_),
    .A2(_0779_),
    .Y(_0075_),
    .B1(net312));
 sg13g2_nor2_1 _1676_ (.A(net327),
    .B(_0726_),
    .Y(_0780_));
 sg13g2_nor2_1 _1677_ (.A(\adc_data3[12] ),
    .B(net363),
    .Y(_0781_));
 sg13g2_a21oi_1 _1678_ (.A1(_0089_),
    .A2(net363),
    .Y(_0782_),
    .B1(_0781_));
 sg13g2_a21oi_1 _1679_ (.A1(net347),
    .A2(_0782_),
    .Y(_0783_),
    .B1(net307));
 sg13g2_o21ai_1 _1680_ (.B1(_0783_),
    .Y(_0784_),
    .A1(net348),
    .A2(_0766_));
 sg13g2_o21ai_1 _1681_ (.B1(_0784_),
    .Y(_0785_),
    .A1(net304),
    .A2(_0751_));
 sg13g2_o21ai_1 _1682_ (.B1(net288),
    .Y(_0786_),
    .A1(_0780_),
    .A2(_0785_));
 sg13g2_o21ai_1 _1683_ (.B1(_0786_),
    .Y(_0787_),
    .A1(net158),
    .A2(net274));
 sg13g2_a221oi_1 _1684_ (.B2(net262),
    .C1(net314),
    .B1(_0787_),
    .A1(_0089_),
    .Y(_0076_),
    .A2(net258));
 sg13g2_nor2_1 _1685_ (.A(net327),
    .B(_0733_),
    .Y(_0788_));
 sg13g2_mux4_1 _1686_ (.S0(net363),
    .A0(\adc_data3[11] ),
    .A1(\adc_data3[12] ),
    .A2(\adc_data3[13] ),
    .A3(\adc_data3[14] ),
    .S1(net354),
    .X(_0789_));
 sg13g2_or2_1 _1687_ (.X(_0790_),
    .B(_0789_),
    .A(net307));
 sg13g2_o21ai_1 _1688_ (.B1(_0790_),
    .Y(_0791_),
    .A1(net304),
    .A2(_0757_));
 sg13g2_o21ai_1 _1689_ (.B1(net288),
    .Y(_0792_),
    .A1(_0788_),
    .A2(_0791_));
 sg13g2_o21ai_1 _1690_ (.B1(_0792_),
    .Y(_0793_),
    .A1(\adc_data3[13] ),
    .A2(net275));
 sg13g2_a221oi_1 _1691_ (.B2(net262),
    .C1(net314),
    .B1(_0793_),
    .A1(_0088_),
    .Y(_0077_),
    .A2(net258));
 sg13g2_nor2_1 _1692_ (.A(_0161_),
    .B(net287),
    .Y(_0794_));
 sg13g2_nand2_2 _1693_ (.Y(_0795_),
    .A(_0160_),
    .B(net291));
 sg13g2_a21oi_1 _1694_ (.A1(net271),
    .A2(_0795_),
    .Y(_0796_),
    .B1(net117));
 sg13g2_a221oi_1 _1695_ (.B2(net325),
    .C1(net308),
    .B1(_0458_),
    .A1(\adc_data0[14] ),
    .Y(_0797_),
    .A2(_0186_));
 sg13g2_or2_1 _1696_ (.X(_0798_),
    .B(_0443_),
    .A(net306));
 sg13g2_o21ai_1 _1697_ (.B1(_0798_),
    .Y(_0799_),
    .A1(net330),
    .A2(_0414_));
 sg13g2_o21ai_1 _1698_ (.B1(net290),
    .Y(_0800_),
    .A1(_0797_),
    .A2(_0799_));
 sg13g2_a22oi_1 _1699_ (.Y(_0801_),
    .B1(net272),
    .B2(_0087_),
    .A2(net283),
    .A1(_0120_));
 sg13g2_a221oi_1 _1700_ (.B2(_0801_),
    .C1(_0347_),
    .B1(_0800_),
    .A1(_0160_),
    .Y(_0802_),
    .A2(net291));
 sg13g2_nor3_1 _1701_ (.A(net317),
    .B(_0796_),
    .C(_0802_),
    .Y(_0078_));
 sg13g2_nor2_1 _1702_ (.A(net305),
    .B(_0550_),
    .Y(_0803_));
 sg13g2_a221oi_1 _1703_ (.B2(net323),
    .C1(net310),
    .B1(_0564_),
    .A1(\adc_data1[14] ),
    .Y(_0804_),
    .A2(_0186_));
 sg13g2_nor2_1 _1704_ (.A(_0803_),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_o21ai_1 _1705_ (.B1(_0805_),
    .Y(_0806_),
    .A1(net332),
    .A2(_0521_));
 sg13g2_nor3_1 _1706_ (.A(net106),
    .B(net289),
    .C(net282),
    .Y(_0807_));
 sg13g2_a221oi_1 _1707_ (.B2(net292),
    .C1(_0807_),
    .B1(_0806_),
    .A1(_0109_),
    .Y(_0808_),
    .A2(net284));
 sg13g2_nor3_1 _1708_ (.A(_0472_),
    .B(_0794_),
    .C(_0808_),
    .Y(_0809_));
 sg13g2_a21oi_1 _1709_ (.A1(net267),
    .A2(_0795_),
    .Y(_0810_),
    .B1(net106));
 sg13g2_nor3_1 _1710_ (.A(net313),
    .B(_0809_),
    .C(_0810_),
    .Y(_0079_));
 sg13g2_nor2_1 _1711_ (.A(net305),
    .B(_0662_),
    .Y(_0811_));
 sg13g2_a221oi_1 _1712_ (.B2(net323),
    .C1(net310),
    .B1(_0677_),
    .A1(\adc_data2[14] ),
    .Y(_0812_),
    .A2(_0186_));
 sg13g2_nor2_1 _1713_ (.A(_0811_),
    .B(_0812_),
    .Y(_0813_));
 sg13g2_o21ai_1 _1714_ (.B1(_0813_),
    .Y(_0814_),
    .A1(net334),
    .A2(_0632_));
 sg13g2_a22oi_1 _1715_ (.Y(_0815_),
    .B1(_0814_),
    .B2(net293),
    .A2(net285),
    .A1(_0099_));
 sg13g2_o21ai_1 _1716_ (.B1(_0815_),
    .Y(_0816_),
    .A1(net112),
    .A2(_0361_));
 sg13g2_and3_1 _1717_ (.X(_0817_),
    .A(net265),
    .B(_0795_),
    .C(_0816_));
 sg13g2_a21oi_1 _1718_ (.A1(net265),
    .A2(_0795_),
    .Y(_0818_),
    .B1(net112));
 sg13g2_nor3_1 _1719_ (.A(net318),
    .B(_0817_),
    .C(_0818_),
    .Y(_0080_));
 sg13g2_nor3_1 _1720_ (.A(net119),
    .B(net289),
    .C(net282),
    .Y(_0819_));
 sg13g2_nor2_1 _1721_ (.A(net304),
    .B(_0768_),
    .Y(_0820_));
 sg13g2_a221oi_1 _1722_ (.B2(net322),
    .C1(net307),
    .B1(_0782_),
    .A1(\adc_data3[14] ),
    .Y(_0821_),
    .A2(_0186_));
 sg13g2_nor2_1 _1723_ (.A(_0820_),
    .B(_0821_),
    .Y(_0082_));
 sg13g2_o21ai_1 _1724_ (.B1(_0082_),
    .Y(_0083_),
    .A1(net327),
    .A2(_0739_));
 sg13g2_a221oi_1 _1725_ (.B2(net289),
    .C1(_0819_),
    .B1(_0083_),
    .A1(_0088_),
    .Y(_0084_),
    .A2(net282));
 sg13g2_nor3_1 _1726_ (.A(_0691_),
    .B(_0794_),
    .C(_0084_),
    .Y(_0085_));
 sg13g2_a21oi_1 _1727_ (.A1(net262),
    .A2(_0795_),
    .Y(_0086_),
    .B1(net119));
 sg13g2_nor3_1 _1728_ (.A(net314),
    .B(_0085_),
    .C(_0086_),
    .Y(_0081_));
 sg13g2_dfrbpq_2 _1729_ (.RESET_B(net34),
    .D(_0000_),
    .Q(\cycle[0] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_2 _1730_ (.RESET_B(net69),
    .D(net130),
    .Q(\cycle[1] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_2 _1731_ (.RESET_B(net67),
    .D(net209),
    .Q(\cycle[2] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_2 _1732_ (.RESET_B(net65),
    .D(_0003_),
    .Q(\cycle[3] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_2 _1733_ (.RESET_B(net63),
    .D(_0004_),
    .Q(\cycle[4] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_2 _1734_ (.RESET_B(net61),
    .D(_0005_),
    .Q(\cycle[5] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_2 _1735_ (.RESET_B(net59),
    .D(_0006_),
    .Q(\tx_cycle[0] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _1736_ (.RESET_B(net57),
    .D(_0007_),
    .Q(\tx_cycle[1] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_1 _1737_ (.RESET_B(net55),
    .D(_0008_),
    .Q(\tx_cycle[2] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_2 _1738_ (.RESET_B(net53),
    .D(_0009_),
    .Q(\tx_cycle[3] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_2 _1739_ (.RESET_B(net51),
    .D(_0010_),
    .Q(\tx_cycle[4] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_2 _1740_ (.RESET_B(net49),
    .D(_0011_),
    .Q(\tx_cycle[5] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_2 _1741_ (.RESET_B(net47),
    .D(_0012_),
    .Q(\tx_cycle[6] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_2 _1742_ (.RESET_B(net45),
    .D(_0013_),
    .Q(adc_sclk),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_2 _1743_ (.RESET_B(net43),
    .D(_0014_),
    .Q(\clk_div[0] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_2 _1744_ (.RESET_B(net41),
    .D(_0015_),
    .Q(\clk_div[1] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_2 _1745_ (.RESET_B(net39),
    .D(_0016_),
    .Q(\clk_div[2] ),
    .CLK(clknet_4_15_0_clk_regs));
 sg13g2_dfrbpq_1 _1746_ (.RESET_B(net37),
    .D(_0017_),
    .Q(\clk_div[3] ),
    .CLK(clknet_4_13_0_clk_regs));
 sg13g2_dfrbpq_2 _1747_ (.RESET_B(net35),
    .D(_0018_),
    .Q(\adc_data0[0] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _1748_ (.RESET_B(net33),
    .D(_0019_),
    .Q(\adc_data0[1] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _1749_ (.RESET_B(net31),
    .D(net116),
    .Q(\adc_data0[2] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_1 _1750_ (.RESET_B(net29),
    .D(_0021_),
    .Q(\adc_data0[3] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _1751_ (.RESET_B(net27),
    .D(_0022_),
    .Q(\adc_data0[4] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_2 _1752_ (.RESET_B(net25),
    .D(_0023_),
    .Q(\adc_data0[5] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_2 _1753_ (.RESET_B(net23),
    .D(_0024_),
    .Q(\adc_data0[6] ),
    .CLK(clknet_4_7_0_clk_regs));
 sg13g2_dfrbpq_2 _1754_ (.RESET_B(net21),
    .D(net191),
    .Q(\adc_data0[7] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_2 _1755_ (.RESET_B(net101),
    .D(net151),
    .Q(\adc_data0[8] ),
    .CLK(clknet_4_5_0_clk_regs));
 sg13g2_dfrbpq_1 _1756_ (.RESET_B(net99),
    .D(_0027_),
    .Q(\adc_data0[9] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_2 _1757_ (.RESET_B(net97),
    .D(net157),
    .Q(\adc_data0[10] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_2 _1758_ (.RESET_B(net95),
    .D(_0029_),
    .Q(\adc_data0[11] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_2 _1759_ (.RESET_B(net93),
    .D(_0030_),
    .Q(\adc_data0[12] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_2 _1760_ (.RESET_B(net91),
    .D(net135),
    .Q(\adc_data0[13] ),
    .CLK(clknet_4_4_0_clk_regs));
 sg13g2_dfrbpq_1 _1761_ (.RESET_B(net89),
    .D(_0032_),
    .Q(\adc_data0[14] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_2 _1762_ (.RESET_B(net87),
    .D(_0033_),
    .Q(\adc_data1[0] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _1763_ (.RESET_B(net85),
    .D(_0034_),
    .Q(\adc_data1[1] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _1764_ (.RESET_B(net83),
    .D(_0035_),
    .Q(\adc_data1[2] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _1765_ (.RESET_B(net81),
    .D(_0036_),
    .Q(\adc_data1[3] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _1766_ (.RESET_B(net79),
    .D(net167),
    .Q(\adc_data1[4] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_2 _1767_ (.RESET_B(net77),
    .D(_0038_),
    .Q(\adc_data1[5] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _1768_ (.RESET_B(net75),
    .D(_0039_),
    .Q(\adc_data1[6] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_2 _1769_ (.RESET_B(net73),
    .D(net187),
    .Q(\adc_data1[7] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_2 _1770_ (.RESET_B(net71),
    .D(net163),
    .Q(\adc_data1[8] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _1771_ (.RESET_B(net68),
    .D(_0042_),
    .Q(\adc_data1[9] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_2 _1772_ (.RESET_B(net64),
    .D(net184),
    .Q(\adc_data1[10] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _1773_ (.RESET_B(net60),
    .D(_0044_),
    .Q(\adc_data1[11] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_2 _1774_ (.RESET_B(net56),
    .D(net148),
    .Q(\adc_data1[12] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _1775_ (.RESET_B(net52),
    .D(_0046_),
    .Q(\adc_data1[13] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _1776_ (.RESET_B(net48),
    .D(_0047_),
    .Q(\adc_data1[14] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_2 _1777_ (.RESET_B(net44),
    .D(_0048_),
    .Q(\adc_data2[0] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _1778_ (.RESET_B(net40),
    .D(_0049_),
    .Q(\adc_data2[1] ),
    .CLK(clknet_4_12_0_clk_regs));
 sg13g2_dfrbpq_1 _1779_ (.RESET_B(net36),
    .D(net109),
    .Q(\adc_data2[2] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_1 _1780_ (.RESET_B(net32),
    .D(_0051_),
    .Q(\adc_data2[3] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_2 _1781_ (.RESET_B(net28),
    .D(net140),
    .Q(\adc_data2[4] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_2 _1782_ (.RESET_B(net24),
    .D(_0053_),
    .Q(\adc_data2[5] ),
    .CLK(clknet_4_14_0_clk_regs));
 sg13g2_dfrbpq_2 _1783_ (.RESET_B(net20),
    .D(net144),
    .Q(\adc_data2[6] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_2 _1784_ (.RESET_B(net98),
    .D(net133),
    .Q(\adc_data2[7] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_2 _1785_ (.RESET_B(net94),
    .D(_0056_),
    .Q(\adc_data2[8] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_2 _1786_ (.RESET_B(net90),
    .D(_0057_),
    .Q(\adc_data2[9] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_2 _1787_ (.RESET_B(net86),
    .D(_0058_),
    .Q(\adc_data2[10] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_2 _1788_ (.RESET_B(net82),
    .D(net161),
    .Q(\adc_data2[11] ),
    .CLK(clknet_4_11_0_clk_regs));
 sg13g2_dfrbpq_2 _1789_ (.RESET_B(net78),
    .D(_0060_),
    .Q(\adc_data2[12] ),
    .CLK(clknet_4_10_0_clk_regs));
 sg13g2_dfrbpq_1 _1790_ (.RESET_B(net74),
    .D(_0061_),
    .Q(\adc_data2[13] ),
    .CLK(clknet_4_8_0_clk_regs));
 sg13g2_dfrbpq_1 _1791_ (.RESET_B(net70),
    .D(_0062_),
    .Q(\adc_data2[14] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_2 _1792_ (.RESET_B(net62),
    .D(_0063_),
    .Q(\adc_data3[0] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _1793_ (.RESET_B(net54),
    .D(_0064_),
    .Q(\adc_data3[1] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _1794_ (.RESET_B(net46),
    .D(_0065_),
    .Q(\adc_data3[2] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _1795_ (.RESET_B(net38),
    .D(_0066_),
    .Q(\adc_data3[3] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _1796_ (.RESET_B(net30),
    .D(_0067_),
    .Q(\adc_data3[4] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_2 _1797_ (.RESET_B(net22),
    .D(net155),
    .Q(\adc_data3[5] ),
    .CLK(clknet_4_1_0_clk_regs));
 sg13g2_dfrbpq_1 _1798_ (.RESET_B(net96),
    .D(_0069_),
    .Q(\adc_data3[6] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _1799_ (.RESET_B(net88),
    .D(_0070_),
    .Q(\adc_data3[7] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_2 _1800_ (.RESET_B(net80),
    .D(net153),
    .Q(\adc_data3[8] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_2 _1801_ (.RESET_B(net72),
    .D(_0072_),
    .Q(\adc_data3[9] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_1 _1802_ (.RESET_B(net58),
    .D(_0073_),
    .Q(\adc_data3[10] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_2 _1803_ (.RESET_B(net42),
    .D(net165),
    .Q(\adc_data3[11] ),
    .CLK(clknet_4_0_0_clk_regs));
 sg13g2_dfrbpq_2 _1804_ (.RESET_B(net26),
    .D(net159),
    .Q(\adc_data3[12] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _1805_ (.RESET_B(net92),
    .D(_0076_),
    .Q(\adc_data3[13] ),
    .CLK(clknet_4_2_0_clk_regs));
 sg13g2_dfrbpq_1 _1806_ (.RESET_B(net76),
    .D(net173),
    .Q(\adc_data3[14] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_dfrbpq_1 _1807_ (.RESET_B(net50),
    .D(net118),
    .Q(\adc_data0[15] ),
    .CLK(clknet_4_6_0_clk_regs));
 sg13g2_dfrbpq_1 _1808_ (.RESET_B(net100),
    .D(net107),
    .Q(\adc_data1[15] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _1809_ (.RESET_B(net66),
    .D(_0080_),
    .Q(\adc_data2[15] ),
    .CLK(clknet_4_9_0_clk_regs));
 sg13g2_dfrbpq_1 _1810_ (.RESET_B(net84),
    .D(net120),
    .Q(\adc_data3[15] ),
    .CLK(clknet_4_3_0_clk_regs));
 sg13g2_tiehi _1754__21 (.L_HI(net21));
 sg13g2_tiehi _1797__22 (.L_HI(net22));
 sg13g2_tiehi _1753__23 (.L_HI(net23));
 sg13g2_tiehi _1782__24 (.L_HI(net24));
 sg13g2_tiehi _1752__25 (.L_HI(net25));
 sg13g2_tiehi _1804__26 (.L_HI(net26));
 sg13g2_tiehi _1751__27 (.L_HI(net27));
 sg13g2_tiehi _1781__28 (.L_HI(net28));
 sg13g2_tiehi _1750__29 (.L_HI(net29));
 sg13g2_tiehi _1796__30 (.L_HI(net30));
 sg13g2_tiehi _1749__31 (.L_HI(net31));
 sg13g2_tiehi _1780__32 (.L_HI(net32));
 sg13g2_tiehi _1748__33 (.L_HI(net33));
 sg13g2_tiehi _1729__34 (.L_HI(net34));
 sg13g2_tiehi _1747__35 (.L_HI(net35));
 sg13g2_tiehi _1779__36 (.L_HI(net36));
 sg13g2_tiehi _1746__37 (.L_HI(net37));
 sg13g2_tiehi _1795__38 (.L_HI(net38));
 sg13g2_tiehi _1745__39 (.L_HI(net39));
 sg13g2_tiehi _1778__40 (.L_HI(net40));
 sg13g2_tiehi _1744__41 (.L_HI(net41));
 sg13g2_tiehi _1803__42 (.L_HI(net42));
 sg13g2_tiehi _1743__43 (.L_HI(net43));
 sg13g2_tiehi _1777__44 (.L_HI(net44));
 sg13g2_tiehi _1742__45 (.L_HI(net45));
 sg13g2_tiehi _1794__46 (.L_HI(net46));
 sg13g2_tiehi _1741__47 (.L_HI(net47));
 sg13g2_tiehi _1776__48 (.L_HI(net48));
 sg13g2_tiehi _1740__49 (.L_HI(net49));
 sg13g2_tiehi _1807__50 (.L_HI(net50));
 sg13g2_tiehi _1739__51 (.L_HI(net51));
 sg13g2_tiehi _1775__52 (.L_HI(net52));
 sg13g2_tiehi _1738__53 (.L_HI(net53));
 sg13g2_tiehi _1793__54 (.L_HI(net54));
 sg13g2_tiehi _1737__55 (.L_HI(net55));
 sg13g2_tiehi _1774__56 (.L_HI(net56));
 sg13g2_tiehi _1736__57 (.L_HI(net57));
 sg13g2_tiehi _1802__58 (.L_HI(net58));
 sg13g2_tiehi _1735__59 (.L_HI(net59));
 sg13g2_tiehi _1773__60 (.L_HI(net60));
 sg13g2_tiehi _1734__61 (.L_HI(net61));
 sg13g2_tiehi _1792__62 (.L_HI(net62));
 sg13g2_tiehi _1733__63 (.L_HI(net63));
 sg13g2_tiehi _1772__64 (.L_HI(net64));
 sg13g2_tiehi _1732__65 (.L_HI(net65));
 sg13g2_tiehi _1809__66 (.L_HI(net66));
 sg13g2_tiehi _1731__67 (.L_HI(net67));
 sg13g2_tiehi _1771__68 (.L_HI(net68));
 sg13g2_tiehi _1730__69 (.L_HI(net69));
 sg13g2_tiehi _1791__70 (.L_HI(net70));
 sg13g2_tiehi _1770__71 (.L_HI(net71));
 sg13g2_tiehi _1801__72 (.L_HI(net72));
 sg13g2_tiehi _1769__73 (.L_HI(net73));
 sg13g2_tiehi _1790__74 (.L_HI(net74));
 sg13g2_tiehi _1768__75 (.L_HI(net75));
 sg13g2_tiehi _1806__76 (.L_HI(net76));
 sg13g2_tiehi _1767__77 (.L_HI(net77));
 sg13g2_tiehi _1789__78 (.L_HI(net78));
 sg13g2_tiehi _1766__79 (.L_HI(net79));
 sg13g2_tiehi _1800__80 (.L_HI(net80));
 sg13g2_tiehi _1765__81 (.L_HI(net81));
 sg13g2_tiehi _1788__82 (.L_HI(net82));
 sg13g2_tiehi _1764__83 (.L_HI(net83));
 sg13g2_tiehi _1810__84 (.L_HI(net84));
 sg13g2_tiehi _1763__85 (.L_HI(net85));
 sg13g2_tiehi _1787__86 (.L_HI(net86));
 sg13g2_tiehi _1762__87 (.L_HI(net87));
 sg13g2_tiehi _1799__88 (.L_HI(net88));
 sg13g2_tiehi _1761__89 (.L_HI(net89));
 sg13g2_tiehi _1786__90 (.L_HI(net90));
 sg13g2_tiehi _1760__91 (.L_HI(net91));
 sg13g2_tiehi _1805__92 (.L_HI(net92));
 sg13g2_tiehi _1759__93 (.L_HI(net93));
 sg13g2_tiehi _1785__94 (.L_HI(net94));
 sg13g2_tiehi _1758__95 (.L_HI(net95));
 sg13g2_tiehi _1798__96 (.L_HI(net96));
 sg13g2_tiehi _1757__97 (.L_HI(net97));
 sg13g2_tiehi _1784__98 (.L_HI(net98));
 sg13g2_tiehi _1756__99 (.L_HI(net99));
 sg13g2_tiehi _1808__100 (.L_HI(net100));
 sg13g2_tiehi _1755__101 (.L_HI(net101));
 sg13g2_tiehi tt_um_spi_aggregator_102 (.L_HI(net102));
 sg13g2_tiehi tt_um_spi_aggregator_103 (.L_HI(net103));
 sg13g2_tiehi tt_um_spi_aggregator_104 (.L_HI(net104));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_tielo tt_um_spi_aggregator_11 (.L_LO(net11));
 sg13g2_tielo tt_um_spi_aggregator_12 (.L_LO(net12));
 sg13g2_tielo tt_um_spi_aggregator_13 (.L_LO(net13));
 sg13g2_tielo tt_um_spi_aggregator_14 (.L_LO(net14));
 sg13g2_tielo tt_um_spi_aggregator_15 (.L_LO(net15));
 sg13g2_tielo tt_um_spi_aggregator_16 (.L_LO(net16));
 sg13g2_tielo tt_um_spi_aggregator_17 (.L_LO(net17));
 sg13g2_tielo tt_um_spi_aggregator_18 (.L_LO(net18));
 sg13g2_tielo tt_um_spi_aggregator_19 (.L_LO(net19));
 sg13g2_tiehi _1783__20 (.L_HI(net20));
 sg13g2_buf_1 _1906_ (.A(net299),
    .X(uio_out[4]));
 sg13g2_buf_1 _1907_ (.A(net296),
    .X(uio_out[5]));
 sg13g2_buf_1 _1908_ (.A(tx_cs_n),
    .X(uio_out[6]));
 sg13g2_buf_1 _1909_ (.A(net299),
    .X(uo_out[0]));
 sg13g2_buf_1 _1910_ (.A(adc_cs_n),
    .X(uo_out[1]));
 sg13g2_buf_1 _1911_ (.A(net299),
    .X(uo_out[2]));
 sg13g2_buf_1 _1912_ (.A(tx_mosi),
    .X(uo_out[3]));
 sg13g2_buf_1 _1913_ (.A(clknet_1_0__leaf_clk),
    .X(uo_out[4]));
 sg13g2_buf_1 _1914_ (.A(tx_cs_n),
    .X(uo_out[5]));
 sg13g2_buf_1 _1915_ (.A(net299),
    .X(uo_out[6]));
 sg13g2_buf_1 _1916_ (.A(tx_cs_n),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout257 (.A(net258),
    .X(net257));
 sg13g2_buf_1 fanout258 (.A(_0694_),
    .X(net258));
 sg13g2_buf_8 fanout259 (.A(_0475_),
    .X(net259));
 sg13g2_buf_8 fanout260 (.A(_0362_),
    .X(net260));
 sg13g2_buf_8 fanout261 (.A(net262),
    .X(net261));
 sg13g2_buf_8 fanout262 (.A(_0690_),
    .X(net262));
 sg13g2_buf_8 fanout263 (.A(net264),
    .X(net263));
 sg13g2_buf_8 fanout264 (.A(_0580_),
    .X(net264));
 sg13g2_buf_8 fanout265 (.A(_0579_),
    .X(net265));
 sg13g2_buf_1 fanout266 (.A(_0579_),
    .X(net266));
 sg13g2_buf_8 fanout267 (.A(_0471_),
    .X(net267));
 sg13g2_buf_8 fanout268 (.A(_0471_),
    .X(net268));
 sg13g2_buf_8 fanout269 (.A(net270),
    .X(net269));
 sg13g2_buf_8 fanout270 (.A(net271),
    .X(net270));
 sg13g2_buf_8 fanout271 (.A(_0346_),
    .X(net271));
 sg13g2_buf_8 fanout272 (.A(_0360_),
    .X(net272));
 sg13g2_buf_8 fanout273 (.A(_0360_),
    .X(net273));
 sg13g2_buf_8 fanout274 (.A(net275),
    .X(net274));
 sg13g2_buf_8 fanout275 (.A(net280),
    .X(net275));
 sg13g2_buf_8 fanout276 (.A(net277),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(net280),
    .X(net277));
 sg13g2_buf_8 fanout278 (.A(net280),
    .X(net278));
 sg13g2_buf_1 fanout279 (.A(net280),
    .X(net279));
 sg13g2_buf_8 fanout280 (.A(_0358_),
    .X(net280));
 sg13g2_buf_8 fanout281 (.A(_0353_),
    .X(net281));
 sg13g2_buf_8 fanout282 (.A(_0359_),
    .X(net282));
 sg13g2_buf_1 fanout283 (.A(_0359_),
    .X(net283));
 sg13g2_buf_8 fanout284 (.A(net285),
    .X(net284));
 sg13g2_buf_8 fanout285 (.A(_0359_),
    .X(net285));
 sg13g2_buf_8 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_8 fanout287 (.A(_0275_),
    .X(net287));
 sg13g2_buf_8 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_8 fanout289 (.A(_0274_),
    .X(net289));
 sg13g2_buf_8 fanout290 (.A(net291),
    .X(net290));
 sg13g2_buf_8 fanout291 (.A(_0274_),
    .X(net291));
 sg13g2_buf_8 fanout292 (.A(net293),
    .X(net292));
 sg13g2_buf_8 fanout293 (.A(net294),
    .X(net293));
 sg13g2_buf_8 fanout294 (.A(_0274_),
    .X(net294));
 sg13g2_buf_8 fanout295 (.A(_0193_),
    .X(net295));
 sg13g2_buf_8 fanout296 (.A(adc_cs_n),
    .X(net296));
 sg13g2_buf_8 fanout297 (.A(_0183_),
    .X(net297));
 sg13g2_buf_8 fanout298 (.A(_0163_),
    .X(net298));
 sg13g2_buf_8 fanout299 (.A(net222),
    .X(net299));
 sg13g2_buf_8 fanout300 (.A(net219),
    .X(net300));
 sg13g2_buf_8 fanout301 (.A(net221),
    .X(net301));
 sg13g2_buf_8 fanout302 (.A(net220),
    .X(net302));
 sg13g2_buf_8 fanout303 (.A(net218),
    .X(net303));
 sg13g2_buf_8 fanout304 (.A(net306),
    .X(net304));
 sg13g2_buf_8 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_8 fanout306 (.A(_0429_),
    .X(net306));
 sg13g2_buf_8 fanout307 (.A(_0159_),
    .X(net307));
 sg13g2_buf_8 fanout308 (.A(_0159_),
    .X(net308));
 sg13g2_buf_8 fanout309 (.A(net310),
    .X(net309));
 sg13g2_buf_8 fanout310 (.A(net311),
    .X(net310));
 sg13g2_buf_8 fanout311 (.A(_0159_),
    .X(net311));
 sg13g2_buf_8 fanout312 (.A(net313),
    .X(net312));
 sg13g2_buf_8 fanout313 (.A(net321),
    .X(net313));
 sg13g2_buf_1 fanout314 (.A(net321),
    .X(net314));
 sg13g2_buf_8 fanout315 (.A(net317),
    .X(net315));
 sg13g2_buf_1 fanout316 (.A(net317),
    .X(net316));
 sg13g2_buf_8 fanout317 (.A(net321),
    .X(net317));
 sg13g2_buf_8 fanout318 (.A(net319),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(net320),
    .X(net319));
 sg13g2_buf_8 fanout320 (.A(net321),
    .X(net320));
 sg13g2_buf_8 fanout321 (.A(_0147_),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(net325),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(net325),
    .X(net323));
 sg13g2_buf_2 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_8 fanout325 (.A(_0141_),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(_0140_),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(net331),
    .X(net327));
 sg13g2_buf_8 fanout328 (.A(net331),
    .X(net328));
 sg13g2_buf_8 fanout329 (.A(net330),
    .X(net329));
 sg13g2_buf_1 fanout330 (.A(net331),
    .X(net330));
 sg13g2_buf_8 fanout331 (.A(ui_in[3]),
    .X(net331));
 sg13g2_buf_8 fanout332 (.A(net334),
    .X(net332));
 sg13g2_buf_1 fanout333 (.A(net334),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(net336),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(net336),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(ui_in[3]),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(net338),
    .X(net337));
 sg13g2_buf_8 fanout338 (.A(ui_in[2]),
    .X(net338));
 sg13g2_buf_8 fanout339 (.A(net340),
    .X(net339));
 sg13g2_buf_8 fanout340 (.A(net341),
    .X(net340));
 sg13g2_buf_8 fanout341 (.A(ui_in[2]),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(net343),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(net346),
    .X(net343));
 sg13g2_buf_8 fanout344 (.A(net345),
    .X(net344));
 sg13g2_buf_1 fanout345 (.A(net346),
    .X(net345));
 sg13g2_buf_8 fanout346 (.A(ui_in[2]),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(net349),
    .X(net348));
 sg13g2_buf_8 fanout349 (.A(net354),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net351),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(net352),
    .X(net351));
 sg13g2_buf_8 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_1 fanout353 (.A(net354),
    .X(net353));
 sg13g2_buf_8 fanout354 (.A(ui_in[1]),
    .X(net354));
 sg13g2_buf_8 fanout355 (.A(net357),
    .X(net355));
 sg13g2_buf_8 fanout356 (.A(net357),
    .X(net356));
 sg13g2_buf_8 fanout357 (.A(ui_in[1]),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(net359),
    .X(net358));
 sg13g2_buf_8 fanout359 (.A(ui_in[1]),
    .X(net359));
 sg13g2_buf_8 fanout360 (.A(net361),
    .X(net360));
 sg13g2_buf_8 fanout361 (.A(net362),
    .X(net361));
 sg13g2_buf_8 fanout362 (.A(net378),
    .X(net362));
 sg13g2_buf_8 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net378),
    .X(net364));
 sg13g2_buf_8 fanout365 (.A(net368),
    .X(net365));
 sg13g2_buf_8 fanout366 (.A(net368),
    .X(net366));
 sg13g2_buf_1 fanout367 (.A(net368),
    .X(net367));
 sg13g2_buf_8 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_1 fanout369 (.A(net378),
    .X(net369));
 sg13g2_buf_8 fanout370 (.A(net371),
    .X(net370));
 sg13g2_buf_8 fanout371 (.A(net378),
    .X(net371));
 sg13g2_buf_8 fanout372 (.A(net373),
    .X(net372));
 sg13g2_buf_8 fanout373 (.A(net374),
    .X(net373));
 sg13g2_buf_8 fanout374 (.A(net378),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(net377),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(net378),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(ui_in[0]),
    .X(net378));
 sg13g2_buf_8 fanout379 (.A(net380),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(net1),
    .X(net380));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_tielo tt_um_spi_aggregator_10 (.L_LO(net10));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_8_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_8_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_9_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_9_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_10_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_10_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_11_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_11_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_12_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_12_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_13_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_13_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_14_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_14_0_clk_regs));
 sg13g2_buf_8 clkbuf_4_15_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_4_15_0_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk_regs));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk_regs));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk_regs));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk_regs));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk_regs));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk_regs));
 sg13g2_inv_1 clkload7 (.A(clknet_4_9_0_clk_regs));
 sg13g2_inv_1 clkload8 (.A(clknet_4_10_0_clk_regs));
 sg13g2_inv_1 clkload9 (.A(clknet_4_11_0_clk_regs));
 sg13g2_inv_1 clkload10 (.A(clknet_4_12_0_clk_regs));
 sg13g2_inv_1 clkload11 (.A(clknet_4_13_0_clk_regs));
 sg13g2_inv_1 clkload12 (.A(clknet_4_14_0_clk_regs));
 sg13g2_inv_1 clkload13 (.A(clknet_4_15_0_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\cycle[5] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold2 (.A(\adc_data1[15] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold3 (.A(_0079_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold4 (.A(\adc_data2[2] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0050_),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold6 (.A(\cycle[4] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0258_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold8 (.A(\adc_data2[15] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold9 (.A(\adc_data2[0] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0576_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold11 (.A(\adc_data0[2] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0020_),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold13 (.A(\adc_data0[15] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0078_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold15 (.A(\adc_data3[15] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0081_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold17 (.A(\adc_data1[0] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold18 (.A(_0470_),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold19 (.A(\adc_data1[1] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold20 (.A(\adc_data3[0] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0689_),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold22 (.A(\adc_data0[0] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0354_),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold24 (.A(\cycle[1] ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0252_),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0001_),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold27 (.A(\adc_data3[1] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold28 (.A(\adc_data2[7] ),
    .X(net132));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0055_),
    .X(net133));
 sg13g2_dlygate4sd3_1 hold30 (.A(\adc_data0[13] ),
    .X(net134));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0031_),
    .X(net135));
 sg13g2_dlygate4sd3_1 hold32 (.A(\adc_data2[1] ),
    .X(net136));
 sg13g2_dlygate4sd3_1 hold33 (.A(\adc_data3[2] ),
    .X(net137));
 sg13g2_dlygate4sd3_1 hold34 (.A(\adc_data1[2] ),
    .X(net138));
 sg13g2_dlygate4sd3_1 hold35 (.A(\adc_data2[4] ),
    .X(net139));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0052_),
    .X(net140));
 sg13g2_dlygate4sd3_1 hold37 (.A(\adc_data0[3] ),
    .X(net141));
 sg13g2_dlygate4sd3_1 hold38 (.A(\adc_data2[8] ),
    .X(net142));
 sg13g2_dlygate4sd3_1 hold39 (.A(\adc_data2[6] ),
    .X(net143));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0054_),
    .X(net144));
 sg13g2_dlygate4sd3_1 hold41 (.A(\adc_data2[5] ),
    .X(net145));
 sg13g2_dlygate4sd3_1 hold42 (.A(\adc_data2[9] ),
    .X(net146));
 sg13g2_dlygate4sd3_1 hold43 (.A(\adc_data1[12] ),
    .X(net147));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0045_),
    .X(net148));
 sg13g2_dlygate4sd3_1 hold45 (.A(\adc_data2[3] ),
    .X(net149));
 sg13g2_dlygate4sd3_1 hold46 (.A(\adc_data0[8] ),
    .X(net150));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0026_),
    .X(net151));
 sg13g2_dlygate4sd3_1 hold48 (.A(\adc_data3[8] ),
    .X(net152));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0071_),
    .X(net153));
 sg13g2_dlygate4sd3_1 hold50 (.A(\adc_data3[5] ),
    .X(net154));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0068_),
    .X(net155));
 sg13g2_dlygate4sd3_1 hold52 (.A(\adc_data0[10] ),
    .X(net156));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0028_),
    .X(net157));
 sg13g2_dlygate4sd3_1 hold54 (.A(\adc_data3[12] ),
    .X(net158));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0075_),
    .X(net159));
 sg13g2_dlygate4sd3_1 hold56 (.A(\adc_data2[11] ),
    .X(net160));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0059_),
    .X(net161));
 sg13g2_dlygate4sd3_1 hold58 (.A(\adc_data1[8] ),
    .X(net162));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0041_),
    .X(net163));
 sg13g2_dlygate4sd3_1 hold60 (.A(\adc_data3[11] ),
    .X(net164));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0074_),
    .X(net165));
 sg13g2_dlygate4sd3_1 hold62 (.A(\adc_data1[4] ),
    .X(net166));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0037_),
    .X(net167));
 sg13g2_dlygate4sd3_1 hold64 (.A(\adc_data1[3] ),
    .X(net168));
 sg13g2_dlygate4sd3_1 hold65 (.A(\adc_data2[12] ),
    .X(net169));
 sg13g2_dlygate4sd3_1 hold66 (.A(\adc_data1[13] ),
    .X(net170));
 sg13g2_dlygate4sd3_1 hold67 (.A(\adc_data0[4] ),
    .X(net171));
 sg13g2_dlygate4sd3_1 hold68 (.A(\adc_data3[14] ),
    .X(net172));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0077_),
    .X(net173));
 sg13g2_dlygate4sd3_1 hold70 (.A(\adc_data3[9] ),
    .X(net174));
 sg13g2_dlygate4sd3_1 hold71 (.A(\clk_div[2] ),
    .X(net175));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0306_),
    .X(net176));
 sg13g2_dlygate4sd3_1 hold73 (.A(\adc_data3[3] ),
    .X(net177));
 sg13g2_dlygate4sd3_1 hold74 (.A(\adc_data2[13] ),
    .X(net178));
 sg13g2_dlygate4sd3_1 hold75 (.A(\adc_data2[10] ),
    .X(net179));
 sg13g2_dlygate4sd3_1 hold76 (.A(\adc_data3[13] ),
    .X(net180));
 sg13g2_dlygate4sd3_1 hold77 (.A(\adc_data2[14] ),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold78 (.A(\adc_data0[14] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold79 (.A(\adc_data1[10] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0043_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold81 (.A(\adc_data0[11] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold82 (.A(\adc_data1[7] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0040_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold84 (.A(\clk_div[3] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0308_),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold86 (.A(\adc_data0[7] ),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0025_),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold88 (.A(\adc_data0[1] ),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold89 (.A(\adc_data1[5] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold90 (.A(\clk_div[0] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold91 (.A(\adc_data0[12] ),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold92 (.A(\adc_data3[6] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold93 (.A(\adc_data1[6] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold94 (.A(\adc_data3[10] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold95 (.A(\clk_div[1] ),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold96 (.A(\cycle[3] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0257_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold98 (.A(\adc_data3[7] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold99 (.A(\adc_data0[9] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold100 (.A(\adc_data1[9] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold101 (.A(\adc_data3[4] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold102 (.A(\adc_data0[5] ),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold103 (.A(\cycle[2] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0255_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0002_),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold106 (.A(\adc_data1[11] ),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold107 (.A(\cycle[0] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold108 (.A(\adc_data1[14] ),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold109 (.A(\tx_cycle[0] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold110 (.A(\tx_cycle[6] ),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0297_),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold112 (.A(\adc_data0[6] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold113 (.A(\tx_cycle[5] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold114 (.A(\tx_cycle[1] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold115 (.A(\tx_cycle[4] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold116 (.A(\tx_cycle[2] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold117 (.A(\tx_cycle[3] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold118 (.A(adc_sclk),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0299_),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold120 (.A(adc_sclk),
    .X(net224));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_4 FILLER_5_231 ();
 sg13g2_fill_2 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_264 ();
 sg13g2_decap_8 FILLER_5_271 ();
 sg13g2_decap_8 FILLER_5_278 ();
 sg13g2_decap_8 FILLER_5_285 ();
 sg13g2_decap_8 FILLER_5_292 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_8 FILLER_5_306 ();
 sg13g2_decap_8 FILLER_5_313 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_4 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_197 ();
 sg13g2_decap_8 FILLER_6_204 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_240 ();
 sg13g2_decap_8 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_fill_1 FILLER_6_261 ();
 sg13g2_decap_8 FILLER_6_290 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_decap_8 FILLER_6_304 ();
 sg13g2_decap_8 FILLER_6_311 ();
 sg13g2_decap_8 FILLER_6_318 ();
 sg13g2_decap_8 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_332 ();
 sg13g2_decap_8 FILLER_6_339 ();
 sg13g2_decap_8 FILLER_6_346 ();
 sg13g2_decap_8 FILLER_6_353 ();
 sg13g2_decap_8 FILLER_6_360 ();
 sg13g2_decap_8 FILLER_6_367 ();
 sg13g2_decap_8 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_381 ();
 sg13g2_decap_8 FILLER_6_388 ();
 sg13g2_decap_8 FILLER_6_395 ();
 sg13g2_decap_8 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_8 FILLER_7_67 ();
 sg13g2_decap_8 FILLER_7_74 ();
 sg13g2_decap_8 FILLER_7_81 ();
 sg13g2_decap_8 FILLER_7_88 ();
 sg13g2_decap_8 FILLER_7_95 ();
 sg13g2_decap_8 FILLER_7_102 ();
 sg13g2_decap_8 FILLER_7_109 ();
 sg13g2_decap_8 FILLER_7_116 ();
 sg13g2_decap_8 FILLER_7_123 ();
 sg13g2_decap_8 FILLER_7_130 ();
 sg13g2_decap_8 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_151 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_4 FILLER_7_165 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_decap_8 FILLER_7_174 ();
 sg13g2_decap_8 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_229 ();
 sg13g2_decap_4 FILLER_7_235 ();
 sg13g2_decap_4 FILLER_7_246 ();
 sg13g2_decap_4 FILLER_7_272 ();
 sg13g2_decap_4 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_316 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_4 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_36 ();
 sg13g2_fill_2 FILLER_8_43 ();
 sg13g2_fill_1 FILLER_8_45 ();
 sg13g2_decap_8 FILLER_8_78 ();
 sg13g2_decap_8 FILLER_8_85 ();
 sg13g2_decap_8 FILLER_8_92 ();
 sg13g2_decap_4 FILLER_8_99 ();
 sg13g2_decap_8 FILLER_8_107 ();
 sg13g2_decap_8 FILLER_8_114 ();
 sg13g2_decap_8 FILLER_8_121 ();
 sg13g2_decap_8 FILLER_8_128 ();
 sg13g2_decap_8 FILLER_8_135 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_fill_1 FILLER_8_202 ();
 sg13g2_fill_2 FILLER_8_224 ();
 sg13g2_decap_4 FILLER_8_256 ();
 sg13g2_fill_1 FILLER_8_260 ();
 sg13g2_decap_8 FILLER_8_285 ();
 sg13g2_fill_1 FILLER_8_292 ();
 sg13g2_fill_2 FILLER_8_306 ();
 sg13g2_fill_1 FILLER_8_308 ();
 sg13g2_fill_2 FILLER_8_318 ();
 sg13g2_fill_1 FILLER_8_320 ();
 sg13g2_decap_8 FILLER_8_330 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_351 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_decap_8 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_372 ();
 sg13g2_decap_8 FILLER_8_379 ();
 sg13g2_decap_8 FILLER_8_386 ();
 sg13g2_decap_8 FILLER_8_393 ();
 sg13g2_decap_8 FILLER_8_400 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_fill_2 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_54 ();
 sg13g2_decap_8 FILLER_9_61 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_153 ();
 sg13g2_decap_4 FILLER_9_160 ();
 sg13g2_fill_2 FILLER_9_181 ();
 sg13g2_fill_1 FILLER_9_191 ();
 sg13g2_fill_1 FILLER_9_251 ();
 sg13g2_decap_4 FILLER_9_270 ();
 sg13g2_fill_2 FILLER_9_274 ();
 sg13g2_decap_8 FILLER_9_337 ();
 sg13g2_decap_8 FILLER_9_344 ();
 sg13g2_decap_8 FILLER_9_351 ();
 sg13g2_decap_8 FILLER_9_358 ();
 sg13g2_decap_8 FILLER_9_365 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_decap_4 FILLER_10_10 ();
 sg13g2_fill_1 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_49 ();
 sg13g2_fill_2 FILLER_10_58 ();
 sg13g2_fill_1 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_163 ();
 sg13g2_fill_2 FILLER_10_175 ();
 sg13g2_fill_2 FILLER_10_203 ();
 sg13g2_fill_2 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_225 ();
 sg13g2_decap_4 FILLER_10_242 ();
 sg13g2_fill_1 FILLER_10_246 ();
 sg13g2_fill_2 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_254 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_fill_2 FILLER_10_283 ();
 sg13g2_fill_1 FILLER_10_285 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_59 ();
 sg13g2_fill_2 FILLER_11_66 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_130 ();
 sg13g2_fill_1 FILLER_11_132 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_fill_2 FILLER_11_165 ();
 sg13g2_decap_4 FILLER_11_179 ();
 sg13g2_fill_1 FILLER_11_183 ();
 sg13g2_fill_2 FILLER_11_197 ();
 sg13g2_fill_1 FILLER_11_199 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_fill_2 FILLER_11_234 ();
 sg13g2_decap_8 FILLER_11_241 ();
 sg13g2_fill_1 FILLER_11_248 ();
 sg13g2_fill_2 FILLER_11_293 ();
 sg13g2_fill_2 FILLER_11_309 ();
 sg13g2_fill_1 FILLER_11_338 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_fill_2 FILLER_12_10 ();
 sg13g2_fill_2 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_fill_2 FILLER_12_118 ();
 sg13g2_fill_1 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_154 ();
 sg13g2_fill_1 FILLER_12_184 ();
 sg13g2_decap_4 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_209 ();
 sg13g2_fill_1 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_227 ();
 sg13g2_decap_4 FILLER_12_259 ();
 sg13g2_decap_4 FILLER_12_306 ();
 sg13g2_fill_2 FILLER_12_331 ();
 sg13g2_fill_1 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_fill_2 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_386 ();
 sg13g2_decap_8 FILLER_12_393 ();
 sg13g2_decap_8 FILLER_12_400 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_33 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_fill_2 FILLER_13_63 ();
 sg13g2_fill_1 FILLER_13_65 ();
 sg13g2_decap_4 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_124 ();
 sg13g2_fill_2 FILLER_13_144 ();
 sg13g2_fill_1 FILLER_13_146 ();
 sg13g2_decap_4 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_4 FILLER_13_200 ();
 sg13g2_fill_2 FILLER_13_204 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_decap_4 FILLER_13_250 ();
 sg13g2_fill_2 FILLER_13_263 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_4 FILLER_13_321 ();
 sg13g2_decap_8 FILLER_13_330 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_fill_1 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_37 ();
 sg13g2_fill_1 FILLER_14_39 ();
 sg13g2_fill_2 FILLER_14_45 ();
 sg13g2_fill_1 FILLER_14_47 ();
 sg13g2_decap_4 FILLER_14_57 ();
 sg13g2_fill_2 FILLER_14_61 ();
 sg13g2_decap_8 FILLER_14_80 ();
 sg13g2_decap_4 FILLER_14_87 ();
 sg13g2_fill_1 FILLER_14_91 ();
 sg13g2_fill_2 FILLER_14_108 ();
 sg13g2_fill_1 FILLER_14_110 ();
 sg13g2_fill_2 FILLER_14_147 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_decap_8 FILLER_14_163 ();
 sg13g2_decap_4 FILLER_14_195 ();
 sg13g2_fill_2 FILLER_14_199 ();
 sg13g2_fill_1 FILLER_14_215 ();
 sg13g2_fill_2 FILLER_14_221 ();
 sg13g2_fill_1 FILLER_14_223 ();
 sg13g2_fill_2 FILLER_14_233 ();
 sg13g2_decap_4 FILLER_14_244 ();
 sg13g2_fill_2 FILLER_14_248 ();
 sg13g2_fill_1 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_fill_2 FILLER_14_291 ();
 sg13g2_fill_1 FILLER_14_293 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_341 ();
 sg13g2_fill_2 FILLER_14_349 ();
 sg13g2_fill_2 FILLER_14_379 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_29 ();
 sg13g2_fill_2 FILLER_15_45 ();
 sg13g2_fill_1 FILLER_15_47 ();
 sg13g2_fill_2 FILLER_15_58 ();
 sg13g2_fill_1 FILLER_15_60 ();
 sg13g2_fill_1 FILLER_15_71 ();
 sg13g2_decap_4 FILLER_15_77 ();
 sg13g2_fill_2 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_fill_2 FILLER_15_132 ();
 sg13g2_fill_2 FILLER_15_138 ();
 sg13g2_decap_4 FILLER_15_179 ();
 sg13g2_fill_2 FILLER_15_183 ();
 sg13g2_decap_4 FILLER_15_198 ();
 sg13g2_fill_2 FILLER_15_222 ();
 sg13g2_fill_2 FILLER_15_255 ();
 sg13g2_fill_2 FILLER_15_283 ();
 sg13g2_fill_2 FILLER_15_306 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_fill_1 FILLER_15_346 ();
 sg13g2_fill_2 FILLER_15_365 ();
 sg13g2_fill_1 FILLER_15_367 ();
 sg13g2_fill_2 FILLER_15_386 ();
 sg13g2_decap_4 FILLER_15_405 ();
 sg13g2_decap_4 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_10 ();
 sg13g2_decap_8 FILLER_16_17 ();
 sg13g2_fill_1 FILLER_16_24 ();
 sg13g2_fill_1 FILLER_16_39 ();
 sg13g2_fill_1 FILLER_16_45 ();
 sg13g2_fill_2 FILLER_16_56 ();
 sg13g2_fill_1 FILLER_16_58 ();
 sg13g2_fill_1 FILLER_16_79 ();
 sg13g2_fill_1 FILLER_16_91 ();
 sg13g2_decap_4 FILLER_16_97 ();
 sg13g2_fill_2 FILLER_16_101 ();
 sg13g2_fill_2 FILLER_16_134 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_fill_2 FILLER_16_211 ();
 sg13g2_decap_4 FILLER_16_217 ();
 sg13g2_fill_2 FILLER_16_221 ();
 sg13g2_decap_4 FILLER_16_232 ();
 sg13g2_decap_4 FILLER_16_242 ();
 sg13g2_fill_2 FILLER_16_246 ();
 sg13g2_fill_2 FILLER_16_289 ();
 sg13g2_fill_1 FILLER_16_301 ();
 sg13g2_fill_1 FILLER_16_323 ();
 sg13g2_fill_1 FILLER_16_336 ();
 sg13g2_fill_2 FILLER_16_346 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_2 FILLER_16_379 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_decap_4 FILLER_17_63 ();
 sg13g2_fill_1 FILLER_17_67 ();
 sg13g2_fill_2 FILLER_17_89 ();
 sg13g2_fill_1 FILLER_17_91 ();
 sg13g2_decap_4 FILLER_17_111 ();
 sg13g2_fill_1 FILLER_17_162 ();
 sg13g2_fill_2 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_171 ();
 sg13g2_fill_1 FILLER_17_185 ();
 sg13g2_decap_8 FILLER_17_199 ();
 sg13g2_decap_4 FILLER_17_206 ();
 sg13g2_fill_2 FILLER_17_210 ();
 sg13g2_decap_4 FILLER_17_216 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_fill_2 FILLER_17_284 ();
 sg13g2_fill_2 FILLER_17_296 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_4 FILLER_17_315 ();
 sg13g2_fill_1 FILLER_17_319 ();
 sg13g2_decap_4 FILLER_17_325 ();
 sg13g2_decap_4 FILLER_17_366 ();
 sg13g2_decap_8 FILLER_17_401 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_10 ();
 sg13g2_fill_2 FILLER_18_17 ();
 sg13g2_fill_1 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_161 ();
 sg13g2_decap_4 FILLER_18_193 ();
 sg13g2_fill_1 FILLER_18_197 ();
 sg13g2_fill_1 FILLER_18_273 ();
 sg13g2_fill_1 FILLER_18_278 ();
 sg13g2_fill_2 FILLER_18_284 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_decap_4 FILLER_18_307 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_360 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_45 ();
 sg13g2_fill_1 FILLER_19_47 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_87 ();
 sg13g2_decap_8 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_108 ();
 sg13g2_fill_1 FILLER_19_171 ();
 sg13g2_decap_8 FILLER_19_208 ();
 sg13g2_decap_8 FILLER_19_215 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_4 FILLER_19_242 ();
 sg13g2_fill_2 FILLER_19_246 ();
 sg13g2_decap_8 FILLER_19_261 ();
 sg13g2_fill_2 FILLER_19_268 ();
 sg13g2_fill_1 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_decap_4 FILLER_19_329 ();
 sg13g2_fill_2 FILLER_19_364 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_fill_2 FILLER_20_18 ();
 sg13g2_fill_2 FILLER_20_56 ();
 sg13g2_fill_1 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_85 ();
 sg13g2_decap_8 FILLER_20_92 ();
 sg13g2_fill_2 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_fill_1 FILLER_20_152 ();
 sg13g2_fill_1 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_195 ();
 sg13g2_fill_2 FILLER_20_200 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_234 ();
 sg13g2_fill_1 FILLER_20_236 ();
 sg13g2_fill_1 FILLER_20_277 ();
 sg13g2_fill_1 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_4 FILLER_20_357 ();
 sg13g2_fill_2 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_366 ();
 sg13g2_fill_1 FILLER_20_377 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_29 ();
 sg13g2_fill_1 FILLER_21_31 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_51 ();
 sg13g2_decap_8 FILLER_21_55 ();
 sg13g2_decap_8 FILLER_21_62 ();
 sg13g2_fill_1 FILLER_21_69 ();
 sg13g2_decap_4 FILLER_21_90 ();
 sg13g2_fill_2 FILLER_21_94 ();
 sg13g2_fill_1 FILLER_21_108 ();
 sg13g2_fill_2 FILLER_21_122 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_decap_8 FILLER_21_239 ();
 sg13g2_decap_4 FILLER_21_246 ();
 sg13g2_fill_1 FILLER_21_250 ();
 sg13g2_decap_4 FILLER_21_268 ();
 sg13g2_fill_2 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_4 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_fill_2 FILLER_21_336 ();
 sg13g2_fill_1 FILLER_21_338 ();
 sg13g2_decap_4 FILLER_21_369 ();
 sg13g2_fill_2 FILLER_21_373 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_4 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_65 ();
 sg13g2_decap_8 FILLER_22_72 ();
 sg13g2_decap_4 FILLER_22_79 ();
 sg13g2_fill_2 FILLER_22_115 ();
 sg13g2_fill_1 FILLER_22_136 ();
 sg13g2_fill_1 FILLER_22_226 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_300 ();
 sg13g2_decap_4 FILLER_22_314 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_4 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_352 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_fill_1 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_fill_1 FILLER_23_16 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_decap_4 FILLER_23_43 ();
 sg13g2_fill_1 FILLER_23_47 ();
 sg13g2_decap_4 FILLER_23_92 ();
 sg13g2_fill_2 FILLER_23_128 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_fill_1 FILLER_23_165 ();
 sg13g2_fill_2 FILLER_23_192 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_1 FILLER_23_246 ();
 sg13g2_fill_2 FILLER_23_260 ();
 sg13g2_fill_2 FILLER_23_275 ();
 sg13g2_fill_2 FILLER_23_290 ();
 sg13g2_fill_1 FILLER_23_292 ();
 sg13g2_fill_2 FILLER_23_312 ();
 sg13g2_decap_4 FILLER_23_357 ();
 sg13g2_fill_1 FILLER_23_361 ();
 sg13g2_fill_2 FILLER_23_380 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_11 ();
 sg13g2_decap_4 FILLER_24_66 ();
 sg13g2_decap_4 FILLER_24_79 ();
 sg13g2_decap_4 FILLER_24_96 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_2 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_fill_2 FILLER_24_193 ();
 sg13g2_decap_4 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_231 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_decap_8 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_decap_4 FILLER_24_304 ();
 sg13g2_decap_4 FILLER_24_311 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_330 ();
 sg13g2_fill_1 FILLER_24_332 ();
 sg13g2_decap_4 FILLER_24_344 ();
 sg13g2_fill_1 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_29 ();
 sg13g2_fill_2 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_fill_1 FILLER_25_105 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_167 ();
 sg13g2_fill_1 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_decap_4 FILLER_25_211 ();
 sg13g2_fill_1 FILLER_25_215 ();
 sg13g2_fill_1 FILLER_25_221 ();
 sg13g2_fill_1 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_fill_2 FILLER_25_272 ();
 sg13g2_fill_1 FILLER_25_293 ();
 sg13g2_decap_4 FILLER_25_324 ();
 sg13g2_fill_2 FILLER_25_328 ();
 sg13g2_decap_4 FILLER_25_350 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_fill_2 FILLER_26_10 ();
 sg13g2_decap_8 FILLER_26_89 ();
 sg13g2_decap_4 FILLER_26_96 ();
 sg13g2_fill_1 FILLER_26_100 ();
 sg13g2_decap_4 FILLER_26_111 ();
 sg13g2_fill_1 FILLER_26_115 ();
 sg13g2_fill_2 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_183 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_4 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_250 ();
 sg13g2_fill_2 FILLER_26_269 ();
 sg13g2_decap_4 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_294 ();
 sg13g2_fill_1 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_302 ();
 sg13g2_fill_2 FILLER_26_308 ();
 sg13g2_fill_2 FILLER_26_328 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_decap_4 FILLER_26_392 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_4 ();
 sg13g2_decap_4 FILLER_27_10 ();
 sg13g2_fill_2 FILLER_27_30 ();
 sg13g2_fill_1 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_96 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_fill_2 FILLER_27_119 ();
 sg13g2_decap_4 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_155 ();
 sg13g2_fill_1 FILLER_27_160 ();
 sg13g2_fill_2 FILLER_27_169 ();
 sg13g2_fill_1 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_209 ();
 sg13g2_decap_8 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_223 ();
 sg13g2_fill_2 FILLER_27_243 ();
 sg13g2_decap_8 FILLER_27_264 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_fill_2 FILLER_27_293 ();
 sg13g2_fill_1 FILLER_27_295 ();
 sg13g2_fill_1 FILLER_27_305 ();
 sg13g2_fill_1 FILLER_27_319 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_fill_1 FILLER_27_379 ();
 sg13g2_decap_4 FILLER_27_393 ();
 sg13g2_fill_1 FILLER_27_397 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_29 ();
 sg13g2_fill_2 FILLER_28_44 ();
 sg13g2_fill_1 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_95 ();
 sg13g2_decap_4 FILLER_28_103 ();
 sg13g2_fill_1 FILLER_28_107 ();
 sg13g2_decap_8 FILLER_28_129 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_184 ();
 sg13g2_decap_8 FILLER_28_235 ();
 sg13g2_decap_4 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_288 ();
 sg13g2_fill_1 FILLER_28_337 ();
 sg13g2_fill_2 FILLER_28_359 ();
 sg13g2_decap_4 FILLER_28_390 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_14 ();
 sg13g2_decap_4 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_53 ();
 sg13g2_fill_1 FILLER_29_59 ();
 sg13g2_decap_4 FILLER_29_65 ();
 sg13g2_fill_2 FILLER_29_69 ();
 sg13g2_decap_8 FILLER_29_94 ();
 sg13g2_decap_8 FILLER_29_115 ();
 sg13g2_decap_8 FILLER_29_122 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_fill_1 FILLER_29_131 ();
 sg13g2_decap_4 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_200 ();
 sg13g2_fill_1 FILLER_29_202 ();
 sg13g2_fill_2 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_decap_8 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_322 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_decap_4 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_60 ();
 sg13g2_fill_1 FILLER_30_62 ();
 sg13g2_decap_4 FILLER_30_80 ();
 sg13g2_fill_1 FILLER_30_84 ();
 sg13g2_decap_4 FILLER_30_150 ();
 sg13g2_fill_2 FILLER_30_159 ();
 sg13g2_fill_1 FILLER_30_161 ();
 sg13g2_decap_4 FILLER_30_171 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_decap_4 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_215 ();
 sg13g2_decap_4 FILLER_30_221 ();
 sg13g2_decap_4 FILLER_30_241 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_fill_1 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_fill_1 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_313 ();
 sg13g2_fill_2 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_decap_8 FILLER_30_397 ();
 sg13g2_decap_4 FILLER_30_404 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_4 ();
 sg13g2_fill_2 FILLER_31_26 ();
 sg13g2_decap_4 FILLER_31_49 ();
 sg13g2_fill_1 FILLER_31_53 ();
 sg13g2_fill_1 FILLER_31_63 ();
 sg13g2_fill_2 FILLER_31_69 ();
 sg13g2_decap_4 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_105 ();
 sg13g2_decap_4 FILLER_31_118 ();
 sg13g2_fill_1 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_166 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_180 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_4 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_fill_2 FILLER_31_238 ();
 sg13g2_fill_2 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_266 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_375 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_55 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_108 ();
 sg13g2_decap_8 FILLER_32_115 ();
 sg13g2_decap_4 FILLER_32_148 ();
 sg13g2_fill_1 FILLER_32_180 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_215 ();
 sg13g2_decap_4 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_265 ();
 sg13g2_decap_8 FILLER_32_272 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_4 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_329 ();
 sg13g2_decap_4 FILLER_32_346 ();
 sg13g2_fill_2 FILLER_32_350 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_10 ();
 sg13g2_fill_1 FILLER_33_17 ();
 sg13g2_decap_8 FILLER_33_47 ();
 sg13g2_decap_8 FILLER_33_54 ();
 sg13g2_decap_4 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_65 ();
 sg13g2_decap_4 FILLER_33_82 ();
 sg13g2_decap_4 FILLER_33_95 ();
 sg13g2_decap_4 FILLER_33_110 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_fill_1 FILLER_33_145 ();
 sg13g2_fill_1 FILLER_33_169 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_fill_2 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_4 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_4 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_290 ();
 sg13g2_decap_8 FILLER_33_312 ();
 sg13g2_decap_8 FILLER_33_319 ();
 sg13g2_decap_8 FILLER_33_337 ();
 sg13g2_fill_2 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_32 ();
 sg13g2_fill_2 FILLER_34_51 ();
 sg13g2_fill_1 FILLER_34_53 ();
 sg13g2_fill_2 FILLER_34_67 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_1 FILLER_34_93 ();
 sg13g2_fill_2 FILLER_34_104 ();
 sg13g2_fill_2 FILLER_34_127 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_175 ();
 sg13g2_fill_1 FILLER_34_182 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_238 ();
 sg13g2_fill_1 FILLER_34_245 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_decap_8 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_280 ();
 sg13g2_fill_2 FILLER_34_294 ();
 sg13g2_decap_8 FILLER_34_304 ();
 sg13g2_decap_4 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_341 ();
 sg13g2_fill_2 FILLER_34_351 ();
 sg13g2_fill_1 FILLER_34_366 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_13 ();
 sg13g2_decap_4 FILLER_35_20 ();
 sg13g2_fill_2 FILLER_35_24 ();
 sg13g2_fill_2 FILLER_35_42 ();
 sg13g2_fill_1 FILLER_35_44 ();
 sg13g2_decap_4 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_89 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_156 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_fill_1 FILLER_35_174 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_fill_1 FILLER_35_181 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_fill_1 FILLER_35_241 ();
 sg13g2_decap_4 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_263 ();
 sg13g2_decap_8 FILLER_35_267 ();
 sg13g2_decap_8 FILLER_35_274 ();
 sg13g2_decap_4 FILLER_35_281 ();
 sg13g2_fill_2 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_334 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_fill_1 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_decap_4 FILLER_36_74 ();
 sg13g2_fill_2 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_89 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_decap_4 FILLER_36_103 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_135 ();
 sg13g2_fill_2 FILLER_36_164 ();
 sg13g2_fill_1 FILLER_36_166 ();
 sg13g2_fill_2 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_206 ();
 sg13g2_fill_1 FILLER_36_217 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_254 ();
 sg13g2_fill_2 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_263 ();
 sg13g2_decap_4 FILLER_36_280 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_fill_2 FILLER_36_304 ();
 sg13g2_fill_2 FILLER_36_333 ();
 sg13g2_fill_1 FILLER_36_339 ();
 sg13g2_fill_2 FILLER_36_391 ();
 sg13g2_fill_1 FILLER_36_393 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_14 ();
 sg13g2_decap_4 FILLER_37_32 ();
 sg13g2_fill_1 FILLER_37_36 ();
 sg13g2_decap_8 FILLER_37_128 ();
 sg13g2_decap_4 FILLER_37_135 ();
 sg13g2_fill_2 FILLER_37_139 ();
 sg13g2_decap_8 FILLER_37_145 ();
 sg13g2_decap_8 FILLER_37_152 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_decap_4 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_170 ();
 sg13g2_fill_1 FILLER_37_176 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_188 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_decap_4 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_243 ();
 sg13g2_decap_4 FILLER_37_259 ();
 sg13g2_fill_1 FILLER_37_294 ();
 sg13g2_fill_2 FILLER_37_315 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_4 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_18 ();
 sg13g2_decap_8 FILLER_38_32 ();
 sg13g2_decap_8 FILLER_38_39 ();
 sg13g2_fill_2 FILLER_38_46 ();
 sg13g2_fill_1 FILLER_38_48 ();
 sg13g2_fill_2 FILLER_38_53 ();
 sg13g2_fill_1 FILLER_38_55 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_116 ();
 sg13g2_fill_1 FILLER_38_118 ();
 sg13g2_decap_8 FILLER_38_127 ();
 sg13g2_decap_8 FILLER_38_134 ();
 sg13g2_decap_8 FILLER_38_141 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_273 ();
 sg13g2_fill_1 FILLER_38_275 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_fill_1 FILLER_38_324 ();
 sg13g2_fill_2 FILLER_38_362 ();
 sg13g2_fill_1 FILLER_38_364 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net10;
 assign uio_oe[1] = net11;
 assign uio_oe[2] = net12;
 assign uio_oe[3] = net13;
 assign uio_oe[4] = net102;
 assign uio_oe[5] = net103;
 assign uio_oe[6] = net104;
 assign uio_oe[7] = net14;
 assign uio_out[0] = net15;
 assign uio_out[1] = net16;
 assign uio_out[2] = net17;
 assign uio_out[3] = net18;
 assign uio_out[7] = net19;
endmodule
