module tt_um_urish_rings (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire clknet_0_clk;
 wire \abs_x[0] ;
 wire \abs_y[0] ;
 wire \anim_offset[1] ;
 wire \anim_offset[2] ;
 wire \anim_offset[3] ;
 wire \anim_offset[4] ;
 wire \anim_offset[5] ;
 wire \anim_offset[6] ;
 wire \anim_offset[7] ;
 wire \cx[1] ;
 wire \cx[2] ;
 wire \cx[3] ;
 wire \cx[4] ;
 wire \cx[5] ;
 wire \cy[1] ;
 wire \cy[2] ;
 wire \cy[3] ;
 wire \hpos[6] ;
 wire \hpos[7] ;
 wire \hpos[8] ;
 wire \hpos[9] ;
 wire hsync;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net1;
 wire net2;
 wire net3;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sg13g2_inv_1 _326_ (.Y(_270_),
    .A(net39));
 sg13g2_inv_2 _327_ (.Y(_271_),
    .A(net80));
 sg13g2_inv_1 _328_ (.Y(_272_),
    .A(net42));
 sg13g2_inv_2 _329_ (.Y(_273_),
    .A(net40));
 sg13g2_inv_1 _330_ (.Y(_274_),
    .A(net91));
 sg13g2_inv_1 _331_ (.Y(_275_),
    .A(net70));
 sg13g2_inv_2 _332_ (.Y(_276_),
    .A(net74));
 sg13g2_inv_1 _333_ (.Y(_277_),
    .A(net2));
 sg13g2_inv_2 _334_ (.Y(_278_),
    .A(net77));
 sg13g2_and4_1 _335_ (.A(net36),
    .B(net78),
    .C(net76),
    .D(net68),
    .X(_279_));
 sg13g2_nand2_2 _336_ (.Y(_280_),
    .A(net70),
    .B(net72));
 sg13g2_nor4_1 _337_ (.A(_274_),
    .B(_275_),
    .C(net38),
    .D(net79),
    .Y(_281_));
 sg13g2_nand3_1 _338_ (.B(_280_),
    .C(_281_),
    .A(_279_),
    .Y(_001_));
 sg13g2_nor2_1 _339_ (.A(net80),
    .B(net83),
    .Y(_282_));
 sg13g2_nand4_1 _340_ (.B(net83),
    .C(net41),
    .A(net80),
    .Y(_283_),
    .D(net42));
 sg13g2_a21oi_1 _341_ (.A1(_272_),
    .A2(_282_),
    .Y(_284_),
    .B1(net85));
 sg13g2_nand4_1 _342_ (.B(net40),
    .C(_283_),
    .A(net41),
    .Y(_000_),
    .D(_284_));
 sg13g2_nand2_1 _343_ (.Y(_285_),
    .A(net36),
    .B(net37));
 sg13g2_and4_1 _344_ (.A(net36),
    .B(net37),
    .C(\hvsync_gen.vpos[7] ),
    .D(\hvsync_gen.vpos[6] ),
    .X(_286_));
 sg13g2_nand4_1 _345_ (.B(net37),
    .C(\hvsync_gen.vpos[7] ),
    .A(net36),
    .Y(_287_),
    .D(\hvsync_gen.vpos[6] ));
 sg13g2_nor2_1 _346_ (.A(\hvsync_gen.vpos[8] ),
    .B(\hvsync_gen.vpos[9] ),
    .Y(_288_));
 sg13g2_or2_1 _347_ (.X(_289_),
    .B(\hvsync_gen.vpos[9] ),
    .A(\hvsync_gen.vpos[8] ));
 sg13g2_or2_1 _348_ (.X(_290_),
    .B(\cy[1] ),
    .A(net39));
 sg13g2_nor3_1 _349_ (.A(net39),
    .B(\cy[1] ),
    .C(\cy[2] ),
    .Y(_291_));
 sg13g2_nor4_1 _350_ (.A(net39),
    .B(\cy[1] ),
    .C(\cy[3] ),
    .D(\cy[2] ),
    .Y(_292_));
 sg13g2_nor3_2 _351_ (.A(_286_),
    .B(_289_),
    .C(_292_),
    .Y(_293_));
 sg13g2_xnor2_1 _352_ (.Y(_294_),
    .A(net38),
    .B(_293_));
 sg13g2_nor2_1 _353_ (.A(net41),
    .B(net42),
    .Y(_295_));
 sg13g2_nor2b_1 _354_ (.A(_295_),
    .B_N(\hpos[8] ),
    .Y(_296_));
 sg13g2_o21ai_1 _355_ (.B1(\hpos[8] ),
    .Y(_297_),
    .A1(net41),
    .A2(net42));
 sg13g2_nand2_1 _356_ (.Y(_298_),
    .A(_273_),
    .B(_297_));
 sg13g2_or2_1 _357_ (.X(_299_),
    .B(\cx[1] ),
    .A(\abs_x[0] ));
 sg13g2_or3_1 _358_ (.A(net43),
    .B(\cx[1] ),
    .C(\cx[2] ),
    .X(_300_));
 sg13g2_nor4_1 _359_ (.A(net43),
    .B(\cx[1] ),
    .C(\cx[2] ),
    .D(\cx[3] ),
    .Y(_301_));
 sg13g2_or4_1 _360_ (.A(net43),
    .B(\cx[1] ),
    .C(\cx[2] ),
    .D(\cx[3] ),
    .X(_302_));
 sg13g2_nand2_2 _361_ (.Y(_303_),
    .A(_282_),
    .B(_301_));
 sg13g2_nor2b_1 _362_ (.A(_298_),
    .B_N(_303_),
    .Y(_029_));
 sg13g2_xnor2_1 _363_ (.Y(_030_),
    .A(net42),
    .B(_029_));
 sg13g2_xnor2_1 _364_ (.Y(_031_),
    .A(_272_),
    .B(_029_));
 sg13g2_a21o_2 _365_ (.A2(_288_),
    .A1(_285_),
    .B1(_293_),
    .X(_032_));
 sg13g2_and3_1 _366_ (.X(_033_),
    .A(net36),
    .B(net37),
    .C(\hvsync_gen.vpos[6] ));
 sg13g2_xor2_1 _367_ (.B(_285_),
    .A(\hvsync_gen.vpos[6] ),
    .X(_034_));
 sg13g2_nor2_1 _368_ (.A(_289_),
    .B(_033_),
    .Y(_035_));
 sg13g2_nor2_1 _369_ (.A(_293_),
    .B(_035_),
    .Y(_036_));
 sg13g2_xnor2_1 _370_ (.Y(_037_),
    .A(_032_),
    .B(_034_));
 sg13g2_inv_1 _371_ (.Y(_038_),
    .A(_037_));
 sg13g2_xor2_1 _372_ (.B(net38),
    .A(net36),
    .X(_039_));
 sg13g2_inv_1 _373_ (.Y(_040_),
    .A(_039_));
 sg13g2_o21ai_1 _374_ (.B1(_039_),
    .Y(_041_),
    .A1(net38),
    .A2(_289_));
 sg13g2_nor2_1 _375_ (.A(_293_),
    .B(_041_),
    .Y(_042_));
 sg13g2_a21oi_2 _376_ (.B1(_042_),
    .Y(_043_),
    .A2(_040_),
    .A1(_032_));
 sg13g2_a21o_1 _377_ (.A2(_040_),
    .A1(_032_),
    .B1(_042_),
    .X(_044_));
 sg13g2_nand3_1 _378_ (.B(_297_),
    .C(_302_),
    .A(_273_),
    .Y(_045_));
 sg13g2_a21oi_1 _379_ (.A1(_271_),
    .A2(_301_),
    .Y(_046_),
    .B1(_298_));
 sg13g2_xor2_1 _380_ (.B(_046_),
    .A(\cx[5] ),
    .X(_047_));
 sg13g2_xnor2_1 _381_ (.Y(_048_),
    .A(\cx[5] ),
    .B(_046_));
 sg13g2_a22oi_1 _382_ (.Y(_049_),
    .B1(_044_),
    .B2(_048_),
    .A2(_037_),
    .A1(_031_));
 sg13g2_xnor2_1 _383_ (.Y(_050_),
    .A(_271_),
    .B(_045_));
 sg13g2_nor2_1 _384_ (.A(_294_),
    .B(_050_),
    .Y(_051_));
 sg13g2_a21oi_1 _385_ (.A1(_043_),
    .A2(_047_),
    .Y(_052_),
    .B1(_051_));
 sg13g2_a21o_1 _386_ (.A2(_047_),
    .A1(_043_),
    .B1(_051_),
    .X(_053_));
 sg13g2_xnor2_1 _387_ (.Y(_054_),
    .A(net41),
    .B(\hpos[6] ));
 sg13g2_nand3_1 _388_ (.B(_282_),
    .C(_301_),
    .A(\hpos[6] ),
    .Y(_055_));
 sg13g2_nor2b_1 _389_ (.A(_298_),
    .B_N(_055_),
    .Y(_056_));
 sg13g2_xnor2_1 _390_ (.Y(_057_),
    .A(_054_),
    .B(_056_));
 sg13g2_o21ai_1 _391_ (.B1(_287_),
    .Y(_058_),
    .A1(\hvsync_gen.vpos[7] ),
    .A2(_033_));
 sg13g2_xor2_1 _392_ (.B(_058_),
    .A(_036_),
    .X(_059_));
 sg13g2_nor2_1 _393_ (.A(_057_),
    .B(_059_),
    .Y(_060_));
 sg13g2_a221oi_1 _394_ (.B2(_053_),
    .C1(_060_),
    .B1(_049_),
    .A1(_030_),
    .Y(_061_),
    .A2(_038_));
 sg13g2_nand3_1 _395_ (.B(_288_),
    .C(_290_),
    .A(_287_),
    .Y(_062_));
 sg13g2_xnor2_1 _396_ (.Y(_063_),
    .A(\cy[2] ),
    .B(_062_));
 sg13g2_nand3_1 _397_ (.B(_297_),
    .C(_299_),
    .A(_273_),
    .Y(_064_));
 sg13g2_xor2_1 _398_ (.B(_064_),
    .A(\cx[2] ),
    .X(_065_));
 sg13g2_nand2b_1 _399_ (.Y(_066_),
    .B(net39),
    .A_N(\abs_x[0] ));
 sg13g2_xnor2_1 _400_ (.Y(_067_),
    .A(net43),
    .B(net98));
 sg13g2_nand3_1 _401_ (.B(_297_),
    .C(_067_),
    .A(_273_),
    .Y(_068_));
 sg13g2_a21o_1 _402_ (.A2(_297_),
    .A1(_273_),
    .B1(\cx[1] ),
    .X(_069_));
 sg13g2_and2_1 _403_ (.A(_068_),
    .B(_069_),
    .X(_070_));
 sg13g2_nand3_1 _404_ (.B(_068_),
    .C(_069_),
    .A(_066_),
    .Y(_071_));
 sg13g2_nand2_1 _405_ (.Y(_072_),
    .A(net39),
    .B(net91));
 sg13g2_xor2_1 _406_ (.B(net91),
    .A(net39),
    .X(_073_));
 sg13g2_nor3_1 _407_ (.A(_286_),
    .B(_289_),
    .C(_073_),
    .Y(_074_));
 sg13g2_a21oi_1 _408_ (.A1(_287_),
    .A2(_288_),
    .Y(_075_),
    .B1(\cy[1] ));
 sg13g2_nor2_1 _409_ (.A(_074_),
    .B(_075_),
    .Y(_076_));
 sg13g2_or2_1 _410_ (.X(_077_),
    .B(_299_),
    .A(_270_));
 sg13g2_o21ai_1 _411_ (.B1(_077_),
    .Y(_078_),
    .A1(_074_),
    .A2(_075_));
 sg13g2_a22oi_1 _412_ (.Y(_079_),
    .B1(_071_),
    .B2(_078_),
    .A2(_065_),
    .A1(_063_));
 sg13g2_nor2_1 _413_ (.A(_063_),
    .B(_065_),
    .Y(_080_));
 sg13g2_nand3_1 _414_ (.B(_297_),
    .C(_300_),
    .A(_273_),
    .Y(_081_));
 sg13g2_xor2_1 _415_ (.B(_081_),
    .A(\cx[3] ),
    .X(_082_));
 sg13g2_nor3_1 _416_ (.A(_286_),
    .B(_289_),
    .C(_291_),
    .Y(_083_));
 sg13g2_xnor2_1 _417_ (.Y(_084_),
    .A(\cy[3] ),
    .B(_083_));
 sg13g2_nor2b_1 _418_ (.A(_082_),
    .B_N(_084_),
    .Y(_085_));
 sg13g2_or3_1 _419_ (.A(_079_),
    .B(_080_),
    .C(_085_),
    .X(_086_));
 sg13g2_nor2b_1 _420_ (.A(_084_),
    .B_N(_082_),
    .Y(_087_));
 sg13g2_a21oi_1 _421_ (.A1(_294_),
    .A2(_050_),
    .Y(_088_),
    .B1(_087_));
 sg13g2_nand4_1 _422_ (.B(_052_),
    .C(_086_),
    .A(_049_),
    .Y(_089_),
    .D(_088_));
 sg13g2_nor3_1 _423_ (.A(net41),
    .B(\hpos[6] ),
    .C(\hpos[8] ),
    .Y(_090_));
 sg13g2_nor2_1 _424_ (.A(net40),
    .B(_090_),
    .Y(_091_));
 sg13g2_o21ai_1 _425_ (.B1(_091_),
    .Y(_092_),
    .A1(\hpos[7] ),
    .A2(_055_));
 sg13g2_a21oi_1 _426_ (.A1(net40),
    .A2(_090_),
    .Y(_093_),
    .B1(_296_));
 sg13g2_and2_1 _427_ (.A(_092_),
    .B(_093_),
    .X(_094_));
 sg13g2_nor2_1 _428_ (.A(\hvsync_gen.vpos[8] ),
    .B(_286_),
    .Y(_095_));
 sg13g2_a22oi_1 _429_ (.Y(_096_),
    .B1(_095_),
    .B2(\hvsync_gen.vpos[9] ),
    .A2(_279_),
    .A1(net38));
 sg13g2_o21ai_1 _430_ (.B1(\hvsync_gen.vpos[9] ),
    .Y(_097_),
    .A1(\hvsync_gen.vpos[8] ),
    .A2(_286_));
 sg13g2_a21o_1 _431_ (.A2(_296_),
    .A1(\hpos[9] ),
    .B1(_097_),
    .X(_098_));
 sg13g2_o21ai_1 _432_ (.B1(_098_),
    .Y(_099_),
    .A1(_094_),
    .A2(_096_));
 sg13g2_a21o_1 _433_ (.A2(_059_),
    .A1(_057_),
    .B1(_099_),
    .X(_100_));
 sg13g2_a21oi_1 _434_ (.A1(_061_),
    .A2(_089_),
    .Y(_101_),
    .B1(_100_));
 sg13g2_a21o_2 _435_ (.A2(_089_),
    .A1(_061_),
    .B1(_100_),
    .X(_102_));
 sg13g2_nand3_1 _436_ (.B(_296_),
    .C(_097_),
    .A(\hpos[9] ),
    .Y(_103_));
 sg13g2_nand3_1 _437_ (.B(_096_),
    .C(_098_),
    .A(_094_),
    .Y(_104_));
 sg13g2_and2_1 _438_ (.A(_103_),
    .B(_104_),
    .X(_105_));
 sg13g2_nand2_1 _439_ (.Y(_106_),
    .A(_103_),
    .B(_104_));
 sg13g2_nand2_1 _440_ (.Y(_107_),
    .A(_102_),
    .B(_105_));
 sg13g2_nor3_1 _441_ (.A(_050_),
    .B(_101_),
    .C(_106_),
    .Y(_108_));
 sg13g2_a21oi_2 _442_ (.B1(_108_),
    .Y(_109_),
    .A2(net33),
    .A1(_294_));
 sg13g2_mux2_1 _443_ (.A0(_084_),
    .A1(_082_),
    .S(net33),
    .X(_110_));
 sg13g2_nand3b_1 _444_ (.B(_102_),
    .C(_105_),
    .Y(_111_),
    .A_N(_065_));
 sg13g2_o21ai_1 _445_ (.B1(_063_),
    .Y(_112_),
    .A1(_101_),
    .A2(_106_));
 sg13g2_nand3_1 _446_ (.B(_102_),
    .C(_105_),
    .A(_076_),
    .Y(_113_));
 sg13g2_o21ai_1 _447_ (.B1(_070_),
    .Y(_114_),
    .A1(_101_),
    .A2(_106_));
 sg13g2_a22oi_1 _448_ (.Y(_115_),
    .B1(_113_),
    .B2(_114_),
    .A2(_112_),
    .A1(_111_));
 sg13g2_nand4_1 _449_ (.B(_112_),
    .C(_113_),
    .A(_111_),
    .Y(_116_),
    .D(_114_));
 sg13g2_nor2b_1 _450_ (.A(_115_),
    .B_N(_116_),
    .Y(_117_));
 sg13g2_and2_1 _451_ (.A(net43),
    .B(_076_),
    .X(_118_));
 sg13g2_and2_1 _452_ (.A(net39),
    .B(_070_),
    .X(_119_));
 sg13g2_mux2_1 _453_ (.A0(_119_),
    .A1(_118_),
    .S(net33),
    .X(_120_));
 sg13g2_a21oi_1 _454_ (.A1(_116_),
    .A2(_120_),
    .Y(_121_),
    .B1(_115_));
 sg13g2_mux2_1 _455_ (.A0(_082_),
    .A1(_084_),
    .S(net33),
    .X(_122_));
 sg13g2_a21oi_1 _456_ (.A1(_102_),
    .A2(_105_),
    .Y(_123_),
    .B1(_065_));
 sg13g2_nand3_1 _457_ (.B(_102_),
    .C(_105_),
    .A(_063_),
    .Y(_124_));
 sg13g2_nor2b_2 _458_ (.A(_123_),
    .B_N(_124_),
    .Y(_125_));
 sg13g2_or2_1 _459_ (.X(_126_),
    .B(_125_),
    .A(_122_));
 sg13g2_and2_1 _460_ (.A(_122_),
    .B(_125_),
    .X(_127_));
 sg13g2_xor2_1 _461_ (.B(_125_),
    .A(_122_),
    .X(_128_));
 sg13g2_nand2b_1 _462_ (.Y(_129_),
    .B(_128_),
    .A_N(_121_));
 sg13g2_or2_1 _463_ (.X(_130_),
    .B(_110_),
    .A(_109_));
 sg13g2_and2_1 _464_ (.A(_126_),
    .B(_130_),
    .X(_131_));
 sg13g2_a22oi_1 _465_ (.Y(_132_),
    .B1(_129_),
    .B2(_131_),
    .A2(_110_),
    .A1(_109_));
 sg13g2_nand2_1 _466_ (.Y(_133_),
    .A(_043_),
    .B(net32));
 sg13g2_o21ai_1 _467_ (.B1(_133_),
    .Y(_134_),
    .A1(_047_),
    .A2(net33));
 sg13g2_nor2_1 _468_ (.A(_294_),
    .B(net33),
    .Y(_135_));
 sg13g2_a21oi_1 _469_ (.A1(_050_),
    .A2(net33),
    .Y(_136_),
    .B1(_135_));
 sg13g2_nor2b_1 _470_ (.A(_134_),
    .B_N(_136_),
    .Y(_137_));
 sg13g2_xor2_1 _471_ (.B(_136_),
    .A(_134_),
    .X(_138_));
 sg13g2_a221oi_1 _472_ (.B2(_131_),
    .C1(_138_),
    .B1(_129_),
    .A1(_109_),
    .Y(_139_),
    .A2(_110_));
 sg13g2_xor2_1 _473_ (.B(_138_),
    .A(_132_),
    .X(_140_));
 sg13g2_nand2_1 _474_ (.Y(_141_),
    .A(\anim_offset[1] ),
    .B(_277_));
 sg13g2_nor2_1 _475_ (.A(\anim_offset[1] ),
    .B(\anim_offset[2] ),
    .Y(_142_));
 sg13g2_nor2_1 _476_ (.A(net2),
    .B(_142_),
    .Y(_143_));
 sg13g2_a21oi_1 _477_ (.A1(_276_),
    .A2(_142_),
    .Y(_144_),
    .B1(net2));
 sg13g2_xnor2_1 _478_ (.Y(_145_),
    .A(\anim_offset[4] ),
    .B(_144_));
 sg13g2_nand2b_1 _479_ (.Y(_146_),
    .B(_145_),
    .A_N(_140_));
 sg13g2_xor2_1 _480_ (.B(_145_),
    .A(_140_),
    .X(_147_));
 sg13g2_xnor2_1 _481_ (.Y(_148_),
    .A(_276_),
    .B(_143_));
 sg13g2_xnor2_1 _482_ (.Y(_149_),
    .A(_117_),
    .B(_120_));
 sg13g2_xnor2_1 _483_ (.Y(_150_),
    .A(\anim_offset[2] ),
    .B(_141_));
 sg13g2_nand3_1 _484_ (.B(_149_),
    .C(_150_),
    .A(\anim_offset[1] ),
    .Y(_151_));
 sg13g2_a21oi_1 _485_ (.A1(\anim_offset[1] ),
    .A2(_149_),
    .Y(_152_),
    .B1(_150_));
 sg13g2_xnor2_1 _486_ (.Y(_153_),
    .A(_121_),
    .B(_128_));
 sg13g2_a21o_1 _487_ (.A2(_153_),
    .A1(_151_),
    .B1(_152_),
    .X(_154_));
 sg13g2_xor2_1 _488_ (.B(_110_),
    .A(_109_),
    .X(_155_));
 sg13g2_o21ai_1 _489_ (.B1(_126_),
    .Y(_156_),
    .A1(_121_),
    .A2(_127_));
 sg13g2_xnor2_1 _490_ (.Y(_157_),
    .A(_155_),
    .B(_156_));
 sg13g2_nor2_1 _491_ (.A(_148_),
    .B(_157_),
    .Y(_158_));
 sg13g2_nand2_1 _492_ (.Y(_159_),
    .A(_148_),
    .B(_157_));
 sg13g2_a21oi_1 _493_ (.A1(_154_),
    .A2(_159_),
    .Y(_160_),
    .B1(_158_));
 sg13g2_or2_1 _494_ (.X(_161_),
    .B(_160_),
    .A(_147_));
 sg13g2_o21ai_1 _495_ (.B1(\hpos[9] ),
    .Y(_162_),
    .A1(\hpos[7] ),
    .A2(\hpos[8] ));
 sg13g2_inv_1 _496_ (.Y(_163_),
    .A(_162_));
 sg13g2_nor3_2 _497_ (.A(\hvsync_gen.vpos[9] ),
    .B(_279_),
    .C(_163_),
    .Y(_164_));
 sg13g2_nand2_1 _498_ (.Y(_165_),
    .A(_161_),
    .B(_164_));
 sg13g2_a21oi_1 _499_ (.A1(_147_),
    .A2(_160_),
    .Y(uo_out[4]),
    .B1(_165_));
 sg13g2_nand2_1 _500_ (.Y(_166_),
    .A(_037_),
    .B(net31));
 sg13g2_o21ai_1 _501_ (.B1(_166_),
    .Y(_167_),
    .A1(_031_),
    .A2(net31));
 sg13g2_nor2_1 _502_ (.A(_043_),
    .B(net32),
    .Y(_168_));
 sg13g2_a21oi_1 _503_ (.A1(_047_),
    .A2(net32),
    .Y(_169_),
    .B1(_168_));
 sg13g2_inv_1 _504_ (.Y(_170_),
    .A(_169_));
 sg13g2_nand2_1 _505_ (.Y(_171_),
    .A(_167_),
    .B(_170_));
 sg13g2_xnor2_1 _506_ (.Y(_172_),
    .A(_167_),
    .B(_169_));
 sg13g2_nor3_1 _507_ (.A(_137_),
    .B(_139_),
    .C(_172_),
    .Y(_173_));
 sg13g2_o21ai_1 _508_ (.B1(_172_),
    .Y(_174_),
    .A1(_137_),
    .A2(_139_));
 sg13g2_nand2b_1 _509_ (.Y(_175_),
    .B(_174_),
    .A_N(_173_));
 sg13g2_nor3_1 _510_ (.A(\anim_offset[4] ),
    .B(\anim_offset[3] ),
    .C(_143_),
    .Y(_176_));
 sg13g2_nor2_1 _511_ (.A(net2),
    .B(_176_),
    .Y(_177_));
 sg13g2_xnor2_1 _512_ (.Y(_178_),
    .A(_278_),
    .B(_177_));
 sg13g2_nor2_1 _513_ (.A(_175_),
    .B(_178_),
    .Y(_179_));
 sg13g2_xnor2_1 _514_ (.Y(_180_),
    .A(_175_),
    .B(_178_));
 sg13g2_a21oi_1 _515_ (.A1(_146_),
    .A2(_161_),
    .Y(_181_),
    .B1(_180_));
 sg13g2_nand3_1 _516_ (.B(_161_),
    .C(_180_),
    .A(_146_),
    .Y(_182_));
 sg13g2_nand2_1 _517_ (.Y(_183_),
    .A(_164_),
    .B(_182_));
 sg13g2_nor2_2 _518_ (.A(_181_),
    .B(_183_),
    .Y(uo_out[5]));
 sg13g2_nor2_1 _519_ (.A(_057_),
    .B(net31),
    .Y(_184_));
 sg13g2_a21oi_1 _520_ (.A1(_059_),
    .A2(net31),
    .Y(_185_),
    .B1(_184_));
 sg13g2_nor2_1 _521_ (.A(_037_),
    .B(net31),
    .Y(_186_));
 sg13g2_a21oi_1 _522_ (.A1(_031_),
    .A2(net31),
    .Y(_187_),
    .B1(_186_));
 sg13g2_nor2b_1 _523_ (.A(_185_),
    .B_N(_187_),
    .Y(_188_));
 sg13g2_xor2_1 _524_ (.B(_187_),
    .A(_185_),
    .X(_189_));
 sg13g2_and3_1 _525_ (.X(_190_),
    .A(_171_),
    .B(_174_),
    .C(_189_));
 sg13g2_a21oi_1 _526_ (.A1(_171_),
    .A2(_174_),
    .Y(_191_),
    .B1(_189_));
 sg13g2_or2_1 _527_ (.X(_192_),
    .B(_191_),
    .A(_190_));
 sg13g2_a21oi_1 _528_ (.A1(_278_),
    .A2(_176_),
    .Y(_193_),
    .B1(net2));
 sg13g2_xor2_1 _529_ (.B(_193_),
    .A(\anim_offset[6] ),
    .X(_194_));
 sg13g2_or2_1 _530_ (.X(_195_),
    .B(_194_),
    .A(_192_));
 sg13g2_xor2_1 _531_ (.B(_194_),
    .A(_192_),
    .X(_196_));
 sg13g2_o21ai_1 _532_ (.B1(_196_),
    .Y(_197_),
    .A1(_179_),
    .A2(_181_));
 sg13g2_or3_1 _533_ (.A(_179_),
    .B(_181_),
    .C(_196_),
    .X(_198_));
 sg13g2_and3_2 _534_ (.X(uo_out[6]),
    .A(_164_),
    .B(_197_),
    .C(_198_));
 sg13g2_nor2_1 _535_ (.A(_188_),
    .B(_191_),
    .Y(_199_));
 sg13g2_xor2_1 _536_ (.B(_094_),
    .A(_059_),
    .X(_200_));
 sg13g2_nor2_1 _537_ (.A(net31),
    .B(_200_),
    .Y(_201_));
 sg13g2_xnor2_1 _538_ (.Y(_202_),
    .A(_057_),
    .B(_096_));
 sg13g2_a21oi_1 _539_ (.A1(net31),
    .A2(_202_),
    .Y(_203_),
    .B1(_201_));
 sg13g2_o21ai_1 _540_ (.B1(_277_),
    .Y(_204_),
    .A1(\anim_offset[6] ),
    .A2(_193_));
 sg13g2_xor2_1 _541_ (.B(_204_),
    .A(\anim_offset[7] ),
    .X(_205_));
 sg13g2_xnor2_1 _542_ (.Y(_206_),
    .A(_203_),
    .B(_205_));
 sg13g2_xnor2_1 _543_ (.Y(_207_),
    .A(_199_),
    .B(_206_));
 sg13g2_nand3_1 _544_ (.B(_197_),
    .C(_207_),
    .A(_195_),
    .Y(_208_));
 sg13g2_a21o_1 _545_ (.A2(_197_),
    .A1(_195_),
    .B1(_207_),
    .X(_209_));
 sg13g2_and3_1 _546_ (.X(uo_out[2]),
    .A(_164_),
    .B(_208_),
    .C(_209_));
 sg13g2_and3_2 _547_ (.X(_210_),
    .A(net43),
    .B(net99),
    .C(net65));
 sg13g2_and2_1 _548_ (.A(net89),
    .B(_210_),
    .X(_211_));
 sg13g2_nand2_1 _549_ (.Y(_212_),
    .A(net89),
    .B(_210_));
 sg13g2_nor2_1 _550_ (.A(_271_),
    .B(_212_),
    .Y(_213_));
 sg13g2_nor3_1 _551_ (.A(net83),
    .B(net41),
    .C(net42),
    .Y(_214_));
 sg13g2_and4_1 _552_ (.A(net85),
    .B(net40),
    .C(_213_),
    .D(_214_),
    .X(_215_));
 sg13g2_nor2b_2 _553_ (.A(_215_),
    .B_N(net44),
    .Y(_216_));
 sg13g2_nand2b_2 _554_ (.Y(_217_),
    .B(net44),
    .A_N(_215_));
 sg13g2_nor2_1 _555_ (.A(net43),
    .B(_217_),
    .Y(_002_));
 sg13g2_nor2_1 _556_ (.A(_067_),
    .B(_217_),
    .Y(_003_));
 sg13g2_a21oi_1 _557_ (.A1(net43),
    .A2(\cx[1] ),
    .Y(_218_),
    .B1(net65));
 sg13g2_nor3_1 _558_ (.A(_210_),
    .B(_217_),
    .C(net66),
    .Y(_004_));
 sg13g2_o21ai_1 _559_ (.B1(net44),
    .Y(_219_),
    .A1(net89),
    .A2(_210_));
 sg13g2_nor2_1 _560_ (.A(_211_),
    .B(net90),
    .Y(_005_));
 sg13g2_o21ai_1 _561_ (.B1(net44),
    .Y(_220_),
    .A1(net80),
    .A2(_211_));
 sg13g2_nor2_1 _562_ (.A(_213_),
    .B(net81),
    .Y(_006_));
 sg13g2_and2_1 _563_ (.A(net83),
    .B(_213_),
    .X(_221_));
 sg13g2_nor2_1 _564_ (.A(net83),
    .B(_213_),
    .Y(_222_));
 sg13g2_nor3_1 _565_ (.A(_217_),
    .B(_221_),
    .C(net84),
    .Y(_007_));
 sg13g2_xnor2_1 _566_ (.Y(_223_),
    .A(net42),
    .B(_221_));
 sg13g2_nor2_1 _567_ (.A(_217_),
    .B(_223_),
    .Y(_008_));
 sg13g2_a21oi_1 _568_ (.A1(net42),
    .A2(_221_),
    .Y(_224_),
    .B1(net41));
 sg13g2_nor2_1 _569_ (.A(_283_),
    .B(_212_),
    .Y(_225_));
 sg13g2_nor3_1 _570_ (.A(_217_),
    .B(_224_),
    .C(_225_),
    .Y(_009_));
 sg13g2_nor2_1 _571_ (.A(net85),
    .B(_225_),
    .Y(_226_));
 sg13g2_and2_1 _572_ (.A(net85),
    .B(_225_),
    .X(_227_));
 sg13g2_nor3_1 _573_ (.A(_217_),
    .B(net86),
    .C(_227_),
    .Y(_010_));
 sg13g2_o21ai_1 _574_ (.B1(net35),
    .Y(_228_),
    .A1(net40),
    .A2(_227_));
 sg13g2_a21oi_1 _575_ (.A1(net40),
    .A2(_227_),
    .Y(_011_),
    .B1(_228_));
 sg13g2_nor4_1 _576_ (.A(net36),
    .B(net37),
    .C(\hvsync_gen.vpos[7] ),
    .D(\hvsync_gen.vpos[6] ),
    .Y(_229_));
 sg13g2_inv_1 _577_ (.Y(_230_),
    .A(_229_));
 sg13g2_nor2_1 _578_ (.A(net40),
    .B(_289_),
    .Y(_231_));
 sg13g2_nand4_1 _579_ (.B(_090_),
    .C(_229_),
    .A(_292_),
    .Y(_232_),
    .D(_231_));
 sg13g2_nor3_1 _580_ (.A(net1),
    .B(_303_),
    .C(_232_),
    .Y(_233_));
 sg13g2_xor2_1 _581_ (.B(_233_),
    .A(net62),
    .X(_012_));
 sg13g2_nor2_1 _582_ (.A(net62),
    .B(net1),
    .Y(_234_));
 sg13g2_nor3_1 _583_ (.A(_303_),
    .B(_232_),
    .C(_234_),
    .Y(_235_));
 sg13g2_and2_1 _584_ (.A(net58),
    .B(_235_),
    .X(_236_));
 sg13g2_xor2_1 _585_ (.B(_235_),
    .A(net58),
    .X(_013_));
 sg13g2_and2_1 _586_ (.A(net74),
    .B(_236_),
    .X(_237_));
 sg13g2_xnor2_1 _587_ (.Y(_014_),
    .A(_276_),
    .B(_236_));
 sg13g2_and2_1 _588_ (.A(net56),
    .B(_237_),
    .X(_238_));
 sg13g2_xor2_1 _589_ (.B(_237_),
    .A(net56),
    .X(_015_));
 sg13g2_xnor2_1 _590_ (.Y(_016_),
    .A(_278_),
    .B(_238_));
 sg13g2_nand3_1 _591_ (.B(net93),
    .C(_238_),
    .A(net77),
    .Y(_239_));
 sg13g2_a21o_1 _592_ (.A2(_238_),
    .A1(net77),
    .B1(net93),
    .X(_240_));
 sg13g2_and2_1 _593_ (.A(_239_),
    .B(_240_),
    .X(_017_));
 sg13g2_xnor2_1 _594_ (.Y(_018_),
    .A(net60),
    .B(_239_));
 sg13g2_nor4_1 _595_ (.A(_280_),
    .B(_290_),
    .C(_096_),
    .D(_230_),
    .Y(_241_));
 sg13g2_nand3b_1 _596_ (.B(_215_),
    .C(net44),
    .Y(_242_),
    .A_N(_241_));
 sg13g2_inv_1 _597_ (.Y(_243_),
    .A(net34));
 sg13g2_nand2_1 _598_ (.Y(_244_),
    .A(net64),
    .B(net35));
 sg13g2_o21ai_1 _599_ (.B1(_244_),
    .Y(_019_),
    .A1(net64),
    .A2(net34));
 sg13g2_nand3_1 _600_ (.B(_073_),
    .C(_215_),
    .A(net44),
    .Y(_245_));
 sg13g2_o21ai_1 _601_ (.B1(_245_),
    .Y(_020_),
    .A1(_274_),
    .A2(_217_));
 sg13g2_nand2_1 _602_ (.Y(_246_),
    .A(net72),
    .B(net35));
 sg13g2_nand3_1 _603_ (.B(\cy[1] ),
    .C(\cy[2] ),
    .A(net64),
    .Y(_247_));
 sg13g2_xor2_1 _604_ (.B(_072_),
    .A(net72),
    .X(_248_));
 sg13g2_o21ai_1 _605_ (.B1(_246_),
    .Y(_021_),
    .A1(net34),
    .A2(_248_));
 sg13g2_nand2_1 _606_ (.Y(_249_),
    .A(net70),
    .B(net35));
 sg13g2_nor2_1 _607_ (.A(_280_),
    .B(_072_),
    .Y(_250_));
 sg13g2_or2_1 _608_ (.X(_251_),
    .B(_072_),
    .A(_280_));
 sg13g2_xor2_1 _609_ (.B(_247_),
    .A(net70),
    .X(_252_));
 sg13g2_o21ai_1 _610_ (.B1(_249_),
    .Y(_022_),
    .A1(net34),
    .A2(_252_));
 sg13g2_nand2_1 _611_ (.Y(_253_),
    .A(net37),
    .B(net35));
 sg13g2_xnor2_1 _612_ (.Y(_254_),
    .A(net37),
    .B(_250_));
 sg13g2_o21ai_1 _613_ (.B1(_253_),
    .Y(_023_),
    .A1(_242_),
    .A2(_254_));
 sg13g2_nand2_1 _614_ (.Y(_255_),
    .A(net36),
    .B(_216_));
 sg13g2_a21oi_1 _615_ (.A1(net37),
    .A2(_250_),
    .Y(_256_),
    .B1(net97));
 sg13g2_nor2_1 _616_ (.A(_285_),
    .B(_251_),
    .Y(_257_));
 sg13g2_or2_1 _617_ (.X(_258_),
    .B(_257_),
    .A(_256_));
 sg13g2_o21ai_1 _618_ (.B1(_255_),
    .Y(_024_),
    .A1(_242_),
    .A2(_258_));
 sg13g2_nand2_1 _619_ (.Y(_259_),
    .A(net76),
    .B(_216_));
 sg13g2_xnor2_1 _620_ (.Y(_260_),
    .A(net76),
    .B(_257_));
 sg13g2_o21ai_1 _621_ (.B1(_259_),
    .Y(_025_),
    .A1(net34),
    .A2(_260_));
 sg13g2_a21oi_1 _622_ (.A1(_033_),
    .A2(_250_),
    .Y(_261_),
    .B1(net78));
 sg13g2_nor2_1 _623_ (.A(_287_),
    .B(_251_),
    .Y(_262_));
 sg13g2_nor3_1 _624_ (.A(net34),
    .B(_261_),
    .C(_262_),
    .Y(_263_));
 sg13g2_a21o_1 _625_ (.A2(net35),
    .A1(net78),
    .B1(_263_),
    .X(_026_));
 sg13g2_nand2_1 _626_ (.Y(_264_),
    .A(net68),
    .B(_262_));
 sg13g2_nor2b_1 _627_ (.A(net34),
    .B_N(_264_),
    .Y(_265_));
 sg13g2_nor2_1 _628_ (.A(net35),
    .B(_265_),
    .Y(_266_));
 sg13g2_a21oi_1 _629_ (.A1(_243_),
    .A2(_262_),
    .Y(_267_),
    .B1(net68));
 sg13g2_nor2_1 _630_ (.A(_266_),
    .B(net69),
    .Y(_027_));
 sg13g2_o21ai_1 _631_ (.B1(net79),
    .Y(_268_),
    .A1(net35),
    .A2(_265_));
 sg13g2_or2_1 _632_ (.X(_269_),
    .B(_264_),
    .A(net79));
 sg13g2_o21ai_1 _633_ (.B1(_268_),
    .Y(_028_),
    .A1(net34),
    .A2(_269_));
 sg13g2_dfrbpq_2 _634_ (.RESET_B(net30),
    .D(_002_),
    .Q(\abs_x[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _635_ (.RESET_B(net53),
    .D(_003_),
    .Q(\cx[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _636_ (.RESET_B(net52),
    .D(net67),
    .Q(\cx[2] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _637_ (.RESET_B(net51),
    .D(_005_),
    .Q(\cx[3] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _638_ (.RESET_B(net50),
    .D(net82),
    .Q(\cx[4] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _639_ (.RESET_B(net49),
    .D(_007_),
    .Q(\cx[5] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _640_ (.RESET_B(net48),
    .D(_008_),
    .Q(\hpos[6] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _641_ (.RESET_B(net47),
    .D(_009_),
    .Q(\hpos[7] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _642_ (.RESET_B(net46),
    .D(_010_),
    .Q(\hpos[8] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _643_ (.RESET_B(net29),
    .D(_011_),
    .Q(\hpos[9] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _644_ (.RESET_B(net44),
    .D(net63),
    .Q(\anim_offset[1] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _645_ (.RESET_B(net44),
    .D(net59),
    .Q(\anim_offset[2] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _646_ (.RESET_B(net45),
    .D(_014_),
    .Q(\anim_offset[3] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _647_ (.RESET_B(net45),
    .D(net57),
    .Q(\anim_offset[4] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _648_ (.RESET_B(net45),
    .D(_016_),
    .Q(\anim_offset[5] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _649_ (.RESET_B(net45),
    .D(_017_),
    .Q(\anim_offset[6] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _650_ (.RESET_B(net45),
    .D(net61),
    .Q(\anim_offset[7] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _651_ (.RESET_B(net28),
    .D(net88),
    .Q(hsync),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _652_ (.RESET_B(net27),
    .D(_019_),
    .Q(\abs_y[0] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _653_ (.RESET_B(net25),
    .D(_020_),
    .Q(\cy[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _654_ (.RESET_B(net23),
    .D(net73),
    .Q(\cy[2] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _655_ (.RESET_B(net21),
    .D(net71),
    .Q(\cy[3] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _656_ (.RESET_B(net19),
    .D(_023_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_1 _657_ (.RESET_B(net54),
    .D(_024_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _658_ (.RESET_B(net24),
    .D(_025_),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _659_ (.RESET_B(net20),
    .D(_026_),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _660_ (.RESET_B(net26),
    .D(_027_),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _661_ (.RESET_B(net22),
    .D(_028_),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _662_ (.RESET_B(net55),
    .D(net95),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_tiehi _659__20 (.L_HI(net20));
 sg13g2_tiehi _655__21 (.L_HI(net21));
 sg13g2_tiehi _661__22 (.L_HI(net22));
 sg13g2_tiehi _654__23 (.L_HI(net23));
 sg13g2_tiehi _658__24 (.L_HI(net24));
 sg13g2_tiehi _653__25 (.L_HI(net25));
 sg13g2_tiehi _660__26 (.L_HI(net26));
 sg13g2_tiehi _652__27 (.L_HI(net27));
 sg13g2_tiehi _651__28 (.L_HI(net28));
 sg13g2_tiehi _643__29 (.L_HI(net29));
 sg13g2_tiehi _634__30 (.L_HI(net30));
 sg13g2_tiehi _642__31 (.L_HI(net46));
 sg13g2_tiehi _641__32 (.L_HI(net47));
 sg13g2_tiehi _640__33 (.L_HI(net48));
 sg13g2_tiehi _639__34 (.L_HI(net49));
 sg13g2_tiehi _638__35 (.L_HI(net50));
 sg13g2_tiehi _637__36 (.L_HI(net51));
 sg13g2_tiehi _636__37 (.L_HI(net52));
 sg13g2_tiehi _635__38 (.L_HI(net53));
 sg13g2_tiehi _657__39 (.L_HI(net54));
 sg13g2_tiehi _662__40 (.L_HI(net55));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_urish_rings_4 (.L_LO(net4));
 sg13g2_tielo tt_um_urish_rings_5 (.L_LO(net5));
 sg13g2_tielo tt_um_urish_rings_6 (.L_LO(net6));
 sg13g2_tielo tt_um_urish_rings_7 (.L_LO(net7));
 sg13g2_tielo tt_um_urish_rings_8 (.L_LO(net8));
 sg13g2_tielo tt_um_urish_rings_9 (.L_LO(net9));
 sg13g2_tielo tt_um_urish_rings_10 (.L_LO(net10));
 sg13g2_tielo tt_um_urish_rings_11 (.L_LO(net11));
 sg13g2_tielo tt_um_urish_rings_12 (.L_LO(net12));
 sg13g2_tielo tt_um_urish_rings_13 (.L_LO(net13));
 sg13g2_tielo tt_um_urish_rings_14 (.L_LO(net14));
 sg13g2_tielo tt_um_urish_rings_15 (.L_LO(net15));
 sg13g2_tielo tt_um_urish_rings_16 (.L_LO(net16));
 sg13g2_tielo tt_um_urish_rings_17 (.L_LO(net17));
 sg13g2_tielo tt_um_urish_rings_18 (.L_LO(net18));
 sg13g2_tiehi _656__19 (.L_HI(net19));
 sg13g2_buf_1 _701_ (.A(uo_out[5]),
    .X(uo_out[0]));
 sg13g2_buf_1 _702_ (.A(uo_out[6]),
    .X(uo_out[1]));
 sg13g2_buf_1 _703_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _704_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout31 (.A(net32),
    .X(net31));
 sg13g2_buf_1 fanout32 (.A(net33),
    .X(net32));
 sg13g2_buf_8 fanout33 (.A(_107_),
    .X(net33));
 sg13g2_buf_8 fanout34 (.A(_242_),
    .X(net34));
 sg13g2_buf_8 fanout35 (.A(_216_),
    .X(net35));
 sg13g2_buf_8 fanout36 (.A(net97),
    .X(net36));
 sg13g2_buf_8 fanout37 (.A(net94),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(net94),
    .X(net38));
 sg13g2_buf_8 fanout39 (.A(net64),
    .X(net39));
 sg13g2_buf_8 fanout40 (.A(net92),
    .X(net40));
 sg13g2_buf_8 fanout41 (.A(net87),
    .X(net41));
 sg13g2_buf_8 fanout42 (.A(net96),
    .X(net42));
 sg13g2_buf_8 fanout43 (.A(net75),
    .X(net43));
 sg13g2_buf_8 fanout44 (.A(rst_n),
    .X(net44));
 sg13g2_buf_8 fanout45 (.A(rst_n),
    .X(net45));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_tielo tt_um_urish_rings_3 (.L_LO(net3));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_4__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\anim_offset[4] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold2 (.A(_015_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold3 (.A(\anim_offset[2] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold4 (.A(_013_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold5 (.A(\anim_offset[7] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold6 (.A(_018_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold7 (.A(\anim_offset[1] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold8 (.A(_012_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold9 (.A(\abs_y[0] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold10 (.A(\cx[2] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold11 (.A(_218_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold12 (.A(_004_),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold13 (.A(\hvsync_gen.vpos[8] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold14 (.A(_267_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold15 (.A(\cy[3] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold16 (.A(_022_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold17 (.A(\cy[2] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold18 (.A(_021_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold19 (.A(\anim_offset[3] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold20 (.A(\abs_x[0] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold21 (.A(\hvsync_gen.vpos[6] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold22 (.A(\anim_offset[5] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold23 (.A(\hvsync_gen.vpos[7] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.vpos[9] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold25 (.A(\cx[4] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold26 (.A(_220_),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold27 (.A(_006_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold28 (.A(\cx[5] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold29 (.A(_222_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold30 (.A(\hpos[8] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold31 (.A(_226_),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold32 (.A(\hpos[7] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold33 (.A(_000_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold34 (.A(\cx[3] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold35 (.A(_219_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold36 (.A(\cy[1] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold37 (.A(\hpos[9] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold38 (.A(\anim_offset[6] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold39 (.A(\hvsync_gen.vpos[4] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold40 (.A(_001_),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold41 (.A(\hpos[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold42 (.A(\hvsync_gen.vpos[5] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold43 (.A(\cx[1] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold44 (.A(\cx[1] ),
    .X(net99));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_160 ();
 sg13g2_decap_8 FILLER_20_167 ();
 sg13g2_fill_2 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_215 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_decap_8 FILLER_20_232 ();
 sg13g2_decap_8 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_decap_8 FILLER_20_274 ();
 sg13g2_decap_8 FILLER_20_281 ();
 sg13g2_decap_8 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_302 ();
 sg13g2_decap_8 FILLER_20_309 ();
 sg13g2_decap_8 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_20_323 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_20_337 ();
 sg13g2_decap_8 FILLER_20_344 ();
 sg13g2_decap_8 FILLER_20_351 ();
 sg13g2_decap_8 FILLER_20_358 ();
 sg13g2_decap_8 FILLER_20_365 ();
 sg13g2_decap_8 FILLER_20_372 ();
 sg13g2_decap_8 FILLER_20_379 ();
 sg13g2_decap_8 FILLER_20_386 ();
 sg13g2_decap_8 FILLER_20_393 ();
 sg13g2_decap_8 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_147 ();
 sg13g2_fill_1 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_178 ();
 sg13g2_fill_2 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_189 ();
 sg13g2_decap_4 FILLER_21_199 ();
 sg13g2_fill_2 FILLER_21_203 ();
 sg13g2_fill_1 FILLER_21_223 ();
 sg13g2_decap_8 FILLER_21_264 ();
 sg13g2_decap_8 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_278 ();
 sg13g2_decap_8 FILLER_21_285 ();
 sg13g2_decap_8 FILLER_21_292 ();
 sg13g2_decap_8 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_306 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_327 ();
 sg13g2_decap_8 FILLER_21_334 ();
 sg13g2_decap_8 FILLER_21_341 ();
 sg13g2_decap_8 FILLER_21_348 ();
 sg13g2_decap_8 FILLER_21_355 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_138 ();
 sg13g2_decap_4 FILLER_22_170 ();
 sg13g2_decap_8 FILLER_22_192 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_22_211 ();
 sg13g2_decap_8 FILLER_22_222 ();
 sg13g2_fill_1 FILLER_22_229 ();
 sg13g2_fill_2 FILLER_22_239 ();
 sg13g2_fill_1 FILLER_22_241 ();
 sg13g2_decap_4 FILLER_22_246 ();
 sg13g2_decap_4 FILLER_22_281 ();
 sg13g2_decap_8 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_8 FILLER_22_303 ();
 sg13g2_decap_8 FILLER_22_310 ();
 sg13g2_decap_8 FILLER_22_317 ();
 sg13g2_decap_8 FILLER_22_324 ();
 sg13g2_decap_8 FILLER_22_331 ();
 sg13g2_decap_8 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_352 ();
 sg13g2_decap_8 FILLER_22_359 ();
 sg13g2_decap_8 FILLER_22_366 ();
 sg13g2_decap_8 FILLER_22_373 ();
 sg13g2_decap_8 FILLER_22_380 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_8 FILLER_22_394 ();
 sg13g2_decap_8 FILLER_22_401 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_4 FILLER_23_105 ();
 sg13g2_fill_2 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_115 ();
 sg13g2_fill_1 FILLER_23_145 ();
 sg13g2_fill_2 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_1 FILLER_23_221 ();
 sg13g2_decap_4 FILLER_23_239 ();
 sg13g2_fill_2 FILLER_23_243 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_decap_8 FILLER_23_302 ();
 sg13g2_decap_8 FILLER_23_309 ();
 sg13g2_decap_8 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_decap_8 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_344 ();
 sg13g2_decap_8 FILLER_23_351 ();
 sg13g2_decap_8 FILLER_23_358 ();
 sg13g2_decap_8 FILLER_23_365 ();
 sg13g2_decap_8 FILLER_23_372 ();
 sg13g2_decap_8 FILLER_23_379 ();
 sg13g2_decap_8 FILLER_23_386 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_decap_8 FILLER_23_400 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_fill_1 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_4 FILLER_24_159 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_decap_4 FILLER_24_179 ();
 sg13g2_fill_1 FILLER_24_183 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_4 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_4 FILLER_24_221 ();
 sg13g2_fill_1 FILLER_24_225 ();
 sg13g2_decap_4 FILLER_24_234 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_4 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_302 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_decap_8 FILLER_24_323 ();
 sg13g2_decap_8 FILLER_24_330 ();
 sg13g2_decap_8 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_344 ();
 sg13g2_decap_8 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_358 ();
 sg13g2_decap_8 FILLER_24_365 ();
 sg13g2_decap_8 FILLER_24_372 ();
 sg13g2_decap_8 FILLER_24_379 ();
 sg13g2_decap_8 FILLER_24_386 ();
 sg13g2_decap_8 FILLER_24_393 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_135 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_179 ();
 sg13g2_decap_8 FILLER_25_201 ();
 sg13g2_decap_4 FILLER_25_224 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_fill_2 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_263 ();
 sg13g2_fill_2 FILLER_25_277 ();
 sg13g2_fill_1 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_406 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_4 FILLER_26_130 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_decap_4 FILLER_26_160 ();
 sg13g2_fill_2 FILLER_26_164 ();
 sg13g2_decap_4 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_fill_2 FILLER_26_201 ();
 sg13g2_fill_2 FILLER_26_213 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_250 ();
 sg13g2_decap_4 FILLER_26_257 ();
 sg13g2_decap_8 FILLER_26_299 ();
 sg13g2_decap_8 FILLER_26_306 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_decap_8 FILLER_26_320 ();
 sg13g2_decap_8 FILLER_26_327 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_4 FILLER_26_404 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_102 ();
 sg13g2_fill_1 FILLER_27_104 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_163 ();
 sg13g2_decap_8 FILLER_27_172 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_decap_4 FILLER_27_230 ();
 sg13g2_fill_2 FILLER_27_234 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_decap_4 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_332 ();
 sg13g2_decap_8 FILLER_27_339 ();
 sg13g2_decap_8 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_353 ();
 sg13g2_decap_8 FILLER_27_360 ();
 sg13g2_decap_8 FILLER_27_367 ();
 sg13g2_decap_8 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_decap_8 FILLER_27_402 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_fill_2 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_127 ();
 sg13g2_decap_4 FILLER_28_134 ();
 sg13g2_decap_4 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_155 ();
 sg13g2_fill_1 FILLER_28_166 ();
 sg13g2_fill_2 FILLER_28_180 ();
 sg13g2_fill_2 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_194 ();
 sg13g2_fill_1 FILLER_28_205 ();
 sg13g2_decap_8 FILLER_28_215 ();
 sg13g2_decap_8 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_229 ();
 sg13g2_fill_1 FILLER_28_231 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_decap_4 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_decap_8 FILLER_28_282 ();
 sg13g2_fill_2 FILLER_28_298 ();
 sg13g2_fill_1 FILLER_28_300 ();
 sg13g2_fill_2 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_340 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_4 FILLER_29_77 ();
 sg13g2_fill_1 FILLER_29_81 ();
 sg13g2_fill_2 FILLER_29_137 ();
 sg13g2_fill_1 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_183 ();
 sg13g2_fill_1 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_4 FILLER_29_205 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_decap_4 FILLER_29_253 ();
 sg13g2_fill_2 FILLER_29_270 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_decap_4 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_295 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_fill_2 FILLER_29_327 ();
 sg13g2_fill_1 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_fill_2 FILLER_29_406 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_fill_1 FILLER_30_86 ();
 sg13g2_fill_2 FILLER_30_91 ();
 sg13g2_fill_1 FILLER_30_93 ();
 sg13g2_decap_4 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_226 ();
 sg13g2_fill_2 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_fill_2 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_271 ();
 sg13g2_fill_1 FILLER_30_275 ();
 sg13g2_decap_8 FILLER_30_297 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_decap_4 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_365 ();
 sg13g2_decap_8 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_4 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_2 FILLER_31_140 ();
 sg13g2_decap_4 FILLER_31_150 ();
 sg13g2_fill_1 FILLER_31_154 ();
 sg13g2_fill_2 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_173 ();
 sg13g2_decap_4 FILLER_31_180 ();
 sg13g2_fill_2 FILLER_31_184 ();
 sg13g2_decap_8 FILLER_31_197 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_fill_2 FILLER_31_227 ();
 sg13g2_fill_1 FILLER_31_229 ();
 sg13g2_fill_2 FILLER_31_235 ();
 sg13g2_fill_1 FILLER_31_237 ();
 sg13g2_decap_4 FILLER_31_243 ();
 sg13g2_decap_4 FILLER_31_257 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_fill_2 FILLER_31_278 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_fill_1 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_292 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_319 ();
 sg13g2_decap_4 FILLER_31_326 ();
 sg13g2_fill_2 FILLER_31_330 ();
 sg13g2_decap_4 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_340 ();
 sg13g2_decap_4 FILLER_31_345 ();
 sg13g2_fill_1 FILLER_31_349 ();
 sg13g2_decap_8 FILLER_31_355 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_8 FILLER_32_148 ();
 sg13g2_decap_8 FILLER_32_170 ();
 sg13g2_fill_2 FILLER_32_177 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_190 ();
 sg13g2_decap_4 FILLER_32_201 ();
 sg13g2_fill_1 FILLER_32_205 ();
 sg13g2_decap_8 FILLER_32_218 ();
 sg13g2_fill_1 FILLER_32_225 ();
 sg13g2_decap_4 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_253 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_4 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_4 FILLER_32_305 ();
 sg13g2_fill_1 FILLER_32_309 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_343 ();
 sg13g2_fill_1 FILLER_32_352 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_79 ();
 sg13g2_fill_2 FILLER_33_108 ();
 sg13g2_fill_1 FILLER_33_110 ();
 sg13g2_decap_8 FILLER_33_146 ();
 sg13g2_decap_8 FILLER_33_166 ();
 sg13g2_decap_8 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_180 ();
 sg13g2_decap_8 FILLER_33_207 ();
 sg13g2_decap_4 FILLER_33_214 ();
 sg13g2_fill_2 FILLER_33_218 ();
 sg13g2_decap_4 FILLER_33_224 ();
 sg13g2_fill_2 FILLER_33_228 ();
 sg13g2_fill_2 FILLER_33_235 ();
 sg13g2_fill_2 FILLER_33_253 ();
 sg13g2_decap_8 FILLER_33_264 ();
 sg13g2_fill_2 FILLER_33_279 ();
 sg13g2_fill_1 FILLER_33_281 ();
 sg13g2_decap_4 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_320 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_342 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_decap_8 FILLER_33_389 ();
 sg13g2_decap_8 FILLER_33_396 ();
 sg13g2_decap_4 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_407 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_107 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_123 ();
 sg13g2_fill_2 FILLER_34_168 ();
 sg13g2_fill_2 FILLER_34_181 ();
 sg13g2_fill_1 FILLER_34_183 ();
 sg13g2_fill_1 FILLER_34_189 ();
 sg13g2_decap_8 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_213 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_decap_4 FILLER_34_265 ();
 sg13g2_fill_2 FILLER_34_269 ();
 sg13g2_decap_8 FILLER_34_276 ();
 sg13g2_decap_8 FILLER_34_283 ();
 sg13g2_decap_8 FILLER_34_290 ();
 sg13g2_decap_4 FILLER_34_297 ();
 sg13g2_fill_2 FILLER_34_301 ();
 sg13g2_decap_8 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_fill_2 FILLER_34_326 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_decap_4 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_399 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_88 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_fill_1 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_decap_4 FILLER_35_172 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_1 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_decap_4 FILLER_35_242 ();
 sg13g2_fill_2 FILLER_35_246 ();
 sg13g2_decap_4 FILLER_35_253 ();
 sg13g2_fill_1 FILLER_35_261 ();
 sg13g2_decap_4 FILLER_35_273 ();
 sg13g2_fill_2 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_decap_4 FILLER_35_319 ();
 sg13g2_fill_1 FILLER_35_323 ();
 sg13g2_fill_2 FILLER_35_337 ();
 sg13g2_fill_1 FILLER_35_339 ();
 sg13g2_fill_1 FILLER_35_353 ();
 sg13g2_decap_8 FILLER_35_398 ();
 sg13g2_decap_4 FILLER_35_405 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_fill_2 FILLER_36_91 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_2 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_decap_8 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_fill_2 FILLER_36_220 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_fill_2 FILLER_36_233 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_276 ();
 sg13g2_decap_8 FILLER_36_283 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_fill_1 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_4 FILLER_36_322 ();
 sg13g2_decap_4 FILLER_36_334 ();
 sg13g2_fill_2 FILLER_36_355 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_decap_8 FILLER_36_380 ();
 sg13g2_decap_8 FILLER_36_387 ();
 sg13g2_decap_8 FILLER_36_394 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_4 FILLER_37_105 ();
 sg13g2_fill_2 FILLER_37_109 ();
 sg13g2_fill_1 FILLER_37_166 ();
 sg13g2_decap_8 FILLER_37_198 ();
 sg13g2_decap_8 FILLER_37_205 ();
 sg13g2_decap_8 FILLER_37_212 ();
 sg13g2_decap_8 FILLER_37_223 ();
 sg13g2_decap_8 FILLER_37_230 ();
 sg13g2_fill_1 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_251 ();
 sg13g2_decap_4 FILLER_37_258 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_decap_4 FILLER_37_284 ();
 sg13g2_fill_2 FILLER_37_321 ();
 sg13g2_fill_1 FILLER_37_323 ();
 sg13g2_fill_2 FILLER_37_332 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_390 ();
 sg13g2_decap_8 FILLER_37_397 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_151 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_219 ();
 sg13g2_decap_8 FILLER_38_226 ();
 sg13g2_decap_8 FILLER_38_233 ();
 sg13g2_decap_8 FILLER_38_240 ();
 sg13g2_decap_8 FILLER_38_247 ();
 sg13g2_decap_8 FILLER_38_254 ();
 sg13g2_decap_8 FILLER_38_261 ();
 sg13g2_fill_1 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_4 FILLER_38_322 ();
 sg13g2_fill_2 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_395 ();
 sg13g2_decap_8 FILLER_38_402 ();
 assign uio_oe[0] = net3;
 assign uio_oe[1] = net4;
 assign uio_oe[2] = net5;
 assign uio_oe[3] = net6;
 assign uio_oe[4] = net7;
 assign uio_oe[5] = net8;
 assign uio_oe[6] = net9;
 assign uio_oe[7] = net10;
 assign uio_out[0] = net11;
 assign uio_out[1] = net12;
 assign uio_out[2] = net13;
 assign uio_out[3] = net14;
 assign uio_out[4] = net15;
 assign uio_out[5] = net16;
 assign uio_out[6] = net17;
 assign uio_out[7] = net18;
endmodule
