module tt_um_pgfarley_tophat_top (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire clear_cmd;
 wire core_busy;
 wire core_error;
 wire \feature_byte[0] ;
 wire \feature_byte[1] ;
 wire \feature_byte[2] ;
 wire \feature_byte[3] ;
 wire \feature_byte[4] ;
 wire \feature_byte[5] ;
 wire \feature_byte[6] ;
 wire \feature_byte[7] ;
 wire feature_byte_valid;
 wire \feature_vector_flat[0] ;
 wire \feature_vector_flat[10] ;
 wire \feature_vector_flat[11] ;
 wire \feature_vector_flat[12] ;
 wire \feature_vector_flat[13] ;
 wire \feature_vector_flat[14] ;
 wire \feature_vector_flat[15] ;
 wire \feature_vector_flat[16] ;
 wire \feature_vector_flat[17] ;
 wire \feature_vector_flat[18] ;
 wire \feature_vector_flat[19] ;
 wire \feature_vector_flat[1] ;
 wire \feature_vector_flat[20] ;
 wire \feature_vector_flat[21] ;
 wire \feature_vector_flat[22] ;
 wire \feature_vector_flat[23] ;
 wire \feature_vector_flat[24] ;
 wire \feature_vector_flat[25] ;
 wire \feature_vector_flat[26] ;
 wire \feature_vector_flat[27] ;
 wire \feature_vector_flat[28] ;
 wire \feature_vector_flat[29] ;
 wire \feature_vector_flat[2] ;
 wire \feature_vector_flat[30] ;
 wire \feature_vector_flat[31] ;
 wire \feature_vector_flat[32] ;
 wire \feature_vector_flat[33] ;
 wire \feature_vector_flat[34] ;
 wire \feature_vector_flat[35] ;
 wire \feature_vector_flat[36] ;
 wire \feature_vector_flat[37] ;
 wire \feature_vector_flat[38] ;
 wire \feature_vector_flat[39] ;
 wire \feature_vector_flat[3] ;
 wire \feature_vector_flat[40] ;
 wire \feature_vector_flat[41] ;
 wire \feature_vector_flat[42] ;
 wire \feature_vector_flat[43] ;
 wire \feature_vector_flat[44] ;
 wire \feature_vector_flat[45] ;
 wire \feature_vector_flat[46] ;
 wire \feature_vector_flat[47] ;
 wire \feature_vector_flat[48] ;
 wire \feature_vector_flat[49] ;
 wire \feature_vector_flat[4] ;
 wire \feature_vector_flat[50] ;
 wire \feature_vector_flat[51] ;
 wire \feature_vector_flat[52] ;
 wire \feature_vector_flat[53] ;
 wire \feature_vector_flat[54] ;
 wire \feature_vector_flat[55] ;
 wire \feature_vector_flat[56] ;
 wire \feature_vector_flat[57] ;
 wire \feature_vector_flat[58] ;
 wire \feature_vector_flat[59] ;
 wire \feature_vector_flat[5] ;
 wire \feature_vector_flat[60] ;
 wire \feature_vector_flat[61] ;
 wire \feature_vector_flat[62] ;
 wire \feature_vector_flat[63] ;
 wire \feature_vector_flat[6] ;
 wire \feature_vector_flat[7] ;
 wire \feature_vector_flat[8] ;
 wire \feature_vector_flat[9] ;
 wire features_loaded;
 wire io_ready;
 wire \leaf_value_flat[0] ;
 wire \leaf_value_flat[10] ;
 wire \leaf_value_flat[11] ;
 wire \leaf_value_flat[12] ;
 wire \leaf_value_flat[13] ;
 wire \leaf_value_flat[14] ;
 wire \leaf_value_flat[15] ;
 wire \leaf_value_flat[16] ;
 wire \leaf_value_flat[17] ;
 wire \leaf_value_flat[18] ;
 wire \leaf_value_flat[19] ;
 wire \leaf_value_flat[1] ;
 wire \leaf_value_flat[20] ;
 wire \leaf_value_flat[21] ;
 wire \leaf_value_flat[22] ;
 wire \leaf_value_flat[23] ;
 wire \leaf_value_flat[24] ;
 wire \leaf_value_flat[25] ;
 wire \leaf_value_flat[26] ;
 wire \leaf_value_flat[27] ;
 wire \leaf_value_flat[28] ;
 wire \leaf_value_flat[29] ;
 wire \leaf_value_flat[2] ;
 wire \leaf_value_flat[30] ;
 wire \leaf_value_flat[31] ;
 wire \leaf_value_flat[32] ;
 wire \leaf_value_flat[33] ;
 wire \leaf_value_flat[34] ;
 wire \leaf_value_flat[35] ;
 wire \leaf_value_flat[36] ;
 wire \leaf_value_flat[37] ;
 wire \leaf_value_flat[38] ;
 wire \leaf_value_flat[39] ;
 wire \leaf_value_flat[3] ;
 wire \leaf_value_flat[40] ;
 wire \leaf_value_flat[41] ;
 wire \leaf_value_flat[42] ;
 wire \leaf_value_flat[43] ;
 wire \leaf_value_flat[44] ;
 wire \leaf_value_flat[45] ;
 wire \leaf_value_flat[46] ;
 wire \leaf_value_flat[47] ;
 wire \leaf_value_flat[48] ;
 wire \leaf_value_flat[49] ;
 wire \leaf_value_flat[4] ;
 wire \leaf_value_flat[50] ;
 wire \leaf_value_flat[51] ;
 wire \leaf_value_flat[52] ;
 wire \leaf_value_flat[53] ;
 wire \leaf_value_flat[54] ;
 wire \leaf_value_flat[55] ;
 wire \leaf_value_flat[56] ;
 wire \leaf_value_flat[57] ;
 wire \leaf_value_flat[58] ;
 wire \leaf_value_flat[59] ;
 wire \leaf_value_flat[5] ;
 wire \leaf_value_flat[60] ;
 wire \leaf_value_flat[61] ;
 wire \leaf_value_flat[62] ;
 wire \leaf_value_flat[63] ;
 wire \leaf_value_flat[6] ;
 wire \leaf_value_flat[7] ;
 wire \leaf_value_flat[8] ;
 wire \leaf_value_flat[9] ;
 wire \model_byte[0] ;
 wire \model_byte[1] ;
 wire \model_byte[2] ;
 wire \model_byte[3] ;
 wire \model_byte[4] ;
 wire \model_byte[5] ;
 wire \model_byte[6] ;
 wire \model_byte[7] ;
 wire model_byte_valid;
 wire model_loaded;
 wire \node_feature_flat[0] ;
 wire \node_feature_flat[10] ;
 wire \node_feature_flat[11] ;
 wire \node_feature_flat[12] ;
 wire \node_feature_flat[13] ;
 wire \node_feature_flat[14] ;
 wire \node_feature_flat[15] ;
 wire \node_feature_flat[16] ;
 wire \node_feature_flat[17] ;
 wire \node_feature_flat[18] ;
 wire \node_feature_flat[19] ;
 wire \node_feature_flat[1] ;
 wire \node_feature_flat[20] ;
 wire \node_feature_flat[2] ;
 wire \node_feature_flat[3] ;
 wire \node_feature_flat[4] ;
 wire \node_feature_flat[5] ;
 wire \node_feature_flat[6] ;
 wire \node_feature_flat[7] ;
 wire \node_feature_flat[8] ;
 wire \node_feature_flat[9] ;
 wire \node_left_flat[0] ;
 wire \node_left_flat[10] ;
 wire \node_left_flat[11] ;
 wire \node_left_flat[12] ;
 wire \node_left_flat[13] ;
 wire \node_left_flat[14] ;
 wire \node_left_flat[15] ;
 wire \node_left_flat[16] ;
 wire \node_left_flat[17] ;
 wire \node_left_flat[18] ;
 wire \node_left_flat[19] ;
 wire \node_left_flat[1] ;
 wire \node_left_flat[20] ;
 wire \node_left_flat[21] ;
 wire \node_left_flat[22] ;
 wire \node_left_flat[23] ;
 wire \node_left_flat[24] ;
 wire \node_left_flat[25] ;
 wire \node_left_flat[26] ;
 wire \node_left_flat[27] ;
 wire \node_left_flat[2] ;
 wire \node_left_flat[3] ;
 wire \node_left_flat[4] ;
 wire \node_left_flat[5] ;
 wire \node_left_flat[6] ;
 wire \node_left_flat[7] ;
 wire \node_left_flat[8] ;
 wire \node_left_flat[9] ;
 wire \node_right_flat[0] ;
 wire \node_right_flat[10] ;
 wire \node_right_flat[11] ;
 wire \node_right_flat[12] ;
 wire \node_right_flat[13] ;
 wire \node_right_flat[14] ;
 wire \node_right_flat[15] ;
 wire \node_right_flat[16] ;
 wire \node_right_flat[17] ;
 wire \node_right_flat[18] ;
 wire \node_right_flat[19] ;
 wire \node_right_flat[1] ;
 wire \node_right_flat[20] ;
 wire \node_right_flat[21] ;
 wire \node_right_flat[22] ;
 wire \node_right_flat[23] ;
 wire \node_right_flat[24] ;
 wire \node_right_flat[25] ;
 wire \node_right_flat[26] ;
 wire \node_right_flat[27] ;
 wire \node_right_flat[2] ;
 wire \node_right_flat[3] ;
 wire \node_right_flat[4] ;
 wire \node_right_flat[5] ;
 wire \node_right_flat[6] ;
 wire \node_right_flat[7] ;
 wire \node_right_flat[8] ;
 wire \node_right_flat[9] ;
 wire \node_threshold_flat[0] ;
 wire \node_threshold_flat[10] ;
 wire \node_threshold_flat[11] ;
 wire \node_threshold_flat[12] ;
 wire \node_threshold_flat[13] ;
 wire \node_threshold_flat[14] ;
 wire \node_threshold_flat[15] ;
 wire \node_threshold_flat[16] ;
 wire \node_threshold_flat[17] ;
 wire \node_threshold_flat[18] ;
 wire \node_threshold_flat[19] ;
 wire \node_threshold_flat[1] ;
 wire \node_threshold_flat[20] ;
 wire \node_threshold_flat[21] ;
 wire \node_threshold_flat[22] ;
 wire \node_threshold_flat[23] ;
 wire \node_threshold_flat[24] ;
 wire \node_threshold_flat[25] ;
 wire \node_threshold_flat[26] ;
 wire \node_threshold_flat[27] ;
 wire \node_threshold_flat[28] ;
 wire \node_threshold_flat[29] ;
 wire \node_threshold_flat[2] ;
 wire \node_threshold_flat[30] ;
 wire \node_threshold_flat[31] ;
 wire \node_threshold_flat[32] ;
 wire \node_threshold_flat[33] ;
 wire \node_threshold_flat[34] ;
 wire \node_threshold_flat[35] ;
 wire \node_threshold_flat[36] ;
 wire \node_threshold_flat[37] ;
 wire \node_threshold_flat[38] ;
 wire \node_threshold_flat[39] ;
 wire \node_threshold_flat[3] ;
 wire \node_threshold_flat[40] ;
 wire \node_threshold_flat[41] ;
 wire \node_threshold_flat[42] ;
 wire \node_threshold_flat[43] ;
 wire \node_threshold_flat[44] ;
 wire \node_threshold_flat[45] ;
 wire \node_threshold_flat[46] ;
 wire \node_threshold_flat[47] ;
 wire \node_threshold_flat[48] ;
 wire \node_threshold_flat[49] ;
 wire \node_threshold_flat[4] ;
 wire \node_threshold_flat[50] ;
 wire \node_threshold_flat[51] ;
 wire \node_threshold_flat[52] ;
 wire \node_threshold_flat[53] ;
 wire \node_threshold_flat[54] ;
 wire \node_threshold_flat[55] ;
 wire \node_threshold_flat[5] ;
 wire \node_threshold_flat[6] ;
 wire \node_threshold_flat[7] ;
 wire \node_threshold_flat[8] ;
 wire \node_threshold_flat[9] ;
 wire pred_valid;
 wire run_cmd;
 wire \u_feature_loader.feature_idx_q[0] ;
 wire \u_feature_loader.feature_idx_q[1] ;
 wire \u_feature_loader.feature_idx_q[2] ;
 wire \u_feature_loader.feature_idx_q[3] ;
 wire \u_model_loader.byte_idx_q[0] ;
 wire \u_model_loader.byte_idx_q[1] ;
 wire \u_model_loader.byte_idx_q[2] ;
 wire \u_model_loader.byte_idx_q[3] ;
 wire \u_model_loader.byte_idx_q[4] ;
 wire \u_model_loader.byte_idx_q[5] ;
 wire \u_tree_core.current_node_q[0] ;
 wire \u_tree_core.current_node_q[1] ;
 wire \u_tree_core.current_node_q[2] ;
 wire \u_tree_core.depth_q[0] ;
 wire \u_tree_core.depth_q[1] ;
 wire \u_tree_core.state_q[0] ;
 wire \u_tree_core.state_q[1] ;
 wire net14;
 wire net15;
 wire net16;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire clknet_leaf_0_clk;
 wire net17;
 wire net18;
 wire net19;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;

 sg13g2_inv_2 _1468_ (.Y(_0820_),
    .A(\u_tree_core.current_node_q[2] ));
 sg13g2_inv_1 _1469_ (.Y(_0821_),
    .A(\u_tree_core.current_node_q[1] ));
 sg13g2_inv_4 _1470_ (.A(net536),
    .Y(_0822_));
 sg13g2_inv_1 _1471_ (.Y(_0823_),
    .A(net738));
 sg13g2_inv_1 _1472_ (.Y(io_ready),
    .A(net688));
 sg13g2_inv_1 _1473_ (.Y(_0824_),
    .A(\feature_vector_flat[63] ));
 sg13g2_inv_1 _1474_ (.Y(_0825_),
    .A(feature_byte_valid));
 sg13g2_inv_1 _1475_ (.Y(_0826_),
    .A(\feature_vector_flat[61] ));
 sg13g2_inv_1 _1476_ (.Y(_0827_),
    .A(\feature_vector_flat[59] ));
 sg13g2_inv_1 _1477_ (.Y(_0828_),
    .A(\feature_vector_flat[57] ));
 sg13g2_inv_1 _1478_ (.Y(_0829_),
    .A(net617));
 sg13g2_inv_1 _1479_ (.Y(_0830_),
    .A(net339));
 sg13g2_inv_1 _1480_ (.Y(_0831_),
    .A(net591));
 sg13g2_inv_1 _1481_ (.Y(_0832_),
    .A(net588));
 sg13g2_inv_1 _1482_ (.Y(_0833_),
    .A(net563));
 sg13g2_inv_1 _1483_ (.Y(_0834_),
    .A(net348));
 sg13g2_inv_1 _1484_ (.Y(_0835_),
    .A(net631));
 sg13g2_inv_1 _1485_ (.Y(_0836_),
    .A(net346));
 sg13g2_inv_1 _1486_ (.Y(_0837_),
    .A(net567));
 sg13g2_inv_1 _1487_ (.Y(_0838_),
    .A(net570));
 sg13g2_inv_1 _1488_ (.Y(_0839_),
    .A(net565));
 sg13g2_inv_1 _1489_ (.Y(_0840_),
    .A(net359));
 sg13g2_inv_1 _1490_ (.Y(_0841_),
    .A(net354));
 sg13g2_inv_1 _1491_ (.Y(_0842_),
    .A(net350));
 sg13g2_inv_1 _1492_ (.Y(_0843_),
    .A(net345));
 sg13g2_inv_1 _1493_ (.Y(_0844_),
    .A(\node_threshold_flat[15] ));
 sg13g2_inv_1 _1494_ (.Y(_0845_),
    .A(\node_threshold_flat[14] ));
 sg13g2_inv_1 _1495_ (.Y(_0846_),
    .A(\node_threshold_flat[13] ));
 sg13g2_inv_1 _1496_ (.Y(_0847_),
    .A(\node_threshold_flat[12] ));
 sg13g2_inv_1 _1497_ (.Y(_0848_),
    .A(net374));
 sg13g2_inv_1 _1498_ (.Y(_0849_),
    .A(\node_threshold_flat[10] ));
 sg13g2_inv_1 _1499_ (.Y(_0850_),
    .A(\node_threshold_flat[9] ));
 sg13g2_inv_1 _1500_ (.Y(_0851_),
    .A(\node_threshold_flat[8] ));
 sg13g2_inv_1 _1501_ (.Y(_0852_),
    .A(net671));
 sg13g2_inv_1 _1502_ (.Y(_0853_),
    .A(net577));
 sg13g2_inv_1 _1503_ (.Y(_0854_),
    .A(net609));
 sg13g2_inv_1 _1504_ (.Y(_0855_),
    .A(net599));
 sg13g2_inv_1 _1505_ (.Y(_0856_),
    .A(net363));
 sg13g2_inv_1 _1506_ (.Y(_0857_),
    .A(net370));
 sg13g2_inv_1 _1507_ (.Y(_0858_),
    .A(net335));
 sg13g2_inv_1 _1508_ (.Y(_0859_),
    .A(net568));
 sg13g2_inv_1 _1509_ (.Y(_0860_),
    .A(net603));
 sg13g2_inv_1 _1510_ (.Y(_0861_),
    .A(\node_left_flat[14] ));
 sg13g2_inv_1 _1511_ (.Y(_0862_),
    .A(\node_left_flat[13] ));
 sg13g2_inv_1 _1512_ (.Y(_0863_),
    .A(\node_left_flat[12] ));
 sg13g2_inv_1 _1513_ (.Y(_0864_),
    .A(\node_left_flat[8] ));
 sg13g2_inv_1 _1514_ (.Y(_0865_),
    .A(net337));
 sg13g2_inv_1 _1515_ (.Y(_0866_),
    .A(\node_left_flat[4] ));
 sg13g2_inv_1 _1516_ (.Y(_0867_),
    .A(net368));
 sg13g2_inv_1 _1517_ (.Y(_0868_),
    .A(\node_left_flat[0] ));
 sg13g2_inv_1 _1518_ (.Y(_0869_),
    .A(net341));
 sg13g2_inv_1 _1519_ (.Y(_0870_),
    .A(\node_right_flat[26] ));
 sg13g2_inv_1 _1520_ (.Y(_0871_),
    .A(\node_right_flat[24] ));
 sg13g2_inv_1 _1521_ (.Y(_0872_),
    .A(net559));
 sg13g2_inv_1 _1522_ (.Y(_0873_),
    .A(net352));
 sg13g2_inv_1 _1523_ (.Y(_0874_),
    .A(\node_right_flat[15] ));
 sg13g2_inv_1 _1524_ (.Y(_0875_),
    .A(\node_right_flat[14] ));
 sg13g2_inv_1 _1525_ (.Y(_0876_),
    .A(\node_right_flat[13] ));
 sg13g2_inv_1 _1526_ (.Y(_0877_),
    .A(\node_right_flat[12] ));
 sg13g2_inv_1 _1527_ (.Y(_0878_),
    .A(\node_right_flat[8] ));
 sg13g2_inv_1 _1528_ (.Y(_0879_),
    .A(net366));
 sg13g2_inv_1 _1529_ (.Y(_0880_),
    .A(\node_right_flat[4] ));
 sg13g2_inv_1 _1530_ (.Y(_0881_),
    .A(net343));
 sg13g2_inv_1 _1531_ (.Y(_0882_),
    .A(\node_right_flat[0] ));
 sg13g2_inv_1 _1532_ (.Y(_0883_),
    .A(\leaf_value_flat[43] ));
 sg13g2_inv_1 _1533_ (.Y(_0884_),
    .A(\leaf_value_flat[35] ));
 sg13g2_inv_2 _1534_ (.Y(_0885_),
    .A(\u_model_loader.byte_idx_q[2] ));
 sg13g2_inv_1 _1535_ (.Y(_0886_),
    .A(\model_byte[7] ));
 sg13g2_inv_1 _1536_ (.Y(_0887_),
    .A(net9));
 sg13g2_inv_2 _1537_ (.Y(_0888_),
    .A(\model_byte[6] ));
 sg13g2_inv_1 _1538_ (.Y(_0889_),
    .A(net8));
 sg13g2_inv_1 _1539_ (.Y(_0890_),
    .A(\model_byte[5] ));
 sg13g2_inv_1 _1540_ (.Y(_0891_),
    .A(net7));
 sg13g2_inv_2 _1541_ (.Y(_0892_),
    .A(\model_byte[4] ));
 sg13g2_inv_1 _1542_ (.Y(_0893_),
    .A(net6));
 sg13g2_inv_2 _1543_ (.Y(_0894_),
    .A(net548));
 sg13g2_inv_1 _1544_ (.Y(_0895_),
    .A(net5));
 sg13g2_inv_4 _1545_ (.A(net550),
    .Y(_0896_));
 sg13g2_inv_1 _1546_ (.Y(_0897_),
    .A(net4));
 sg13g2_inv_4 _1547_ (.A(net551),
    .Y(_0898_));
 sg13g2_inv_1 _1548_ (.Y(_0899_),
    .A(net3));
 sg13g2_inv_1 _1549_ (.Y(_0900_),
    .A(\model_byte[0] ));
 sg13g2_inv_1 _1550_ (.Y(_0901_),
    .A(net2));
 sg13g2_inv_1 _1551_ (.Y(_0902_),
    .A(\u_tree_core.state_q[0] ));
 sg13g2_inv_1 _1552_ (.Y(_0903_),
    .A(net11));
 sg13g2_nor2b_1 _1553_ (.A(clear_cmd),
    .B_N(net554),
    .Y(_0904_));
 sg13g2_nand2b_2 _1554_ (.Y(_0905_),
    .B(net554),
    .A_N(clear_cmd));
 sg13g2_a21oi_1 _1555_ (.A1(net539),
    .A2(_0845_),
    .Y(_0906_),
    .B1(net534));
 sg13g2_o21ai_1 _1556_ (.B1(_0906_),
    .Y(_0907_),
    .A1(net539),
    .A2(\node_threshold_flat[6] ));
 sg13g2_nor2b_1 _1557_ (.A(net541),
    .B_N(\u_tree_core.current_node_q[1] ),
    .Y(_0908_));
 sg13g2_nand2_2 _1558_ (.Y(_0909_),
    .A(net535),
    .B(_0822_));
 sg13g2_and2_1 _1559_ (.A(net534),
    .B(net542),
    .X(_0910_));
 sg13g2_a221oi_1 _1560_ (.B2(\node_threshold_flat[30] ),
    .C1(net533),
    .B1(net464),
    .A1(\node_threshold_flat[22] ),
    .Y(_0911_),
    .A2(net467));
 sg13g2_mux2_1 _1561_ (.A0(\node_threshold_flat[38] ),
    .A1(\node_threshold_flat[46] ),
    .S(net540),
    .X(_0912_));
 sg13g2_a221oi_1 _1562_ (.B2(net529),
    .C1(net531),
    .B1(_0912_),
    .A1(\node_threshold_flat[54] ),
    .Y(_0913_),
    .A2(net467));
 sg13g2_a21o_2 _1563_ (.A2(_0911_),
    .A1(_0907_),
    .B1(_0913_),
    .X(_0914_));
 sg13g2_nand2b_1 _1564_ (.Y(_0915_),
    .B(net536),
    .A_N(\node_feature_flat[3] ));
 sg13g2_or2_1 _1565_ (.X(_0916_),
    .B(\node_feature_flat[0] ),
    .A(net536));
 sg13g2_nand3_1 _1566_ (.B(_0915_),
    .C(_0916_),
    .A(net527),
    .Y(_0917_));
 sg13g2_a221oi_1 _1567_ (.B2(\node_feature_flat[9] ),
    .C1(net532),
    .B1(net463),
    .A1(\node_feature_flat[6] ),
    .Y(_0918_),
    .A2(net465));
 sg13g2_mux2_1 _1568_ (.A0(\node_feature_flat[12] ),
    .A1(\node_feature_flat[15] ),
    .S(net537),
    .X(_0919_));
 sg13g2_a221oi_1 _1569_ (.B2(net527),
    .C1(net530),
    .B1(_0919_),
    .A1(\node_feature_flat[18] ),
    .Y(_0920_),
    .A2(net465));
 sg13g2_a21oi_1 _1570_ (.A1(_0917_),
    .A2(_0918_),
    .Y(_0921_),
    .B1(_0920_));
 sg13g2_nand2b_1 _1571_ (.Y(_0922_),
    .B(\feature_vector_flat[38] ),
    .A_N(net447));
 sg13g2_nand2b_1 _1572_ (.Y(_0923_),
    .B(net536),
    .A_N(\node_feature_flat[4] ));
 sg13g2_or2_1 _1573_ (.X(_0924_),
    .B(\node_feature_flat[1] ),
    .A(net536));
 sg13g2_nand3_1 _1574_ (.B(_0923_),
    .C(_0924_),
    .A(net527),
    .Y(_0925_));
 sg13g2_a221oi_1 _1575_ (.B2(\node_feature_flat[10] ),
    .C1(net532),
    .B1(net463),
    .A1(\node_feature_flat[7] ),
    .Y(_0926_),
    .A2(net465));
 sg13g2_mux2_1 _1576_ (.A0(\node_feature_flat[13] ),
    .A1(\node_feature_flat[16] ),
    .S(net537),
    .X(_0927_));
 sg13g2_a221oi_1 _1577_ (.B2(net528),
    .C1(net530),
    .B1(_0927_),
    .A1(\node_feature_flat[19] ),
    .Y(_0928_),
    .A2(net465));
 sg13g2_a21oi_2 _1578_ (.B1(_0928_),
    .Y(_0929_),
    .A2(_0926_),
    .A1(_0925_));
 sg13g2_a21o_1 _1579_ (.A2(_0926_),
    .A1(_0925_),
    .B1(_0928_),
    .X(_0930_));
 sg13g2_a21oi_1 _1580_ (.A1(\feature_vector_flat[46] ),
    .A2(net447),
    .Y(_0931_),
    .B1(_0929_));
 sg13g2_mux2_1 _1581_ (.A0(\node_feature_flat[14] ),
    .A1(\node_feature_flat[17] ),
    .S(net537),
    .X(_0932_));
 sg13g2_a221oi_1 _1582_ (.B2(net527),
    .C1(net530),
    .B1(_0932_),
    .A1(\node_feature_flat[20] ),
    .Y(_0933_),
    .A2(net465));
 sg13g2_nor2_1 _1583_ (.A(net526),
    .B(\node_feature_flat[5] ),
    .Y(_0934_));
 sg13g2_o21ai_1 _1584_ (.B1(net527),
    .Y(_0935_),
    .A1(net536),
    .A2(\node_feature_flat[2] ));
 sg13g2_a221oi_1 _1585_ (.B2(\node_feature_flat[11] ),
    .C1(net532),
    .B1(net463),
    .A1(\node_feature_flat[8] ),
    .Y(_0936_),
    .A2(net465));
 sg13g2_o21ai_1 _1586_ (.B1(_0936_),
    .Y(_0937_),
    .A1(_0934_),
    .A2(_0935_));
 sg13g2_nand2b_2 _1587_ (.Y(_0938_),
    .B(_0937_),
    .A_N(_0933_));
 sg13g2_nand2b_1 _1588_ (.Y(_0939_),
    .B(\feature_vector_flat[54] ),
    .A_N(net447));
 sg13g2_a21oi_1 _1589_ (.A1(\feature_vector_flat[62] ),
    .A2(net447),
    .Y(_0940_),
    .B1(net442));
 sg13g2_a221oi_1 _1590_ (.B2(_0940_),
    .C1(net408),
    .B1(_0939_),
    .A1(_0922_),
    .Y(_0941_),
    .A2(_0931_));
 sg13g2_mux4_1 _1591_ (.S0(net442),
    .A0(\feature_vector_flat[22] ),
    .A1(\feature_vector_flat[6] ),
    .A2(\feature_vector_flat[30] ),
    .A3(\feature_vector_flat[14] ),
    .S1(net447),
    .X(_0942_));
 sg13g2_and2_1 _1592_ (.A(net408),
    .B(_0942_),
    .X(_0943_));
 sg13g2_or3_1 _1593_ (.A(_0914_),
    .B(_0941_),
    .C(_0943_),
    .X(_0944_));
 sg13g2_a21oi_1 _1594_ (.A1(net539),
    .A2(_0846_),
    .Y(_0945_),
    .B1(net534));
 sg13g2_o21ai_1 _1595_ (.B1(_0945_),
    .Y(_0946_),
    .A1(net539),
    .A2(\node_threshold_flat[5] ));
 sg13g2_a221oi_1 _1596_ (.B2(\node_threshold_flat[29] ),
    .C1(net533),
    .B1(net464),
    .A1(\node_threshold_flat[21] ),
    .Y(_0947_),
    .A2(net467));
 sg13g2_mux2_1 _1597_ (.A0(\node_threshold_flat[37] ),
    .A1(\node_threshold_flat[45] ),
    .S(net540),
    .X(_0948_));
 sg13g2_a221oi_1 _1598_ (.B2(net529),
    .C1(net531),
    .B1(_0948_),
    .A1(\node_threshold_flat[53] ),
    .Y(_0949_),
    .A2(net467));
 sg13g2_a21oi_1 _1599_ (.A1(_0946_),
    .A2(_0947_),
    .Y(_0950_),
    .B1(_0949_));
 sg13g2_mux2_1 _1600_ (.A0(\feature_vector_flat[37] ),
    .A1(\feature_vector_flat[45] ),
    .S(net447),
    .X(_0951_));
 sg13g2_or2_1 _1601_ (.X(_0952_),
    .B(net447),
    .A(\feature_vector_flat[53] ));
 sg13g2_a21oi_1 _1602_ (.A1(_0826_),
    .A2(net446),
    .Y(_0953_),
    .B1(net442));
 sg13g2_a221oi_1 _1603_ (.B2(_0953_),
    .C1(net408),
    .B1(_0952_),
    .A1(net443),
    .Y(_0954_),
    .A2(_0951_));
 sg13g2_mux4_1 _1604_ (.S0(net442),
    .A0(\feature_vector_flat[21] ),
    .A1(\feature_vector_flat[5] ),
    .A2(\feature_vector_flat[29] ),
    .A3(\feature_vector_flat[13] ),
    .S1(net446),
    .X(_0955_));
 sg13g2_nor2b_1 _1605_ (.A(_0955_),
    .B_N(net408),
    .Y(_0956_));
 sg13g2_or2_1 _1606_ (.X(_0957_),
    .B(_0956_),
    .A(_0954_));
 sg13g2_o21ai_1 _1607_ (.B1(_0950_),
    .Y(_0958_),
    .A1(_0954_),
    .A2(_0956_));
 sg13g2_and2_1 _1608_ (.A(_0944_),
    .B(_0958_),
    .X(_0959_));
 sg13g2_a21oi_1 _1609_ (.A1(net539),
    .A2(_0844_),
    .Y(_0960_),
    .B1(net534));
 sg13g2_o21ai_1 _1610_ (.B1(_0960_),
    .Y(_0961_),
    .A1(net539),
    .A2(\node_threshold_flat[7] ));
 sg13g2_a221oi_1 _1611_ (.B2(\node_threshold_flat[31] ),
    .C1(net533),
    .B1(net464),
    .A1(\node_threshold_flat[23] ),
    .Y(_0962_),
    .A2(net468));
 sg13g2_mux2_1 _1612_ (.A0(\node_threshold_flat[39] ),
    .A1(\node_threshold_flat[47] ),
    .S(net541),
    .X(_0963_));
 sg13g2_a221oi_1 _1613_ (.B2(net529),
    .C1(net531),
    .B1(_0963_),
    .A1(\node_threshold_flat[55] ),
    .Y(_0964_),
    .A2(net467));
 sg13g2_a21oi_1 _1614_ (.A1(_0961_),
    .A2(_0962_),
    .Y(_0965_),
    .B1(_0964_));
 sg13g2_mux2_1 _1615_ (.A0(\feature_vector_flat[39] ),
    .A1(\feature_vector_flat[47] ),
    .S(net446),
    .X(_0966_));
 sg13g2_or2_1 _1616_ (.X(_0967_),
    .B(net448),
    .A(\feature_vector_flat[55] ));
 sg13g2_a21oi_1 _1617_ (.A1(_0824_),
    .A2(net448),
    .Y(_0968_),
    .B1(net442));
 sg13g2_a221oi_1 _1618_ (.B2(_0968_),
    .C1(net408),
    .B1(_0967_),
    .A1(net443),
    .Y(_0969_),
    .A2(_0966_));
 sg13g2_mux4_1 _1619_ (.S0(net442),
    .A0(\feature_vector_flat[23] ),
    .A1(\feature_vector_flat[7] ),
    .A2(\feature_vector_flat[31] ),
    .A3(\feature_vector_flat[15] ),
    .S1(net448),
    .X(_0970_));
 sg13g2_nor2b_1 _1620_ (.A(_0970_),
    .B_N(net408),
    .Y(_0971_));
 sg13g2_o21ai_1 _1621_ (.B1(_0965_),
    .Y(_0972_),
    .A1(_0969_),
    .A2(_0971_));
 sg13g2_a21oi_1 _1622_ (.A1(net539),
    .A2(_0847_),
    .Y(_0973_),
    .B1(net534));
 sg13g2_o21ai_1 _1623_ (.B1(_0973_),
    .Y(_0974_),
    .A1(net539),
    .A2(\node_threshold_flat[4] ));
 sg13g2_a221oi_1 _1624_ (.B2(\node_threshold_flat[28] ),
    .C1(net533),
    .B1(net464),
    .A1(\node_threshold_flat[20] ),
    .Y(_0975_),
    .A2(net468));
 sg13g2_mux2_1 _1625_ (.A0(\node_threshold_flat[36] ),
    .A1(\node_threshold_flat[44] ),
    .S(net540),
    .X(_0976_));
 sg13g2_a221oi_1 _1626_ (.B2(net529),
    .C1(net531),
    .B1(_0976_),
    .A1(\node_threshold_flat[52] ),
    .Y(_0977_),
    .A2(net467));
 sg13g2_a21o_1 _1627_ (.A2(_0975_),
    .A1(_0974_),
    .B1(_0977_),
    .X(_0978_));
 sg13g2_nand2b_1 _1628_ (.Y(_0979_),
    .B(\feature_vector_flat[36] ),
    .A_N(net446));
 sg13g2_a21oi_1 _1629_ (.A1(\feature_vector_flat[44] ),
    .A2(net446),
    .Y(_0980_),
    .B1(_0929_));
 sg13g2_nand2b_1 _1630_ (.Y(_0981_),
    .B(\feature_vector_flat[52] ),
    .A_N(net446));
 sg13g2_a21oi_1 _1631_ (.A1(\feature_vector_flat[60] ),
    .A2(net446),
    .Y(_0982_),
    .B1(net442));
 sg13g2_a221oi_1 _1632_ (.B2(_0982_),
    .C1(net408),
    .B1(_0981_),
    .A1(_0979_),
    .Y(_0983_),
    .A2(_0980_));
 sg13g2_mux4_1 _1633_ (.S0(net442),
    .A0(\feature_vector_flat[20] ),
    .A1(\feature_vector_flat[4] ),
    .A2(\feature_vector_flat[28] ),
    .A3(\feature_vector_flat[12] ),
    .S1(net446),
    .X(_0984_));
 sg13g2_and2_1 _1634_ (.A(net408),
    .B(_0984_),
    .X(_0985_));
 sg13g2_or3_1 _1635_ (.A(_0978_),
    .B(_0983_),
    .C(_0985_),
    .X(_0986_));
 sg13g2_nand4_1 _1636_ (.B(_0958_),
    .C(_0972_),
    .A(_0944_),
    .Y(_0987_),
    .D(_0986_));
 sg13g2_nor3_1 _1637_ (.A(_0965_),
    .B(_0969_),
    .C(_0971_),
    .Y(_0988_));
 sg13g2_o21ai_1 _1638_ (.B1(_0914_),
    .Y(_0989_),
    .A1(_0941_),
    .A2(_0943_));
 sg13g2_nand2b_1 _1639_ (.Y(_0990_),
    .B(_0989_),
    .A_N(_0988_));
 sg13g2_o21ai_1 _1640_ (.B1(_0978_),
    .Y(_0991_),
    .A1(_0983_),
    .A2(_0985_));
 sg13g2_o21ai_1 _1641_ (.B1(_0991_),
    .Y(_0992_),
    .A1(_0950_),
    .A2(_0957_));
 sg13g2_nor3_1 _1642_ (.A(_0987_),
    .B(_0990_),
    .C(_0992_),
    .Y(_0993_));
 sg13g2_a21oi_1 _1643_ (.A1(net542),
    .A2(_0838_),
    .Y(_0994_),
    .B1(net534));
 sg13g2_o21ai_1 _1644_ (.B1(_0994_),
    .Y(_0995_),
    .A1(net542),
    .A2(\node_threshold_flat[35] ));
 sg13g2_a21oi_1 _1645_ (.A1(\node_threshold_flat[51] ),
    .A2(net467),
    .Y(_0996_),
    .B1(_0820_));
 sg13g2_a21oi_1 _1646_ (.A1(net542),
    .A2(_0848_),
    .Y(_0997_),
    .B1(net534));
 sg13g2_o21ai_1 _1647_ (.B1(_0997_),
    .Y(_0998_),
    .A1(net542),
    .A2(\node_threshold_flat[3] ));
 sg13g2_a221oi_1 _1648_ (.B2(\node_threshold_flat[27] ),
    .C1(net533),
    .B1(net464),
    .A1(\node_threshold_flat[19] ),
    .Y(_0999_),
    .A2(net467));
 sg13g2_a22oi_1 _1649_ (.Y(_1000_),
    .B1(_0998_),
    .B2(_0999_),
    .A2(_0996_),
    .A1(_0995_));
 sg13g2_mux2_1 _1650_ (.A0(\feature_vector_flat[35] ),
    .A1(\feature_vector_flat[43] ),
    .S(net444),
    .X(_1001_));
 sg13g2_or2_1 _1651_ (.X(_1002_),
    .B(net448),
    .A(\feature_vector_flat[51] ));
 sg13g2_a21oi_1 _1652_ (.A1(_0827_),
    .A2(net444),
    .Y(_1003_),
    .B1(net441));
 sg13g2_a221oi_1 _1653_ (.B2(_1003_),
    .C1(net407),
    .B1(_1002_),
    .A1(net443),
    .Y(_1004_),
    .A2(_1001_));
 sg13g2_mux4_1 _1654_ (.S0(net441),
    .A0(\feature_vector_flat[19] ),
    .A1(\feature_vector_flat[3] ),
    .A2(\feature_vector_flat[27] ),
    .A3(\feature_vector_flat[11] ),
    .S1(net444),
    .X(_1005_));
 sg13g2_nor2b_1 _1655_ (.A(_1005_),
    .B_N(net407),
    .Y(_1006_));
 sg13g2_o21ai_1 _1656_ (.B1(_1000_),
    .Y(_1007_),
    .A1(_1004_),
    .A2(_1006_));
 sg13g2_inv_1 _1657_ (.Y(_1008_),
    .A(_1007_));
 sg13g2_nor3_1 _1658_ (.A(_1000_),
    .B(_1004_),
    .C(_1006_),
    .Y(_1009_));
 sg13g2_a21oi_1 _1659_ (.A1(net536),
    .A2(_0849_),
    .Y(_1010_),
    .B1(net535));
 sg13g2_o21ai_1 _1660_ (.B1(_1010_),
    .Y(_1011_),
    .A1(net537),
    .A2(\node_threshold_flat[2] ));
 sg13g2_a221oi_1 _1661_ (.B2(\node_threshold_flat[26] ),
    .C1(net532),
    .B1(net463),
    .A1(\node_threshold_flat[18] ),
    .Y(_1012_),
    .A2(net466));
 sg13g2_mux2_1 _1662_ (.A0(\node_threshold_flat[34] ),
    .A1(\node_threshold_flat[42] ),
    .S(net538),
    .X(_1013_));
 sg13g2_a221oi_1 _1663_ (.B2(net528),
    .C1(net531),
    .B1(_1013_),
    .A1(\node_threshold_flat[50] ),
    .Y(_1014_),
    .A2(net466));
 sg13g2_a21o_1 _1664_ (.A2(_1012_),
    .A1(_1011_),
    .B1(_1014_),
    .X(_1015_));
 sg13g2_nand2b_1 _1665_ (.Y(_1016_),
    .B(\feature_vector_flat[34] ),
    .A_N(net444));
 sg13g2_a21oi_1 _1666_ (.A1(\feature_vector_flat[42] ),
    .A2(net444),
    .Y(_1017_),
    .B1(_0929_));
 sg13g2_nand2b_1 _1667_ (.Y(_1018_),
    .B(\feature_vector_flat[50] ),
    .A_N(net444));
 sg13g2_a21oi_1 _1668_ (.A1(\feature_vector_flat[58] ),
    .A2(net444),
    .Y(_1019_),
    .B1(net443));
 sg13g2_a221oi_1 _1669_ (.B2(_1019_),
    .C1(net407),
    .B1(_1018_),
    .A1(_1016_),
    .Y(_1020_),
    .A2(_1017_));
 sg13g2_mux4_1 _1670_ (.S0(net441),
    .A0(\feature_vector_flat[18] ),
    .A1(\feature_vector_flat[2] ),
    .A2(\feature_vector_flat[26] ),
    .A3(\feature_vector_flat[10] ),
    .S1(net445),
    .X(_1021_));
 sg13g2_and2_1 _1671_ (.A(net407),
    .B(_1021_),
    .X(_1022_));
 sg13g2_or2_1 _1672_ (.X(_1023_),
    .B(_1022_),
    .A(_1020_));
 sg13g2_a21oi_1 _1673_ (.A1(_1015_),
    .A2(_1023_),
    .Y(_1024_),
    .B1(_1009_));
 sg13g2_a21oi_1 _1674_ (.A1(net537),
    .A2(_0850_),
    .Y(_1025_),
    .B1(net535));
 sg13g2_o21ai_1 _1675_ (.B1(_1025_),
    .Y(_1026_),
    .A1(net538),
    .A2(\node_threshold_flat[1] ));
 sg13g2_a221oi_1 _1676_ (.B2(\node_threshold_flat[25] ),
    .C1(net532),
    .B1(net463),
    .A1(\node_threshold_flat[17] ),
    .Y(_1027_),
    .A2(net466));
 sg13g2_mux2_1 _1677_ (.A0(\node_threshold_flat[33] ),
    .A1(\node_threshold_flat[41] ),
    .S(net538),
    .X(_1028_));
 sg13g2_a221oi_1 _1678_ (.B2(net528),
    .C1(net531),
    .B1(_1028_),
    .A1(\node_threshold_flat[49] ),
    .Y(_1029_),
    .A2(net466));
 sg13g2_a21oi_1 _1679_ (.A1(_1026_),
    .A2(_1027_),
    .Y(_1030_),
    .B1(_1029_));
 sg13g2_mux2_1 _1680_ (.A0(\feature_vector_flat[33] ),
    .A1(\feature_vector_flat[41] ),
    .S(net445),
    .X(_1031_));
 sg13g2_or2_1 _1681_ (.X(_1032_),
    .B(net448),
    .A(\feature_vector_flat[49] ));
 sg13g2_a21oi_1 _1682_ (.A1(_0828_),
    .A2(net445),
    .Y(_1033_),
    .B1(net441));
 sg13g2_a221oi_1 _1683_ (.B2(_1033_),
    .C1(net407),
    .B1(_1032_),
    .A1(net441),
    .Y(_1034_),
    .A2(_1031_));
 sg13g2_mux4_1 _1684_ (.S0(net441),
    .A0(\feature_vector_flat[17] ),
    .A1(\feature_vector_flat[1] ),
    .A2(\feature_vector_flat[25] ),
    .A3(\feature_vector_flat[9] ),
    .S1(net445),
    .X(_1035_));
 sg13g2_nor2b_1 _1685_ (.A(_1035_),
    .B_N(net407),
    .Y(_1036_));
 sg13g2_nor3_1 _1686_ (.A(_1030_),
    .B(_1034_),
    .C(_1036_),
    .Y(_1037_));
 sg13g2_or3_1 _1687_ (.A(_1015_),
    .B(_1020_),
    .C(_1022_),
    .X(_1038_));
 sg13g2_nand2_1 _1688_ (.Y(_1039_),
    .A(_1037_),
    .B(_1038_));
 sg13g2_a21oi_1 _1689_ (.A1(_1024_),
    .A2(_1039_),
    .Y(_1040_),
    .B1(_1008_));
 sg13g2_a21o_1 _1690_ (.A2(_0992_),
    .A1(_0959_),
    .B1(_0990_),
    .X(_1041_));
 sg13g2_mux2_1 _1691_ (.A0(\node_threshold_flat[32] ),
    .A1(\node_threshold_flat[40] ),
    .S(net537),
    .X(_1042_));
 sg13g2_a221oi_1 _1692_ (.B2(net528),
    .C1(net531),
    .B1(_1042_),
    .A1(\node_threshold_flat[48] ),
    .Y(_1043_),
    .A2(net466));
 sg13g2_a21oi_1 _1693_ (.A1(net536),
    .A2(_0851_),
    .Y(_1044_),
    .B1(net535));
 sg13g2_o21ai_1 _1694_ (.B1(_1044_),
    .Y(_1045_),
    .A1(net537),
    .A2(\node_threshold_flat[0] ));
 sg13g2_a221oi_1 _1695_ (.B2(\node_threshold_flat[24] ),
    .C1(net533),
    .B1(net464),
    .A1(\node_threshold_flat[16] ),
    .Y(_1046_),
    .A2(net466));
 sg13g2_a21oi_1 _1696_ (.A1(_1045_),
    .A2(_1046_),
    .Y(_1047_),
    .B1(_1043_));
 sg13g2_nand2b_1 _1697_ (.Y(_1048_),
    .B(\feature_vector_flat[32] ),
    .A_N(net445));
 sg13g2_a21oi_1 _1698_ (.A1(\feature_vector_flat[40] ),
    .A2(net445),
    .Y(_1049_),
    .B1(_0929_));
 sg13g2_nand2b_1 _1699_ (.Y(_1050_),
    .B(\feature_vector_flat[48] ),
    .A_N(net444));
 sg13g2_a21oi_1 _1700_ (.A1(\feature_vector_flat[56] ),
    .A2(net445),
    .Y(_1051_),
    .B1(net441));
 sg13g2_a221oi_1 _1701_ (.B2(_1051_),
    .C1(net407),
    .B1(_1050_),
    .A1(_1048_),
    .Y(_1052_),
    .A2(_1049_));
 sg13g2_mux4_1 _1702_ (.S0(net441),
    .A0(\feature_vector_flat[16] ),
    .A1(\feature_vector_flat[0] ),
    .A2(\feature_vector_flat[24] ),
    .A3(\feature_vector_flat[8] ),
    .S1(net445),
    .X(_1053_));
 sg13g2_nand2_1 _1703_ (.Y(_1054_),
    .A(net407),
    .B(_1053_));
 sg13g2_nor2b_1 _1704_ (.A(_1052_),
    .B_N(_1054_),
    .Y(_1055_));
 sg13g2_nand3b_1 _1705_ (.B(_1054_),
    .C(_1047_),
    .Y(_1056_),
    .A_N(_1052_));
 sg13g2_o21ai_1 _1706_ (.B1(_1030_),
    .Y(_1057_),
    .A1(_1034_),
    .A2(_1036_));
 sg13g2_nand4_1 _1707_ (.B(_1038_),
    .C(_1056_),
    .A(_1007_),
    .Y(_1058_),
    .D(_1057_));
 sg13g2_nor4_1 _1708_ (.A(_0987_),
    .B(_0990_),
    .C(_0992_),
    .D(_1058_),
    .Y(_1059_));
 sg13g2_a221oi_1 _1709_ (.B2(_0972_),
    .C1(_1059_),
    .B1(_1041_),
    .A1(_0993_),
    .Y(_1060_),
    .A2(_1040_));
 sg13g2_nor2_1 _1710_ (.A(_1047_),
    .B(_1055_),
    .Y(_1061_));
 sg13g2_nor2_1 _1711_ (.A(_1037_),
    .B(_1061_),
    .Y(_1062_));
 sg13g2_and3_2 _1712_ (.X(_1063_),
    .A(_1024_),
    .B(_1059_),
    .C(_1062_));
 sg13g2_nor2_1 _1713_ (.A(_1060_),
    .B(_1063_),
    .Y(_1064_));
 sg13g2_mux4_1 _1714_ (.S0(net526),
    .A0(\node_left_flat[7] ),
    .A1(\node_left_flat[3] ),
    .A2(\node_right_flat[7] ),
    .A3(\node_right_flat[3] ),
    .S1(net383),
    .X(_1065_));
 sg13g2_mux2_1 _1715_ (.A0(_0860_),
    .A1(_0874_),
    .S(net384),
    .X(_1066_));
 sg13g2_o21ai_1 _1716_ (.B1(\node_left_flat[11] ),
    .Y(_1067_),
    .A1(_1060_),
    .A2(_1063_));
 sg13g2_a21oi_1 _1717_ (.A1(\node_right_flat[11] ),
    .A2(net384),
    .Y(_1068_),
    .B1(_0909_));
 sg13g2_a22oi_1 _1718_ (.Y(_1069_),
    .B1(_1067_),
    .B2(_1068_),
    .A2(_1066_),
    .A1(net463));
 sg13g2_o21ai_1 _1719_ (.B1(_1069_),
    .Y(_1070_),
    .A1(net535),
    .A2(_1065_));
 sg13g2_mux4_1 _1720_ (.S0(net526),
    .A0(\node_left_flat[23] ),
    .A1(\node_left_flat[19] ),
    .A2(\node_right_flat[23] ),
    .A3(\node_right_flat[19] ),
    .S1(net383),
    .X(_1071_));
 sg13g2_nor2_1 _1721_ (.A(\node_left_flat[27] ),
    .B(net385),
    .Y(_1072_));
 sg13g2_a21oi_1 _1722_ (.A1(_0869_),
    .A2(net385),
    .Y(_1073_),
    .B1(_1072_));
 sg13g2_a221oi_1 _1723_ (.B2(net465),
    .C1(net530),
    .B1(_1073_),
    .A1(net527),
    .Y(_1074_),
    .A2(_1071_));
 sg13g2_a21oi_2 _1724_ (.B1(_1074_),
    .Y(_1075_),
    .A2(_1070_),
    .A1(net530));
 sg13g2_mux4_1 _1725_ (.S0(net526),
    .A0(\node_left_flat[6] ),
    .A1(\node_left_flat[2] ),
    .A2(\node_right_flat[6] ),
    .A3(\node_right_flat[2] ),
    .S1(net383),
    .X(_1076_));
 sg13g2_or2_1 _1726_ (.X(_1077_),
    .B(_1076_),
    .A(net535));
 sg13g2_mux2_1 _1727_ (.A0(_0861_),
    .A1(_0875_),
    .S(net384),
    .X(_1078_));
 sg13g2_o21ai_1 _1728_ (.B1(\node_left_flat[10] ),
    .Y(_1079_),
    .A1(_1060_),
    .A2(_1063_));
 sg13g2_a21oi_1 _1729_ (.A1(\node_right_flat[10] ),
    .A2(net384),
    .Y(_1080_),
    .B1(_0909_));
 sg13g2_a22oi_1 _1730_ (.Y(_1081_),
    .B1(_1079_),
    .B2(_1080_),
    .A2(_1078_),
    .A1(net463));
 sg13g2_a21oi_1 _1731_ (.A1(_1077_),
    .A2(_1081_),
    .Y(_1082_),
    .B1(net532));
 sg13g2_mux4_1 _1732_ (.S0(net526),
    .A0(\node_left_flat[22] ),
    .A1(\node_left_flat[18] ),
    .A2(\node_right_flat[22] ),
    .A3(\node_right_flat[18] ),
    .S1(net383),
    .X(_1083_));
 sg13g2_or2_1 _1733_ (.X(_1084_),
    .B(net385),
    .A(\node_left_flat[26] ));
 sg13g2_a21oi_1 _1734_ (.A1(_0870_),
    .A2(net385),
    .Y(_1085_),
    .B1(_0909_));
 sg13g2_a221oi_1 _1735_ (.B2(_1085_),
    .C1(net530),
    .B1(_1084_),
    .A1(net527),
    .Y(_1086_),
    .A2(_1083_));
 sg13g2_nor2_2 _1736_ (.A(_1082_),
    .B(_1086_),
    .Y(_1087_));
 sg13g2_or2_1 _1737_ (.X(_1088_),
    .B(_1086_),
    .A(_1082_));
 sg13g2_mux4_1 _1738_ (.S0(net526),
    .A0(\node_left_flat[5] ),
    .A1(\node_left_flat[1] ),
    .A2(\node_right_flat[5] ),
    .A3(\node_right_flat[1] ),
    .S1(net383),
    .X(_1089_));
 sg13g2_or2_1 _1739_ (.X(_1090_),
    .B(_1089_),
    .A(net535));
 sg13g2_mux2_1 _1740_ (.A0(_0862_),
    .A1(_0876_),
    .S(net384),
    .X(_1091_));
 sg13g2_o21ai_1 _1741_ (.B1(\node_left_flat[9] ),
    .Y(_1092_),
    .A1(_1060_),
    .A2(_1063_));
 sg13g2_a21oi_1 _1742_ (.A1(\node_right_flat[9] ),
    .A2(net384),
    .Y(_1093_),
    .B1(_0909_));
 sg13g2_a22oi_1 _1743_ (.Y(_1094_),
    .B1(_1092_),
    .B2(_1093_),
    .A2(_1091_),
    .A1(net463));
 sg13g2_a21o_2 _1744_ (.A2(_1094_),
    .A1(_1090_),
    .B1(net532),
    .X(_1095_));
 sg13g2_mux4_1 _1745_ (.S0(net526),
    .A0(\node_left_flat[21] ),
    .A1(\node_left_flat[17] ),
    .A2(\node_right_flat[21] ),
    .A3(\node_right_flat[17] ),
    .S1(net383),
    .X(_1096_));
 sg13g2_nor3_1 _1746_ (.A(\node_right_flat[25] ),
    .B(_1060_),
    .C(_1063_),
    .Y(_1097_));
 sg13g2_o21ai_1 _1747_ (.B1(net465),
    .Y(_1098_),
    .A1(\node_left_flat[25] ),
    .A2(net385));
 sg13g2_o21ai_1 _1748_ (.B1(net532),
    .Y(_1099_),
    .A1(_1097_),
    .A2(_1098_));
 sg13g2_a21o_2 _1749_ (.A2(_1096_),
    .A1(net528),
    .B1(_1099_),
    .X(_1100_));
 sg13g2_nand2_2 _1750_ (.Y(_1101_),
    .A(_1095_),
    .B(_1100_));
 sg13g2_mux2_1 _1751_ (.A0(_0866_),
    .A1(_0880_),
    .S(net383),
    .X(_1102_));
 sg13g2_mux2_1 _1752_ (.A0(_0868_),
    .A1(_0882_),
    .S(net383),
    .X(_1103_));
 sg13g2_mux2_1 _1753_ (.A0(_0863_),
    .A1(_0877_),
    .S(net384),
    .X(_1104_));
 sg13g2_mux2_1 _1754_ (.A0(_0864_),
    .A1(_0878_),
    .S(net384),
    .X(_1105_));
 sg13g2_mux4_1 _1755_ (.S0(_0822_),
    .A0(_1102_),
    .A1(_1103_),
    .A2(_1104_),
    .A3(_1105_),
    .S1(net535),
    .X(_1106_));
 sg13g2_mux4_1 _1756_ (.S0(net526),
    .A0(\node_left_flat[20] ),
    .A1(\node_left_flat[16] ),
    .A2(\node_right_flat[20] ),
    .A3(\node_right_flat[16] ),
    .S1(net386),
    .X(_1107_));
 sg13g2_or2_1 _1757_ (.X(_1108_),
    .B(net385),
    .A(\node_left_flat[24] ));
 sg13g2_a21oi_1 _1758_ (.A1(_0871_),
    .A2(net385),
    .Y(_1109_),
    .B1(_0909_));
 sg13g2_a221oi_1 _1759_ (.B2(_1109_),
    .C1(net530),
    .B1(_1108_),
    .A1(net527),
    .Y(_1110_),
    .A2(_1107_));
 sg13g2_a21oi_1 _1760_ (.A1(net530),
    .A2(_1106_),
    .Y(_1111_),
    .B1(_1110_));
 sg13g2_and3_2 _1761_ (.X(_1112_),
    .A(_1095_),
    .B(_1100_),
    .C(net380));
 sg13g2_a21o_2 _1762_ (.A2(_1112_),
    .A1(_1087_),
    .B1(_1075_),
    .X(_1113_));
 sg13g2_nor2b_2 _1763_ (.A(net1041),
    .B_N(net593),
    .Y(_1114_));
 sg13g2_nand2b_2 _1764_ (.Y(_1115_),
    .B(net1078),
    .A_N(_1114_));
 sg13g2_or2_1 _1765_ (.X(_1116_),
    .B(_1115_),
    .A(_1113_));
 sg13g2_nand2_1 _1766_ (.Y(_1117_),
    .A(net920),
    .B(net1019));
 sg13g2_nand4_1 _1767_ (.B(net1053),
    .C(net1061),
    .A(net920),
    .Y(_1118_),
    .D(net1019));
 sg13g2_a21oi_1 _1768_ (.A1(_1116_),
    .A2(_1118_),
    .Y(_0001_),
    .B1(net485));
 sg13g2_nor2_1 _1769_ (.A(net485),
    .B(_1115_),
    .Y(_1119_));
 sg13g2_and2_1 _1770_ (.A(\u_tree_core.state_q[1] ),
    .B(_1114_),
    .X(_1120_));
 sg13g2_nand2b_1 _1771_ (.Y(_1121_),
    .B(net1053),
    .A_N(run_cmd));
 sg13g2_nand2_1 _1772_ (.Y(_1122_),
    .A(net509),
    .B(_1121_));
 sg13g2_a221oi_1 _1773_ (.B2(_1113_),
    .C1(_1122_),
    .B1(_1119_),
    .A1(net1053),
    .Y(_1123_),
    .A2(_1117_));
 sg13g2_nand2b_1 _1774_ (.Y(_0000_),
    .B(net1054),
    .A_N(_1120_));
 sg13g2_nand2_2 _1775_ (.Y(uio_out[7]),
    .A(_0823_),
    .B(features_loaded));
 sg13g2_nand3_1 _1776_ (.B(net1),
    .C(net10),
    .A(io_ready),
    .Y(_1124_));
 sg13g2_nor2_1 _1777_ (.A(net11),
    .B(_1124_),
    .Y(_1125_));
 sg13g2_and4_1 _1778_ (.A(net2),
    .B(net553),
    .C(net12),
    .D(_1125_),
    .X(_0002_));
 sg13g2_nor3_2 _1779_ (.A(_0903_),
    .B(net12),
    .C(_1124_),
    .Y(_1126_));
 sg13g2_and2_1 _1780_ (.A(net554),
    .B(net440),
    .X(_0003_));
 sg13g2_o21ai_1 _1781_ (.B1(net554),
    .Y(_1127_),
    .A1(net1065),
    .A2(net439));
 sg13g2_a21oi_1 _1782_ (.A1(_0901_),
    .A2(net439),
    .Y(_0004_),
    .B1(_1127_));
 sg13g2_o21ai_1 _1783_ (.B1(net555),
    .Y(_1128_),
    .A1(net1071),
    .A2(net440));
 sg13g2_a21oi_1 _1784_ (.A1(_0899_),
    .A2(net440),
    .Y(_0005_),
    .B1(_1128_));
 sg13g2_o21ai_1 _1785_ (.B1(net555),
    .Y(_1129_),
    .A1(net1066),
    .A2(net439));
 sg13g2_a21oi_1 _1786_ (.A1(_0897_),
    .A2(net440),
    .Y(_0006_),
    .B1(_1129_));
 sg13g2_o21ai_1 _1787_ (.B1(net555),
    .Y(_1130_),
    .A1(net1069),
    .A2(net440));
 sg13g2_a21oi_1 _1788_ (.A1(_0895_),
    .A2(_1126_),
    .Y(_0007_),
    .B1(_1130_));
 sg13g2_o21ai_1 _1789_ (.B1(net554),
    .Y(_1131_),
    .A1(net1058),
    .A2(net439));
 sg13g2_a21oi_1 _1790_ (.A1(_0893_),
    .A2(net439),
    .Y(_0008_),
    .B1(_1131_));
 sg13g2_o21ai_1 _1791_ (.B1(net555),
    .Y(_1132_),
    .A1(net1064),
    .A2(net440));
 sg13g2_a21oi_1 _1792_ (.A1(_0891_),
    .A2(net440),
    .Y(_0009_),
    .B1(_1132_));
 sg13g2_o21ai_1 _1793_ (.B1(net554),
    .Y(_1133_),
    .A1(net1052),
    .A2(net439));
 sg13g2_a21oi_1 _1794_ (.A1(_0889_),
    .A2(net439),
    .Y(_0010_),
    .B1(_1133_));
 sg13g2_o21ai_1 _1795_ (.B1(net554),
    .Y(_1134_),
    .A1(net1050),
    .A2(_1126_));
 sg13g2_a21oi_1 _1796_ (.A1(_0887_),
    .A2(net439),
    .Y(_0011_),
    .B1(_1134_));
 sg13g2_nor3_2 _1797_ (.A(net11),
    .B(net12),
    .C(_1124_),
    .Y(_1135_));
 sg13g2_and2_1 _1798_ (.A(net553),
    .B(net438),
    .X(_0012_));
 sg13g2_o21ai_1 _1799_ (.B1(net553),
    .Y(_1136_),
    .A1(net1047),
    .A2(net438));
 sg13g2_a21oi_1 _1800_ (.A1(_0901_),
    .A2(net438),
    .Y(_0013_),
    .B1(_1136_));
 sg13g2_o21ai_1 _1801_ (.B1(net553),
    .Y(_1137_),
    .A1(net1048),
    .A2(net437));
 sg13g2_a21oi_1 _1802_ (.A1(_0899_),
    .A2(_1135_),
    .Y(_0014_),
    .B1(_1137_));
 sg13g2_o21ai_1 _1803_ (.B1(net556),
    .Y(_1138_),
    .A1(net1049),
    .A2(net437));
 sg13g2_a21oi_1 _1804_ (.A1(_0897_),
    .A2(net437),
    .Y(_0015_),
    .B1(_1138_));
 sg13g2_o21ai_1 _1805_ (.B1(net553),
    .Y(_1139_),
    .A1(net549),
    .A2(net437));
 sg13g2_a21oi_1 _1806_ (.A1(_0895_),
    .A2(net438),
    .Y(_0016_),
    .B1(_1139_));
 sg13g2_o21ai_1 _1807_ (.B1(net553),
    .Y(_1140_),
    .A1(net1051),
    .A2(net437));
 sg13g2_a21oi_1 _1808_ (.A1(_0893_),
    .A2(net437),
    .Y(_0017_),
    .B1(_1140_));
 sg13g2_o21ai_1 _1809_ (.B1(net556),
    .Y(_1141_),
    .A1(net1059),
    .A2(net437));
 sg13g2_a21oi_1 _1810_ (.A1(_0891_),
    .A2(net437),
    .Y(_0018_),
    .B1(_1141_));
 sg13g2_o21ai_1 _1811_ (.B1(net553),
    .Y(_1142_),
    .A1(net1060),
    .A2(net438));
 sg13g2_a21oi_1 _1812_ (.A1(_0889_),
    .A2(_1135_),
    .Y(_0019_),
    .B1(_1142_));
 sg13g2_o21ai_1 _1813_ (.B1(net553),
    .Y(_1143_),
    .A1(net1063),
    .A2(net438));
 sg13g2_a21oi_1 _1814_ (.A1(_0887_),
    .A2(net438),
    .Y(_0020_),
    .B1(_1143_));
 sg13g2_and2_1 _1815_ (.A(\u_feature_loader.feature_idx_q[1] ),
    .B(\u_feature_loader.feature_idx_q[0] ),
    .X(_1144_));
 sg13g2_and2_1 _1816_ (.A(net586),
    .B(_1144_),
    .X(_1145_));
 sg13g2_nand2_1 _1817_ (.Y(_1146_),
    .A(net544),
    .B(_1145_));
 sg13g2_or2_1 _1818_ (.X(_1147_),
    .B(_1146_),
    .A(net643));
 sg13g2_nor3_2 _1819_ (.A(net544),
    .B(\u_feature_loader.feature_idx_q[1] ),
    .C(\u_feature_loader.feature_idx_q[0] ),
    .Y(_1148_));
 sg13g2_nor2_1 _1820_ (.A(_0825_),
    .B(\u_feature_loader.feature_idx_q[3] ),
    .Y(_1149_));
 sg13g2_nand2b_2 _1821_ (.Y(_1150_),
    .B(_1148_),
    .A_N(\u_feature_loader.feature_idx_q[3] ));
 sg13g2_nand2_2 _1822_ (.Y(_1151_),
    .A(_1148_),
    .B(_1149_));
 sg13g2_nand3b_1 _1823_ (.B(net1019),
    .C(_1151_),
    .Y(_1152_),
    .A_N(run_cmd));
 sg13g2_a21oi_1 _1824_ (.A1(net406),
    .A2(net1020),
    .Y(_0021_),
    .B1(net491));
 sg13g2_a21o_1 _1825_ (.A2(_1113_),
    .A1(\u_tree_core.state_q[1] ),
    .B1(_1120_),
    .X(_1153_));
 sg13g2_nand2_1 _1826_ (.Y(_1154_),
    .A(net508),
    .B(net377));
 sg13g2_inv_1 _1827_ (.Y(_0022_),
    .A(net376));
 sg13g2_o21ai_1 _1828_ (.B1(net494),
    .Y(_1155_),
    .A1(model_byte_valid),
    .A2(net547));
 sg13g2_a21oi_1 _1829_ (.A1(model_byte_valid),
    .A2(net561),
    .Y(_0023_),
    .B1(_1155_));
 sg13g2_a21oi_1 _1830_ (.A1(model_byte_valid),
    .A2(net547),
    .Y(_1156_),
    .B1(net880));
 sg13g2_nand2_1 _1831_ (.Y(_0311_),
    .A(\u_model_loader.byte_idx_q[1] ),
    .B(net547));
 sg13g2_and3_2 _1832_ (.X(_0312_),
    .A(model_byte_valid),
    .B(net880),
    .C(net547));
 sg13g2_nand3_1 _1833_ (.B(net880),
    .C(net547),
    .A(model_byte_valid),
    .Y(_0313_));
 sg13g2_nor3_1 _1834_ (.A(net474),
    .B(net881),
    .C(_0312_),
    .Y(_0024_));
 sg13g2_nand2b_2 _1835_ (.Y(_0314_),
    .B(model_byte_valid),
    .A_N(\u_model_loader.byte_idx_q[5] ));
 sg13g2_nor2_1 _1836_ (.A(\u_model_loader.byte_idx_q[3] ),
    .B(\u_model_loader.byte_idx_q[2] ),
    .Y(_0315_));
 sg13g2_nand2_2 _1837_ (.Y(_0316_),
    .A(net1036),
    .B(net1056));
 sg13g2_nand3_1 _1838_ (.B(\u_model_loader.byte_idx_q[3] ),
    .C(\u_model_loader.byte_idx_q[2] ),
    .A(net545),
    .Y(_0317_));
 sg13g2_nand2b_2 _1839_ (.Y(_0318_),
    .B(_0317_),
    .A_N(\u_model_loader.byte_idx_q[5] ));
 sg13g2_nor3_2 _1840_ (.A(net545),
    .B(\u_model_loader.byte_idx_q[3] ),
    .C(\u_model_loader.byte_idx_q[2] ),
    .Y(_0319_));
 sg13g2_nand2b_1 _1841_ (.Y(_0320_),
    .B(_0315_),
    .A_N(net546));
 sg13g2_xor2_1 _1842_ (.B(_0315_),
    .A(net546),
    .X(_0321_));
 sg13g2_nand2_1 _1843_ (.Y(_0322_),
    .A(\u_model_loader.byte_idx_q[5] ),
    .B(net545));
 sg13g2_nand4_1 _1844_ (.B(_0318_),
    .C(_0321_),
    .A(model_byte_valid),
    .Y(_0323_),
    .D(_0322_));
 sg13g2_nand2b_2 _1845_ (.Y(_0324_),
    .B(_0885_),
    .A_N(_0323_));
 sg13g2_nor2_2 _1846_ (.A(_0311_),
    .B(_0324_),
    .Y(_0325_));
 sg13g2_xnor2_1 _1847_ (.Y(_0326_),
    .A(net1056),
    .B(_0312_));
 sg13g2_nor3_1 _1848_ (.A(net474),
    .B(net402),
    .C(net1057),
    .Y(_0025_));
 sg13g2_a21oi_1 _1849_ (.A1(\u_model_loader.byte_idx_q[2] ),
    .A2(_0312_),
    .Y(_0327_),
    .B1(net1036));
 sg13g2_nor2_2 _1850_ (.A(_0313_),
    .B(_0316_),
    .Y(_0328_));
 sg13g2_nor3_1 _1851_ (.A(net474),
    .B(net1037),
    .C(_0328_),
    .Y(_0026_));
 sg13g2_nor2_1 _1852_ (.A(net545),
    .B(_0328_),
    .Y(_0329_));
 sg13g2_nor2_1 _1853_ (.A(_0313_),
    .B(_0317_),
    .Y(_0330_));
 sg13g2_nor3_1 _1854_ (.A(net474),
    .B(net1073),
    .C(_0330_),
    .Y(_0027_));
 sg13g2_xnor2_1 _1855_ (.Y(_0331_),
    .A(net972),
    .B(_0330_));
 sg13g2_nor3_1 _1856_ (.A(net474),
    .B(net402),
    .C(net973),
    .Y(_0028_));
 sg13g2_or2_1 _1857_ (.X(_0332_),
    .B(_0323_),
    .A(_0885_));
 sg13g2_nor2_1 _1858_ (.A(\u_model_loader.byte_idx_q[1] ),
    .B(net547),
    .Y(_0333_));
 sg13g2_nor2b_2 _1859_ (.A(_0332_),
    .B_N(_0333_),
    .Y(_0334_));
 sg13g2_o21ai_1 _1860_ (.B1(net502),
    .Y(_0335_),
    .A1(net966),
    .A2(net399));
 sg13g2_a21oi_1 _1861_ (.A1(net517),
    .A2(net399),
    .Y(_0029_),
    .B1(_0335_));
 sg13g2_o21ai_1 _1862_ (.B1(net500),
    .Y(_0336_),
    .A1(net968),
    .A2(net399));
 sg13g2_a21oi_1 _1863_ (.A1(net519),
    .A2(net399),
    .Y(_0030_),
    .B1(_0336_));
 sg13g2_o21ai_1 _1864_ (.B1(net493),
    .Y(_0337_),
    .A1(net926),
    .A2(net399));
 sg13g2_a21oi_1 _1865_ (.A1(net520),
    .A2(net399),
    .Y(_0031_),
    .B1(_0337_));
 sg13g2_o21ai_1 _1866_ (.B1(net500),
    .Y(_0338_),
    .A1(net944),
    .A2(net399));
 sg13g2_a21oi_1 _1867_ (.A1(net521),
    .A2(net399),
    .Y(_0032_),
    .B1(_0338_));
 sg13g2_o21ai_1 _1868_ (.B1(net505),
    .Y(_0339_),
    .A1(net865),
    .A2(net400));
 sg13g2_a21oi_1 _1869_ (.A1(net522),
    .A2(net400),
    .Y(_0033_),
    .B1(_0339_));
 sg13g2_o21ai_1 _1870_ (.B1(net505),
    .Y(_0340_),
    .A1(net890),
    .A2(net400));
 sg13g2_a21oi_1 _1871_ (.A1(net523),
    .A2(net400),
    .Y(_0034_),
    .B1(_0340_));
 sg13g2_o21ai_1 _1872_ (.B1(net507),
    .Y(_0341_),
    .A1(net856),
    .A2(net400));
 sg13g2_a21oi_1 _1873_ (.A1(net524),
    .A2(net400),
    .Y(_0035_),
    .B1(_0341_));
 sg13g2_o21ai_1 _1874_ (.B1(net502),
    .Y(_0342_),
    .A1(net980),
    .A2(net400));
 sg13g2_a21oi_1 _1875_ (.A1(net525),
    .A2(net400),
    .Y(_0036_),
    .B1(_0342_));
 sg13g2_nand2b_2 _1876_ (.Y(_0343_),
    .B(net547),
    .A_N(\u_model_loader.byte_idx_q[1] ));
 sg13g2_nor2_2 _1877_ (.A(_0332_),
    .B(_0343_),
    .Y(_0344_));
 sg13g2_o21ai_1 _1878_ (.B1(net502),
    .Y(_0345_),
    .A1(net914),
    .A2(net397));
 sg13g2_a21oi_1 _1879_ (.A1(net517),
    .A2(net397),
    .Y(_0037_),
    .B1(_0345_));
 sg13g2_o21ai_1 _1880_ (.B1(net500),
    .Y(_0346_),
    .A1(net1015),
    .A2(net397));
 sg13g2_a21oi_1 _1881_ (.A1(net519),
    .A2(net397),
    .Y(_0038_),
    .B1(_0346_));
 sg13g2_o21ai_1 _1882_ (.B1(net493),
    .Y(_0347_),
    .A1(net852),
    .A2(net397));
 sg13g2_a21oi_1 _1883_ (.A1(net520),
    .A2(net397),
    .Y(_0039_),
    .B1(_0347_));
 sg13g2_o21ai_1 _1884_ (.B1(net501),
    .Y(_0348_),
    .A1(net945),
    .A2(net397));
 sg13g2_a21oi_1 _1885_ (.A1(net521),
    .A2(net397),
    .Y(_0040_),
    .B1(_0348_));
 sg13g2_o21ai_1 _1886_ (.B1(net505),
    .Y(_0349_),
    .A1(net1002),
    .A2(net398));
 sg13g2_a21oi_1 _1887_ (.A1(net522),
    .A2(net398),
    .Y(_0041_),
    .B1(_0349_));
 sg13g2_o21ai_1 _1888_ (.B1(net505),
    .Y(_0350_),
    .A1(net1034),
    .A2(net398));
 sg13g2_a21oi_1 _1889_ (.A1(net523),
    .A2(net398),
    .Y(_0042_),
    .B1(_0350_));
 sg13g2_o21ai_1 _1890_ (.B1(net507),
    .Y(_0351_),
    .A1(net824),
    .A2(net398));
 sg13g2_a21oi_1 _1891_ (.A1(net524),
    .A2(net398),
    .Y(_0043_),
    .B1(_0351_));
 sg13g2_o21ai_1 _1892_ (.B1(net502),
    .Y(_0352_),
    .A1(net872),
    .A2(net398));
 sg13g2_a21oi_1 _1893_ (.A1(net525),
    .A2(net398),
    .Y(_0044_),
    .B1(_0352_));
 sg13g2_nand2b_2 _1894_ (.Y(_0353_),
    .B(net880),
    .A_N(net547));
 sg13g2_nor2_2 _1895_ (.A(_0332_),
    .B(_0353_),
    .Y(_0354_));
 sg13g2_o21ai_1 _1896_ (.B1(net502),
    .Y(_0355_),
    .A1(net1009),
    .A2(net395));
 sg13g2_a21oi_1 _1897_ (.A1(net517),
    .A2(net395),
    .Y(_0045_),
    .B1(_0355_));
 sg13g2_o21ai_1 _1898_ (.B1(net493),
    .Y(_0356_),
    .A1(net934),
    .A2(net395));
 sg13g2_a21oi_1 _1899_ (.A1(net519),
    .A2(net395),
    .Y(_0046_),
    .B1(_0356_));
 sg13g2_o21ai_1 _1900_ (.B1(net493),
    .Y(_0357_),
    .A1(net860),
    .A2(net395));
 sg13g2_a21oi_1 _1901_ (.A1(net520),
    .A2(net395),
    .Y(_0047_),
    .B1(_0357_));
 sg13g2_o21ai_1 _1902_ (.B1(net500),
    .Y(_0358_),
    .A1(net949),
    .A2(net395));
 sg13g2_a21oi_1 _1903_ (.A1(net521),
    .A2(net395),
    .Y(_0048_),
    .B1(_0358_));
 sg13g2_o21ai_1 _1904_ (.B1(net505),
    .Y(_0359_),
    .A1(net956),
    .A2(net396));
 sg13g2_a21oi_1 _1905_ (.A1(net522),
    .A2(net396),
    .Y(_0049_),
    .B1(_0359_));
 sg13g2_o21ai_1 _1906_ (.B1(net505),
    .Y(_0360_),
    .A1(net901),
    .A2(net396));
 sg13g2_a21oi_1 _1907_ (.A1(net523),
    .A2(net396),
    .Y(_0050_),
    .B1(_0360_));
 sg13g2_o21ai_1 _1908_ (.B1(net507),
    .Y(_0361_),
    .A1(net938),
    .A2(net396));
 sg13g2_a21oi_1 _1909_ (.A1(net524),
    .A2(net396),
    .Y(_0051_),
    .B1(_0361_));
 sg13g2_o21ai_1 _1910_ (.B1(net503),
    .Y(_0362_),
    .A1(net1039),
    .A2(net396));
 sg13g2_a21oi_1 _1911_ (.A1(net525),
    .A2(net396),
    .Y(_0052_),
    .B1(_0362_));
 sg13g2_nor2_2 _1912_ (.A(_0311_),
    .B(_0332_),
    .Y(_0363_));
 sg13g2_o21ai_1 _1913_ (.B1(net502),
    .Y(_0364_),
    .A1(net1024),
    .A2(net393));
 sg13g2_a21oi_1 _1914_ (.A1(net517),
    .A2(net393),
    .Y(_0053_),
    .B1(_0364_));
 sg13g2_o21ai_1 _1915_ (.B1(net500),
    .Y(_0365_),
    .A1(net1022),
    .A2(net393));
 sg13g2_a21oi_1 _1916_ (.A1(net519),
    .A2(net393),
    .Y(_0054_),
    .B1(_0365_));
 sg13g2_o21ai_1 _1917_ (.B1(net493),
    .Y(_0366_),
    .A1(net962),
    .A2(net393));
 sg13g2_a21oi_1 _1918_ (.A1(net520),
    .A2(net393),
    .Y(_0055_),
    .B1(_0366_));
 sg13g2_o21ai_1 _1919_ (.B1(net500),
    .Y(_0367_),
    .A1(net883),
    .A2(net393));
 sg13g2_a21oi_1 _1920_ (.A1(net521),
    .A2(net393),
    .Y(_0056_),
    .B1(_0367_));
 sg13g2_o21ai_1 _1921_ (.B1(net505),
    .Y(_0368_),
    .A1(net822),
    .A2(net394));
 sg13g2_a21oi_1 _1922_ (.A1(net522),
    .A2(net394),
    .Y(_0057_),
    .B1(_0368_));
 sg13g2_o21ai_1 _1923_ (.B1(net505),
    .Y(_0369_),
    .A1(net1017),
    .A2(net394));
 sg13g2_a21oi_1 _1924_ (.A1(net523),
    .A2(net394),
    .Y(_0058_),
    .B1(_0369_));
 sg13g2_o21ai_1 _1925_ (.B1(net507),
    .Y(_0370_),
    .A1(net958),
    .A2(net394));
 sg13g2_a21oi_1 _1926_ (.A1(net524),
    .A2(net394),
    .Y(_0059_),
    .B1(_0370_));
 sg13g2_o21ai_1 _1927_ (.B1(net502),
    .Y(_0371_),
    .A1(net982),
    .A2(net394));
 sg13g2_a21oi_1 _1928_ (.A1(net525),
    .A2(net394),
    .Y(_0060_),
    .B1(_0371_));
 sg13g2_nor2b_2 _1929_ (.A(_0324_),
    .B_N(_0333_),
    .Y(_0372_));
 sg13g2_o21ai_1 _1930_ (.B1(net503),
    .Y(_0373_),
    .A1(net886),
    .A2(net391));
 sg13g2_a21oi_1 _1931_ (.A1(net517),
    .A2(net391),
    .Y(_0061_),
    .B1(_0373_));
 sg13g2_o21ai_1 _1932_ (.B1(net501),
    .Y(_0374_),
    .A1(net846),
    .A2(net391));
 sg13g2_a21oi_1 _1933_ (.A1(net519),
    .A2(net391),
    .Y(_0062_),
    .B1(_0374_));
 sg13g2_o21ai_1 _1934_ (.B1(net493),
    .Y(_0375_),
    .A1(net936),
    .A2(net391));
 sg13g2_a21oi_1 _1935_ (.A1(net520),
    .A2(net391),
    .Y(_0063_),
    .B1(_0375_));
 sg13g2_o21ai_1 _1936_ (.B1(net501),
    .Y(_0376_),
    .A1(net834),
    .A2(net391));
 sg13g2_a21oi_1 _1937_ (.A1(net521),
    .A2(net391),
    .Y(_0064_),
    .B1(_0376_));
 sg13g2_o21ai_1 _1938_ (.B1(net506),
    .Y(_0377_),
    .A1(net918),
    .A2(net392));
 sg13g2_a21oi_1 _1939_ (.A1(net522),
    .A2(net392),
    .Y(_0065_),
    .B1(_0377_));
 sg13g2_o21ai_1 _1940_ (.B1(net506),
    .Y(_0378_),
    .A1(net843),
    .A2(net392));
 sg13g2_a21oi_1 _1941_ (.A1(net523),
    .A2(net392),
    .Y(_0066_),
    .B1(_0378_));
 sg13g2_o21ai_1 _1942_ (.B1(net507),
    .Y(_0379_),
    .A1(net841),
    .A2(net392));
 sg13g2_a21oi_1 _1943_ (.A1(net524),
    .A2(net392),
    .Y(_0067_),
    .B1(_0379_));
 sg13g2_o21ai_1 _1944_ (.B1(net503),
    .Y(_0380_),
    .A1(net837),
    .A2(net392));
 sg13g2_a21oi_1 _1945_ (.A1(net525),
    .A2(net392),
    .Y(_0068_),
    .B1(_0380_));
 sg13g2_nor2_2 _1946_ (.A(_0324_),
    .B(_0343_),
    .Y(_0381_));
 sg13g2_o21ai_1 _1947_ (.B1(net503),
    .Y(_0382_),
    .A1(net888),
    .A2(net389));
 sg13g2_a21oi_1 _1948_ (.A1(net517),
    .A2(net389),
    .Y(_0069_),
    .B1(_0382_));
 sg13g2_o21ai_1 _1949_ (.B1(net500),
    .Y(_0383_),
    .A1(net910),
    .A2(net389));
 sg13g2_a21oi_1 _1950_ (.A1(net519),
    .A2(net389),
    .Y(_0070_),
    .B1(_0383_));
 sg13g2_o21ai_1 _1951_ (.B1(net493),
    .Y(_0384_),
    .A1(net878),
    .A2(net389));
 sg13g2_a21oi_1 _1952_ (.A1(net520),
    .A2(net389),
    .Y(_0071_),
    .B1(_0384_));
 sg13g2_o21ai_1 _1953_ (.B1(net501),
    .Y(_0385_),
    .A1(net996),
    .A2(net389));
 sg13g2_a21oi_1 _1954_ (.A1(net521),
    .A2(net389),
    .Y(_0072_),
    .B1(_0385_));
 sg13g2_o21ai_1 _1955_ (.B1(net506),
    .Y(_0386_),
    .A1(net894),
    .A2(net390));
 sg13g2_a21oi_1 _1956_ (.A1(net522),
    .A2(net390),
    .Y(_0073_),
    .B1(_0386_));
 sg13g2_o21ai_1 _1957_ (.B1(net510),
    .Y(_0387_),
    .A1(net828),
    .A2(net390));
 sg13g2_a21oi_1 _1958_ (.A1(net523),
    .A2(net390),
    .Y(_0074_),
    .B1(_0387_));
 sg13g2_o21ai_1 _1959_ (.B1(net507),
    .Y(_0388_),
    .A1(net839),
    .A2(net390));
 sg13g2_a21oi_1 _1960_ (.A1(net524),
    .A2(net390),
    .Y(_0075_),
    .B1(_0388_));
 sg13g2_o21ai_1 _1961_ (.B1(net504),
    .Y(_0389_),
    .A1(net903),
    .A2(net390));
 sg13g2_a21oi_1 _1962_ (.A1(net525),
    .A2(net390),
    .Y(_0076_),
    .B1(_0389_));
 sg13g2_nor2_2 _1963_ (.A(_0324_),
    .B(_0353_),
    .Y(_0390_));
 sg13g2_o21ai_1 _1964_ (.B1(net503),
    .Y(_0391_),
    .A1(net867),
    .A2(net387));
 sg13g2_a21oi_1 _1965_ (.A1(net517),
    .A2(net388),
    .Y(_0077_),
    .B1(_0391_));
 sg13g2_o21ai_1 _1966_ (.B1(net501),
    .Y(_0392_),
    .A1(net928),
    .A2(net388));
 sg13g2_a21oi_1 _1967_ (.A1(net519),
    .A2(net388),
    .Y(_0078_),
    .B1(_0392_));
 sg13g2_o21ai_1 _1968_ (.B1(net494),
    .Y(_0393_),
    .A1(net990),
    .A2(net388));
 sg13g2_a21oi_1 _1969_ (.A1(net520),
    .A2(net388),
    .Y(_0079_),
    .B1(_0393_));
 sg13g2_o21ai_1 _1970_ (.B1(net504),
    .Y(_0394_),
    .A1(net871),
    .A2(net388));
 sg13g2_a21oi_1 _1971_ (.A1(net521),
    .A2(net388),
    .Y(_0080_),
    .B1(_0394_));
 sg13g2_o21ai_1 _1972_ (.B1(net506),
    .Y(_0395_),
    .A1(net984),
    .A2(net387));
 sg13g2_a21oi_1 _1973_ (.A1(net522),
    .A2(net387),
    .Y(_0081_),
    .B1(_0395_));
 sg13g2_o21ai_1 _1974_ (.B1(net506),
    .Y(_0396_),
    .A1(net942),
    .A2(net387));
 sg13g2_a21oi_1 _1975_ (.A1(net523),
    .A2(net387),
    .Y(_0082_),
    .B1(_0396_));
 sg13g2_o21ai_1 _1976_ (.B1(net507),
    .Y(_0397_),
    .A1(net947),
    .A2(net387));
 sg13g2_a21oi_1 _1977_ (.A1(net524),
    .A2(_0390_),
    .Y(_0083_),
    .B1(_0397_));
 sg13g2_o21ai_1 _1978_ (.B1(net503),
    .Y(_0398_),
    .A1(net924),
    .A2(net387));
 sg13g2_a21oi_1 _1979_ (.A1(net525),
    .A2(net387),
    .Y(_0084_),
    .B1(_0398_));
 sg13g2_o21ai_1 _1980_ (.B1(net503),
    .Y(_0399_),
    .A1(net954),
    .A2(net401));
 sg13g2_a21oi_1 _1981_ (.A1(net518),
    .A2(net401),
    .Y(_0085_),
    .B1(_0399_));
 sg13g2_o21ai_1 _1982_ (.B1(net500),
    .Y(_0400_),
    .A1(net854),
    .A2(net402));
 sg13g2_a21oi_1 _1983_ (.A1(net519),
    .A2(net402),
    .Y(_0086_),
    .B1(_0400_));
 sg13g2_o21ai_1 _1984_ (.B1(net493),
    .Y(_0401_),
    .A1(net1000),
    .A2(net402));
 sg13g2_a21oi_1 _1985_ (.A1(net520),
    .A2(net402),
    .Y(_0087_),
    .B1(_0401_));
 sg13g2_o21ai_1 _1986_ (.B1(net504),
    .Y(_0402_),
    .A1(net876),
    .A2(net402));
 sg13g2_a21oi_1 _1987_ (.A1(_0894_),
    .A2(net402),
    .Y(_0088_),
    .B1(_0402_));
 sg13g2_o21ai_1 _1988_ (.B1(net506),
    .Y(_0403_),
    .A1(net830),
    .A2(net401));
 sg13g2_a21oi_1 _1989_ (.A1(net522),
    .A2(net401),
    .Y(_0089_),
    .B1(_0403_));
 sg13g2_o21ai_1 _1990_ (.B1(net506),
    .Y(_0404_),
    .A1(net932),
    .A2(net401));
 sg13g2_a21oi_1 _1991_ (.A1(net523),
    .A2(net403),
    .Y(_0090_),
    .B1(_0404_));
 sg13g2_o21ai_1 _1992_ (.B1(net507),
    .Y(_0405_),
    .A1(net820),
    .A2(net403));
 sg13g2_a21oi_1 _1993_ (.A1(net524),
    .A2(net403),
    .Y(_0091_),
    .B1(_0405_));
 sg13g2_o21ai_1 _1994_ (.B1(net502),
    .Y(_0406_),
    .A1(net930),
    .A2(net401));
 sg13g2_a21oi_1 _1995_ (.A1(net525),
    .A2(net401),
    .Y(_0092_),
    .B1(_0406_));
 sg13g2_nor2_1 _1996_ (.A(_0313_),
    .B(_0318_),
    .Y(_0407_));
 sg13g2_nand2_2 _1997_ (.Y(_0408_),
    .A(_0319_),
    .B(net431));
 sg13g2_nor2_2 _1998_ (.A(net518),
    .B(net457),
    .Y(_0409_));
 sg13g2_a22oi_1 _1999_ (.Y(_0410_),
    .B1(_0409_),
    .B2(net431),
    .A2(_0408_),
    .A1(net793));
 sg13g2_nor2_1 _2000_ (.A(net470),
    .B(_0410_),
    .Y(_0093_));
 sg13g2_nor2_2 _2001_ (.A(_0898_),
    .B(net458),
    .Y(_0411_));
 sg13g2_a22oi_1 _2002_ (.Y(_0412_),
    .B1(_0411_),
    .B2(net431),
    .A2(_0408_),
    .A1(net725));
 sg13g2_nor2_1 _2003_ (.A(net469),
    .B(_0412_),
    .Y(_0094_));
 sg13g2_nor2_2 _2004_ (.A(_0896_),
    .B(net457),
    .Y(_0413_));
 sg13g2_a22oi_1 _2005_ (.Y(_0414_),
    .B1(_0413_),
    .B2(net431),
    .A2(_0408_),
    .A1(net774));
 sg13g2_nor2_1 _2006_ (.A(net469),
    .B(_0414_),
    .Y(_0095_));
 sg13g2_o21ai_1 _2007_ (.B1(net495),
    .Y(_0415_),
    .A1(net548),
    .A2(_0408_));
 sg13g2_a21oi_1 _2008_ (.A1(_0881_),
    .A2(_0408_),
    .Y(_0096_),
    .B1(_0415_));
 sg13g2_nor2_2 _2009_ (.A(\u_model_loader.byte_idx_q[3] ),
    .B(_0885_),
    .Y(_0416_));
 sg13g2_nor2b_2 _2010_ (.A(net546),
    .B_N(_0416_),
    .Y(_0417_));
 sg13g2_nand2_2 _2011_ (.Y(_0418_),
    .A(net431),
    .B(_0417_));
 sg13g2_and2_1 _2012_ (.A(net552),
    .B(_0417_),
    .X(_0419_));
 sg13g2_a22oi_1 _2013_ (.Y(_0420_),
    .B1(_0419_),
    .B2(net431),
    .A2(_0418_),
    .A1(net851));
 sg13g2_nor2_1 _2014_ (.A(net469),
    .B(_0420_),
    .Y(_0097_));
 sg13g2_and2_1 _2015_ (.A(net551),
    .B(_0417_),
    .X(_0421_));
 sg13g2_a22oi_1 _2016_ (.Y(_0422_),
    .B1(_0421_),
    .B2(net431),
    .A2(_0418_),
    .A1(net775));
 sg13g2_nor2_1 _2017_ (.A(net469),
    .B(_0422_),
    .Y(_0098_));
 sg13g2_and2_1 _2018_ (.A(net550),
    .B(_0417_),
    .X(_0423_));
 sg13g2_a22oi_1 _2019_ (.Y(_0424_),
    .B1(_0423_),
    .B2(net431),
    .A2(_0418_),
    .A1(net810));
 sg13g2_nor2_1 _2020_ (.A(net470),
    .B(_0424_),
    .Y(_0099_));
 sg13g2_o21ai_1 _2021_ (.B1(net495),
    .Y(_0425_),
    .A1(net548),
    .A2(_0418_));
 sg13g2_a21oi_1 _2022_ (.A1(_0879_),
    .A2(_0418_),
    .Y(_0100_),
    .B1(_0425_));
 sg13g2_nor2b_2 _2023_ (.A(\u_model_loader.byte_idx_q[2] ),
    .B_N(\u_model_loader.byte_idx_q[3] ),
    .Y(_0426_));
 sg13g2_nor2b_2 _2024_ (.A(net546),
    .B_N(_0426_),
    .Y(_0427_));
 sg13g2_and2_1 _2025_ (.A(net433),
    .B(net456),
    .X(_0428_));
 sg13g2_nand2_2 _2026_ (.Y(_0429_),
    .A(net433),
    .B(net456));
 sg13g2_a21oi_1 _2027_ (.A1(net552),
    .A2(net457),
    .Y(_0430_),
    .B1(_0429_));
 sg13g2_o21ai_1 _2028_ (.B1(net495),
    .Y(_0431_),
    .A1(net896),
    .A2(_0428_));
 sg13g2_nor2_1 _2029_ (.A(_0430_),
    .B(net897),
    .Y(_0101_));
 sg13g2_a21oi_1 _2030_ (.A1(net551),
    .A2(net457),
    .Y(_0432_),
    .B1(_0429_));
 sg13g2_o21ai_1 _2031_ (.B1(net495),
    .Y(_0433_),
    .A1(net907),
    .A2(_0428_));
 sg13g2_nor2_1 _2032_ (.A(_0432_),
    .B(net908),
    .Y(_0102_));
 sg13g2_a21oi_1 _2033_ (.A1(net550),
    .A2(net457),
    .Y(_0434_),
    .B1(_0429_));
 sg13g2_o21ai_1 _2034_ (.B1(net495),
    .Y(_0435_),
    .A1(net1004),
    .A2(_0428_));
 sg13g2_nor2_1 _2035_ (.A(_0434_),
    .B(net1005),
    .Y(_0103_));
 sg13g2_and2_1 _2036_ (.A(net548),
    .B(_0427_),
    .X(_0436_));
 sg13g2_a22oi_1 _2037_ (.Y(_0437_),
    .B1(_0436_),
    .B2(net433),
    .A2(_0429_),
    .A1(net737));
 sg13g2_nor2_1 _2038_ (.A(net473),
    .B(_0437_),
    .Y(_0104_));
 sg13g2_nor2_2 _2039_ (.A(net545),
    .B(_0316_),
    .Y(_0438_));
 sg13g2_nand2_2 _2040_ (.Y(_0439_),
    .A(net433),
    .B(_0438_));
 sg13g2_nor3_2 _2041_ (.A(net545),
    .B(net518),
    .C(_0316_),
    .Y(_0440_));
 sg13g2_a22oi_1 _2042_ (.Y(_0441_),
    .B1(_0440_),
    .B2(net433),
    .A2(_0439_),
    .A1(net740));
 sg13g2_nor2_1 _2043_ (.A(net470),
    .B(net741),
    .Y(_0105_));
 sg13g2_nor3_2 _2044_ (.A(net545),
    .B(_0898_),
    .C(_0316_),
    .Y(_0442_));
 sg13g2_a22oi_1 _2045_ (.Y(_0443_),
    .B1(_0442_),
    .B2(net433),
    .A2(_0439_),
    .A1(net757));
 sg13g2_nor2_1 _2046_ (.A(net473),
    .B(net758),
    .Y(_0106_));
 sg13g2_nor3_2 _2047_ (.A(net545),
    .B(_0896_),
    .C(_0316_),
    .Y(_0444_));
 sg13g2_a22oi_1 _2048_ (.Y(_0445_),
    .B1(_0444_),
    .B2(net433),
    .A2(_0439_),
    .A1(net721));
 sg13g2_nor2_1 _2049_ (.A(net473),
    .B(net722),
    .Y(_0107_));
 sg13g2_and2_1 _2050_ (.A(net549),
    .B(_0317_),
    .X(_0446_));
 sg13g2_nor2_1 _2051_ (.A(_0894_),
    .B(_0318_),
    .Y(_0447_));
 sg13g2_a22oi_1 _2052_ (.Y(_0448_),
    .B1(_0447_),
    .B2(_0328_),
    .A2(_0439_),
    .A1(net727));
 sg13g2_nor2_1 _2053_ (.A(net473),
    .B(net728),
    .Y(_0108_));
 sg13g2_and2_1 _2054_ (.A(net546),
    .B(_0315_),
    .X(_0449_));
 sg13g2_nand2_2 _2055_ (.Y(_0450_),
    .A(net432),
    .B(_0449_));
 sg13g2_and2_1 _2056_ (.A(net552),
    .B(_0449_),
    .X(_0451_));
 sg13g2_a22oi_1 _2057_ (.Y(_0452_),
    .B1(_0451_),
    .B2(net432),
    .A2(_0450_),
    .A1(net767));
 sg13g2_nor2_1 _2058_ (.A(net478),
    .B(_0452_),
    .Y(_0109_));
 sg13g2_and2_1 _2059_ (.A(net551),
    .B(_0449_),
    .X(_0453_));
 sg13g2_a22oi_1 _2060_ (.Y(_0454_),
    .B1(_0453_),
    .B2(net432),
    .A2(_0450_),
    .A1(net782));
 sg13g2_nor2_1 _2061_ (.A(net478),
    .B(_0454_),
    .Y(_0110_));
 sg13g2_and2_1 _2062_ (.A(net550),
    .B(_0449_),
    .X(_0455_));
 sg13g2_a22oi_1 _2063_ (.Y(_0456_),
    .B1(_0455_),
    .B2(net432),
    .A2(_0450_),
    .A1(net813));
 sg13g2_nor2_1 _2064_ (.A(net471),
    .B(_0456_),
    .Y(_0111_));
 sg13g2_o21ai_1 _2065_ (.B1(net499),
    .Y(_0457_),
    .A1(net548),
    .A2(_0450_));
 sg13g2_a21oi_1 _2066_ (.A1(_0873_),
    .A2(_0450_),
    .Y(_0112_),
    .B1(_0457_));
 sg13g2_and2_1 _2067_ (.A(net546),
    .B(_0416_),
    .X(_0458_));
 sg13g2_nand2_2 _2068_ (.Y(_0459_),
    .A(net432),
    .B(_0458_));
 sg13g2_and2_1 _2069_ (.A(net552),
    .B(_0458_),
    .X(_0460_));
 sg13g2_a22oi_1 _2070_ (.Y(_0461_),
    .B1(_0460_),
    .B2(net432),
    .A2(_0459_),
    .A1(net765));
 sg13g2_nor2_1 _2071_ (.A(net478),
    .B(_0461_),
    .Y(_0113_));
 sg13g2_and2_1 _2072_ (.A(net551),
    .B(_0458_),
    .X(_0462_));
 sg13g2_a22oi_1 _2073_ (.Y(_0463_),
    .B1(_0462_),
    .B2(net432),
    .A2(_0459_),
    .A1(net826));
 sg13g2_nor2_1 _2074_ (.A(net478),
    .B(_0463_),
    .Y(_0114_));
 sg13g2_and2_1 _2075_ (.A(net550),
    .B(_0458_),
    .X(_0464_));
 sg13g2_a22oi_1 _2076_ (.Y(_0465_),
    .B1(_0464_),
    .B2(net432),
    .A2(_0459_),
    .A1(net786));
 sg13g2_nor2_1 _2077_ (.A(net472),
    .B(_0465_),
    .Y(_0115_));
 sg13g2_o21ai_1 _2078_ (.B1(net499),
    .Y(_0466_),
    .A1(net548),
    .A2(_0459_));
 sg13g2_a21oi_1 _2079_ (.A1(_0872_),
    .A2(_0459_),
    .Y(_0116_),
    .B1(_0466_));
 sg13g2_and2_1 _2080_ (.A(net546),
    .B(_0426_),
    .X(_0467_));
 sg13g2_nand2_2 _2081_ (.Y(_0468_),
    .A(net433),
    .B(_0467_));
 sg13g2_and2_1 _2082_ (.A(net552),
    .B(_0467_),
    .X(_0469_));
 sg13g2_a22oi_1 _2083_ (.Y(_0470_),
    .B1(_0469_),
    .B2(net434),
    .A2(_0468_),
    .A1(net790));
 sg13g2_nor2_1 _2084_ (.A(net479),
    .B(_0470_),
    .Y(_0117_));
 sg13g2_and2_1 _2085_ (.A(\model_byte[1] ),
    .B(_0467_),
    .X(_0471_));
 sg13g2_a22oi_1 _2086_ (.Y(_0472_),
    .B1(_0471_),
    .B2(net434),
    .A2(_0468_),
    .A1(net713));
 sg13g2_nor2_1 _2087_ (.A(net479),
    .B(net714),
    .Y(_0118_));
 sg13g2_and2_1 _2088_ (.A(net550),
    .B(_0467_),
    .X(_0473_));
 sg13g2_a22oi_1 _2089_ (.Y(_0474_),
    .B1(_0473_),
    .B2(net434),
    .A2(_0468_),
    .A1(net707));
 sg13g2_nor2_1 _2090_ (.A(net475),
    .B(_0474_),
    .Y(_0119_));
 sg13g2_o21ai_1 _2091_ (.B1(net498),
    .Y(_0475_),
    .A1(net548),
    .A2(_0468_));
 sg13g2_a21oi_1 _2092_ (.A1(_0869_),
    .A2(_0468_),
    .Y(_0120_),
    .B1(_0475_));
 sg13g2_nor2_2 _2093_ (.A(_0314_),
    .B(_0353_),
    .Y(_0476_));
 sg13g2_nand2_2 _2094_ (.Y(_0477_),
    .A(_0319_),
    .B(net453));
 sg13g2_and2_1 _2095_ (.A(_0317_),
    .B(net454),
    .X(_0478_));
 sg13g2_a22oi_1 _2096_ (.Y(_0479_),
    .B1(net428),
    .B2(_0409_),
    .A2(_0477_),
    .A1(net848));
 sg13g2_nor2_1 _2097_ (.A(net470),
    .B(_0479_),
    .Y(_0121_));
 sg13g2_a22oi_1 _2098_ (.Y(_0480_),
    .B1(net428),
    .B2(_0411_),
    .A2(_0477_),
    .A1(net807));
 sg13g2_nor2_1 _2099_ (.A(net469),
    .B(_0480_),
    .Y(_0122_));
 sg13g2_a22oi_1 _2100_ (.Y(_0481_),
    .B1(net428),
    .B2(_0413_),
    .A2(_0477_),
    .A1(net770));
 sg13g2_nor2_1 _2101_ (.A(net469),
    .B(_0481_),
    .Y(_0123_));
 sg13g2_o21ai_1 _2102_ (.B1(net495),
    .Y(_0482_),
    .A1(net455),
    .A2(_0477_));
 sg13g2_a21oi_1 _2103_ (.A1(_0867_),
    .A2(_0477_),
    .Y(_0124_),
    .B1(_0482_));
 sg13g2_nand2_2 _2104_ (.Y(_0483_),
    .A(_0417_),
    .B(net453));
 sg13g2_a22oi_1 _2105_ (.Y(_0484_),
    .B1(_0483_),
    .B2(net628),
    .A2(net428),
    .A1(_0419_));
 sg13g2_nor2_1 _2106_ (.A(net469),
    .B(_0484_),
    .Y(_0125_));
 sg13g2_a22oi_1 _2107_ (.Y(_0485_),
    .B1(_0483_),
    .B2(net590),
    .A2(net428),
    .A1(_0421_));
 sg13g2_nor2_1 _2108_ (.A(net469),
    .B(_0485_),
    .Y(_0126_));
 sg13g2_a22oi_1 _2109_ (.Y(_0486_),
    .B1(_0483_),
    .B2(net648),
    .A2(net428),
    .A1(_0423_));
 sg13g2_nor2_1 _2110_ (.A(net470),
    .B(_0486_),
    .Y(_0127_));
 sg13g2_o21ai_1 _2111_ (.B1(net495),
    .Y(_0487_),
    .A1(net455),
    .A2(_0483_));
 sg13g2_a21oi_1 _2112_ (.A1(_0865_),
    .A2(_0483_),
    .Y(_0128_),
    .B1(_0487_));
 sg13g2_and2_1 _2113_ (.A(net456),
    .B(net453),
    .X(_0488_));
 sg13g2_nand2_1 _2114_ (.Y(_0489_),
    .A(net456),
    .B(net453));
 sg13g2_a21oi_1 _2115_ (.A1(net552),
    .A2(net457),
    .Y(_0490_),
    .B1(_0489_));
 sg13g2_o21ai_1 _2116_ (.B1(net496),
    .Y(_0491_),
    .A1(net1030),
    .A2(_0488_));
 sg13g2_nor2_1 _2117_ (.A(_0490_),
    .B(_0491_),
    .Y(_0129_));
 sg13g2_a21oi_1 _2118_ (.A1(net551),
    .A2(net457),
    .Y(_0492_),
    .B1(_0489_));
 sg13g2_o21ai_1 _2119_ (.B1(net494),
    .Y(_0493_),
    .A1(net970),
    .A2(_0488_));
 sg13g2_nor2_1 _2120_ (.A(_0492_),
    .B(_0493_),
    .Y(_0130_));
 sg13g2_a21oi_1 _2121_ (.A1(net550),
    .A2(net457),
    .Y(_0494_),
    .B1(_0489_));
 sg13g2_o21ai_1 _2122_ (.B1(net494),
    .Y(_0495_),
    .A1(net905),
    .A2(_0488_));
 sg13g2_nor2_1 _2123_ (.A(_0494_),
    .B(_0495_),
    .Y(_0131_));
 sg13g2_a22oi_1 _2124_ (.Y(_0496_),
    .B1(_0489_),
    .B2(net642),
    .A2(net454),
    .A1(_0436_));
 sg13g2_nor2_1 _2125_ (.A(net474),
    .B(_0496_),
    .Y(_0132_));
 sg13g2_nand2_2 _2126_ (.Y(_0497_),
    .A(_0438_),
    .B(net454));
 sg13g2_a22oi_1 _2127_ (.Y(_0498_),
    .B1(_0497_),
    .B2(net686),
    .A2(net453),
    .A1(_0440_));
 sg13g2_nor2_1 _2128_ (.A(net470),
    .B(net687),
    .Y(_0133_));
 sg13g2_a22oi_1 _2129_ (.Y(_0499_),
    .B1(_0497_),
    .B2(net668),
    .A2(net454),
    .A1(_0442_));
 sg13g2_nor2_1 _2130_ (.A(net473),
    .B(net669),
    .Y(_0134_));
 sg13g2_a22oi_1 _2131_ (.Y(_0500_),
    .B1(_0497_),
    .B2(net597),
    .A2(net454),
    .A1(_0444_));
 sg13g2_nor2_1 _2132_ (.A(net473),
    .B(net598),
    .Y(_0135_));
 sg13g2_o21ai_1 _2133_ (.B1(net495),
    .Y(_0501_),
    .A1(net548),
    .A2(_0497_));
 sg13g2_a21oi_1 _2134_ (.A1(_0860_),
    .A2(_0497_),
    .Y(_0136_),
    .B1(_0501_));
 sg13g2_nand2_2 _2135_ (.Y(_0502_),
    .A(_0449_),
    .B(net453));
 sg13g2_a22oi_1 _2136_ (.Y(_0503_),
    .B1(_0502_),
    .B2(net678),
    .A2(net428),
    .A1(_0451_));
 sg13g2_nor2_1 _2137_ (.A(net478),
    .B(_0503_),
    .Y(_0137_));
 sg13g2_a22oi_1 _2138_ (.Y(_0504_),
    .B1(_0502_),
    .B2(net637),
    .A2(net428),
    .A1(_0453_));
 sg13g2_nor2_1 _2139_ (.A(net478),
    .B(_0504_),
    .Y(_0138_));
 sg13g2_a22oi_1 _2140_ (.Y(_0505_),
    .B1(_0502_),
    .B2(net680),
    .A2(net429),
    .A1(_0455_));
 sg13g2_nor2_1 _2141_ (.A(net471),
    .B(_0505_),
    .Y(_0139_));
 sg13g2_o21ai_1 _2142_ (.B1(net499),
    .Y(_0506_),
    .A1(net455),
    .A2(_0502_));
 sg13g2_a21oi_1 _2143_ (.A1(_0859_),
    .A2(_0502_),
    .Y(_0140_),
    .B1(_0506_));
 sg13g2_nand2_2 _2144_ (.Y(_0507_),
    .A(_0458_),
    .B(net453));
 sg13g2_a22oi_1 _2145_ (.Y(_0508_),
    .B1(_0507_),
    .B2(net651),
    .A2(net429),
    .A1(_0460_));
 sg13g2_nor2_1 _2146_ (.A(net471),
    .B(_0508_),
    .Y(_0141_));
 sg13g2_a22oi_1 _2147_ (.Y(_0509_),
    .B1(_0507_),
    .B2(net627),
    .A2(net429),
    .A1(_0462_));
 sg13g2_nor2_1 _2148_ (.A(net471),
    .B(_0509_),
    .Y(_0142_));
 sg13g2_a22oi_1 _2149_ (.Y(_0510_),
    .B1(_0507_),
    .B2(net670),
    .A2(net429),
    .A1(_0464_));
 sg13g2_nor2_1 _2150_ (.A(net471),
    .B(_0510_),
    .Y(_0143_));
 sg13g2_o21ai_1 _2151_ (.B1(net499),
    .Y(_0511_),
    .A1(net455),
    .A2(_0507_));
 sg13g2_a21oi_1 _2152_ (.A1(_0858_),
    .A2(_0507_),
    .Y(_0144_),
    .B1(_0511_));
 sg13g2_nand2_2 _2153_ (.Y(_0512_),
    .A(_0467_),
    .B(net453));
 sg13g2_a22oi_1 _2154_ (.Y(_0513_),
    .B1(_0512_),
    .B2(net629),
    .A2(net430),
    .A1(_0469_));
 sg13g2_nor2_1 _2155_ (.A(net476),
    .B(_0513_),
    .Y(_0145_));
 sg13g2_a22oi_1 _2156_ (.Y(_0514_),
    .B1(_0512_),
    .B2(net614),
    .A2(net430),
    .A1(_0471_));
 sg13g2_nor2_1 _2157_ (.A(net476),
    .B(net615),
    .Y(_0146_));
 sg13g2_a22oi_1 _2158_ (.Y(_0515_),
    .B1(_0512_),
    .B2(net596),
    .A2(net430),
    .A1(_0473_));
 sg13g2_nor2_1 _2159_ (.A(net475),
    .B(_0515_),
    .Y(_0147_));
 sg13g2_o21ai_1 _2160_ (.B1(net498),
    .Y(_0516_),
    .A1(_0446_),
    .A2(_0512_));
 sg13g2_a21oi_1 _2161_ (.A1(_0857_),
    .A2(_0512_),
    .Y(_0148_),
    .B1(_0516_));
 sg13g2_nor2_1 _2162_ (.A(_0314_),
    .B(_0343_),
    .Y(_0517_));
 sg13g2_nand2_2 _2163_ (.Y(_0518_),
    .A(_0319_),
    .B(net451));
 sg13g2_and2_1 _2164_ (.A(_0317_),
    .B(net451),
    .X(_0519_));
 sg13g2_a22oi_1 _2165_ (.Y(_0520_),
    .B1(net424),
    .B2(_0409_),
    .A2(net426),
    .A1(net776));
 sg13g2_nor2_1 _2166_ (.A(net475),
    .B(_0520_),
    .Y(_0149_));
 sg13g2_a22oi_1 _2167_ (.Y(_0521_),
    .B1(net425),
    .B2(_0411_),
    .A2(net426),
    .A1(net708));
 sg13g2_nor2_1 _2168_ (.A(net475),
    .B(_0521_),
    .Y(_0150_));
 sg13g2_a22oi_1 _2169_ (.Y(_0522_),
    .B1(net424),
    .B2(_0413_),
    .A2(net426),
    .A1(net769));
 sg13g2_nor2_1 _2170_ (.A(net475),
    .B(_0522_),
    .Y(_0151_));
 sg13g2_o21ai_1 _2171_ (.B1(net512),
    .Y(_0523_),
    .A1(net455),
    .A2(net426));
 sg13g2_a21oi_1 _2172_ (.A1(_0856_),
    .A2(net426),
    .Y(_0152_),
    .B1(_0523_));
 sg13g2_o21ai_1 _2173_ (.B1(net514),
    .Y(_0524_),
    .A1(\model_byte[4] ),
    .A2(net426));
 sg13g2_a21oi_1 _2174_ (.A1(_0855_),
    .A2(net426),
    .Y(_0153_),
    .B1(_0524_));
 sg13g2_o21ai_1 _2175_ (.B1(net514),
    .Y(_0525_),
    .A1(\model_byte[5] ),
    .A2(net426));
 sg13g2_a21oi_1 _2176_ (.A1(_0854_),
    .A2(net427),
    .Y(_0154_),
    .B1(_0525_));
 sg13g2_o21ai_1 _2177_ (.B1(net514),
    .Y(_0526_),
    .A1(\model_byte[6] ),
    .A2(net427));
 sg13g2_a21oi_1 _2178_ (.A1(_0853_),
    .A2(net427),
    .Y(_0155_),
    .B1(_0526_));
 sg13g2_o21ai_1 _2179_ (.B1(net514),
    .Y(_0527_),
    .A1(\model_byte[7] ),
    .A2(net427));
 sg13g2_a21oi_1 _2180_ (.A1(_0852_),
    .A2(net427),
    .Y(_0156_),
    .B1(_0527_));
 sg13g2_nand2_1 _2181_ (.Y(_0528_),
    .A(_0417_),
    .B(net451));
 sg13g2_a22oi_1 _2182_ (.Y(_0529_),
    .B1(net405),
    .B2(net585),
    .A2(net423),
    .A1(_0419_));
 sg13g2_nor2_1 _2183_ (.A(net472),
    .B(_0529_),
    .Y(_0157_));
 sg13g2_a22oi_1 _2184_ (.Y(_0530_),
    .B1(net405),
    .B2(net647),
    .A2(net423),
    .A1(_0421_));
 sg13g2_nor2_1 _2185_ (.A(net472),
    .B(_0530_),
    .Y(_0158_));
 sg13g2_a22oi_1 _2186_ (.Y(_0531_),
    .B1(net405),
    .B2(net659),
    .A2(net423),
    .A1(_0423_));
 sg13g2_nor2_1 _2187_ (.A(net476),
    .B(_0531_),
    .Y(_0159_));
 sg13g2_o21ai_1 _2188_ (.B1(net512),
    .Y(_0532_),
    .A1(net549),
    .A2(net405));
 sg13g2_a21oi_1 _2189_ (.A1(_0848_),
    .A2(_0528_),
    .Y(_0160_),
    .B1(_0532_));
 sg13g2_and2_1 _2190_ (.A(\model_byte[4] ),
    .B(_0416_),
    .X(_0533_));
 sg13g2_nor2b_2 _2191_ (.A(_0321_),
    .B_N(net451),
    .Y(_0534_));
 sg13g2_a22oi_1 _2192_ (.Y(_0535_),
    .B1(_0533_),
    .B2(_0534_),
    .A2(net405),
    .A1(net805));
 sg13g2_nor2_1 _2193_ (.A(net483),
    .B(net806),
    .Y(_0161_));
 sg13g2_and2_1 _2194_ (.A(\model_byte[5] ),
    .B(_0416_),
    .X(_0536_));
 sg13g2_a22oi_1 _2195_ (.Y(_0537_),
    .B1(_0534_),
    .B2(_0536_),
    .A2(net405),
    .A1(net835));
 sg13g2_nor2_1 _2196_ (.A(net484),
    .B(net836),
    .Y(_0162_));
 sg13g2_and2_1 _2197_ (.A(\model_byte[6] ),
    .B(_0416_),
    .X(_0538_));
 sg13g2_a22oi_1 _2198_ (.Y(_0539_),
    .B1(_0534_),
    .B2(_0538_),
    .A2(net405),
    .A1(net746));
 sg13g2_nor2_1 _2199_ (.A(net483),
    .B(net747),
    .Y(_0163_));
 sg13g2_and2_1 _2200_ (.A(\model_byte[7] ),
    .B(_0416_),
    .X(_0540_));
 sg13g2_a22oi_1 _2201_ (.Y(_0541_),
    .B1(_0534_),
    .B2(_0540_),
    .A2(net405),
    .A1(net711));
 sg13g2_nor2_1 _2202_ (.A(net483),
    .B(net712),
    .Y(_0164_));
 sg13g2_nand2_2 _2203_ (.Y(_0542_),
    .A(_0427_),
    .B(net452));
 sg13g2_a21oi_1 _2204_ (.A1(_0427_),
    .A2(net452),
    .Y(_0543_),
    .B1(net356));
 sg13g2_a21oi_1 _2205_ (.A1(net552),
    .A2(net458),
    .Y(_0544_),
    .B1(_0542_));
 sg13g2_nor3_1 _2206_ (.A(net486),
    .B(net357),
    .C(_0544_),
    .Y(_0165_));
 sg13g2_a21oi_1 _2207_ (.A1(net456),
    .A2(net452),
    .Y(_0545_),
    .B1(net372));
 sg13g2_a21oi_1 _2208_ (.A1(net551),
    .A2(net458),
    .Y(_0546_),
    .B1(_0542_));
 sg13g2_nor3_1 _2209_ (.A(net486),
    .B(_0545_),
    .C(_0546_),
    .Y(_0166_));
 sg13g2_a21oi_1 _2210_ (.A1(net456),
    .A2(net452),
    .Y(_0547_),
    .B1(net581));
 sg13g2_a21oi_1 _2211_ (.A1(net550),
    .A2(net458),
    .Y(_0548_),
    .B1(_0542_));
 sg13g2_nor3_1 _2212_ (.A(net486),
    .B(_0547_),
    .C(_0548_),
    .Y(_0167_));
 sg13g2_a22oi_1 _2213_ (.Y(_0549_),
    .B1(_0542_),
    .B2(net601),
    .A2(net452),
    .A1(_0436_));
 sg13g2_nor2_1 _2214_ (.A(net486),
    .B(_0549_),
    .Y(_0168_));
 sg13g2_and2_1 _2215_ (.A(\model_byte[4] ),
    .B(_0426_),
    .X(_0550_));
 sg13g2_a22oi_1 _2216_ (.Y(_0551_),
    .B1(_0550_),
    .B2(_0534_),
    .A2(_0542_),
    .A1(net780));
 sg13g2_nor2_1 _2217_ (.A(net483),
    .B(net781),
    .Y(_0169_));
 sg13g2_and2_1 _2218_ (.A(\model_byte[5] ),
    .B(_0426_),
    .X(_0552_));
 sg13g2_a22oi_1 _2219_ (.Y(_0553_),
    .B1(_0552_),
    .B2(_0534_),
    .A2(_0542_),
    .A1(net752));
 sg13g2_nor2_1 _2220_ (.A(net483),
    .B(net753),
    .Y(_0170_));
 sg13g2_and2_1 _2221_ (.A(\model_byte[6] ),
    .B(_0426_),
    .X(_0554_));
 sg13g2_a22oi_1 _2222_ (.Y(_0555_),
    .B1(_0554_),
    .B2(_0534_),
    .A2(_0542_),
    .A1(net803));
 sg13g2_nor2_1 _2223_ (.A(net483),
    .B(net804),
    .Y(_0171_));
 sg13g2_and2_1 _2224_ (.A(\model_byte[7] ),
    .B(_0426_),
    .X(_0556_));
 sg13g2_a22oi_1 _2225_ (.Y(_0557_),
    .B1(_0556_),
    .B2(_0534_),
    .A2(_0542_),
    .A1(net731));
 sg13g2_nor2_1 _2226_ (.A(net486),
    .B(net732),
    .Y(_0172_));
 sg13g2_and2_1 _2227_ (.A(_0438_),
    .B(net451),
    .X(_0558_));
 sg13g2_o21ai_1 _2228_ (.B1(net494),
    .Y(_0559_),
    .A1(net940),
    .A2(net421));
 sg13g2_a21oi_1 _2229_ (.A1(net517),
    .A2(net421),
    .Y(_0173_),
    .B1(_0559_));
 sg13g2_o21ai_1 _2230_ (.B1(net504),
    .Y(_0560_),
    .A1(net986),
    .A2(net421));
 sg13g2_a21oi_1 _2231_ (.A1(_0898_),
    .A2(net421),
    .Y(_0174_),
    .B1(_0560_));
 sg13g2_o21ai_1 _2232_ (.B1(net494),
    .Y(_0561_),
    .A1(net1007),
    .A2(net421));
 sg13g2_a21oi_1 _2233_ (.A1(_0896_),
    .A2(net421),
    .Y(_0175_),
    .B1(_0561_));
 sg13g2_o21ai_1 _2234_ (.B1(net504),
    .Y(_0562_),
    .A1(net946),
    .A2(net421));
 sg13g2_a21oi_1 _2235_ (.A1(net521),
    .A2(net422),
    .Y(_0176_),
    .B1(_0562_));
 sg13g2_o21ai_1 _2236_ (.B1(net509),
    .Y(_0563_),
    .A1(net1045),
    .A2(net422));
 sg13g2_a21oi_1 _2237_ (.A1(_0892_),
    .A2(net422),
    .Y(_0177_),
    .B1(_0563_));
 sg13g2_o21ai_1 _2238_ (.B1(net509),
    .Y(_0564_),
    .A1(net1043),
    .A2(net422));
 sg13g2_a21oi_1 _2239_ (.A1(_0890_),
    .A2(net422),
    .Y(_0178_),
    .B1(_0564_));
 sg13g2_o21ai_1 _2240_ (.B1(net509),
    .Y(_0565_),
    .A1(net1032),
    .A2(net422));
 sg13g2_a21oi_1 _2241_ (.A1(_0888_),
    .A2(net422),
    .Y(_0179_),
    .B1(_0565_));
 sg13g2_o21ai_1 _2242_ (.B1(net504),
    .Y(_0566_),
    .A1(net992),
    .A2(net421));
 sg13g2_a21oi_1 _2243_ (.A1(_0886_),
    .A2(_0558_),
    .Y(_0180_),
    .B1(_0566_));
 sg13g2_nand2_1 _2244_ (.Y(_0567_),
    .A(_0449_),
    .B(net451));
 sg13g2_a22oi_1 _2245_ (.Y(_0568_),
    .B1(net420),
    .B2(net662),
    .A2(net423),
    .A1(_0451_));
 sg13g2_nor2_1 _2246_ (.A(net477),
    .B(_0568_),
    .Y(_0181_));
 sg13g2_a22oi_1 _2247_ (.Y(_0569_),
    .B1(net420),
    .B2(net693),
    .A2(net423),
    .A1(_0453_));
 sg13g2_nor2_1 _2248_ (.A(net477),
    .B(_0569_),
    .Y(_0182_));
 sg13g2_a22oi_1 _2249_ (.Y(_0570_),
    .B1(net420),
    .B2(net661),
    .A2(net423),
    .A1(_0455_));
 sg13g2_nor2_1 _2250_ (.A(net472),
    .B(_0570_),
    .Y(_0183_));
 sg13g2_o21ai_1 _2251_ (.B1(net512),
    .Y(_0571_),
    .A1(net455),
    .A2(net419));
 sg13g2_a21oi_1 _2252_ (.A1(_0843_),
    .A2(net419),
    .Y(_0184_),
    .B1(_0571_));
 sg13g2_o21ai_1 _2253_ (.B1(net514),
    .Y(_0572_),
    .A1(\model_byte[4] ),
    .A2(net419));
 sg13g2_a21oi_1 _2254_ (.A1(_0842_),
    .A2(net419),
    .Y(_0185_),
    .B1(_0572_));
 sg13g2_o21ai_1 _2255_ (.B1(net514),
    .Y(_0573_),
    .A1(\model_byte[5] ),
    .A2(net419));
 sg13g2_a21oi_1 _2256_ (.A1(_0841_),
    .A2(net419),
    .Y(_0186_),
    .B1(_0573_));
 sg13g2_o21ai_1 _2257_ (.B1(net512),
    .Y(_0574_),
    .A1(\model_byte[6] ),
    .A2(net419));
 sg13g2_a21oi_1 _2258_ (.A1(_0840_),
    .A2(net419),
    .Y(_0187_),
    .B1(_0574_));
 sg13g2_o21ai_1 _2259_ (.B1(net512),
    .Y(_0575_),
    .A1(\model_byte[7] ),
    .A2(net420));
 sg13g2_a21oi_1 _2260_ (.A1(_0839_),
    .A2(net420),
    .Y(_0188_),
    .B1(_0575_));
 sg13g2_nand2_1 _2261_ (.Y(_0576_),
    .A(_0458_),
    .B(net451));
 sg13g2_a22oi_1 _2262_ (.Y(_0577_),
    .B1(net404),
    .B2(net605),
    .A2(net423),
    .A1(_0460_));
 sg13g2_nor2_1 _2263_ (.A(net477),
    .B(_0577_),
    .Y(_0189_));
 sg13g2_a22oi_1 _2264_ (.Y(_0578_),
    .B1(net404),
    .B2(net667),
    .A2(net423),
    .A1(_0462_));
 sg13g2_nor2_1 _2265_ (.A(net477),
    .B(_0578_),
    .Y(_0190_));
 sg13g2_a22oi_1 _2266_ (.Y(_0579_),
    .B1(net404),
    .B2(net613),
    .A2(net424),
    .A1(_0464_));
 sg13g2_nor2_1 _2267_ (.A(net472),
    .B(_0579_),
    .Y(_0191_));
 sg13g2_o21ai_1 _2268_ (.B1(net512),
    .Y(_0580_),
    .A1(net455),
    .A2(net404));
 sg13g2_a21oi_1 _2269_ (.A1(_0838_),
    .A2(_0576_),
    .Y(_0192_),
    .B1(_0580_));
 sg13g2_and2_1 _2270_ (.A(_0321_),
    .B(net425),
    .X(_0581_));
 sg13g2_a22oi_1 _2271_ (.Y(_0582_),
    .B1(_0581_),
    .B2(_0533_),
    .A2(net404),
    .A1(net759));
 sg13g2_nor2_1 _2272_ (.A(net483),
    .B(net760),
    .Y(_0193_));
 sg13g2_a22oi_1 _2273_ (.Y(_0583_),
    .B1(_0581_),
    .B2(_0536_),
    .A2(net404),
    .A1(net787));
 sg13g2_nor2_1 _2274_ (.A(net491),
    .B(net788),
    .Y(_0194_));
 sg13g2_a22oi_1 _2275_ (.Y(_0584_),
    .B1(_0581_),
    .B2(_0538_),
    .A2(net404),
    .A1(net700));
 sg13g2_nor2_1 _2276_ (.A(net491),
    .B(net701),
    .Y(_0195_));
 sg13g2_a22oi_1 _2277_ (.Y(_0585_),
    .B1(_0581_),
    .B2(_0540_),
    .A2(net404),
    .A1(net777));
 sg13g2_nor2_1 _2278_ (.A(net486),
    .B(net778),
    .Y(_0196_));
 sg13g2_nand2_2 _2279_ (.Y(_0586_),
    .A(_0467_),
    .B(net451));
 sg13g2_a22oi_1 _2280_ (.Y(_0587_),
    .B1(net418),
    .B2(net675),
    .A2(net425),
    .A1(_0469_));
 sg13g2_nor2_1 _2281_ (.A(net479),
    .B(_0587_),
    .Y(_0197_));
 sg13g2_a22oi_1 _2282_ (.Y(_0588_),
    .B1(net418),
    .B2(net635),
    .A2(net425),
    .A1(_0471_));
 sg13g2_nor2_1 _2283_ (.A(net479),
    .B(net636),
    .Y(_0198_));
 sg13g2_a22oi_1 _2284_ (.Y(_0589_),
    .B1(net418),
    .B2(net606),
    .A2(net425),
    .A1(_0473_));
 sg13g2_nor2_1 _2285_ (.A(net486),
    .B(_0589_),
    .Y(_0199_));
 sg13g2_o21ai_1 _2286_ (.B1(net512),
    .Y(_0590_),
    .A1(net455),
    .A2(net418));
 sg13g2_a21oi_1 _2287_ (.A1(_0837_),
    .A2(net418),
    .Y(_0200_),
    .B1(_0590_));
 sg13g2_a22oi_1 _2288_ (.Y(_0591_),
    .B1(net418),
    .B2(net673),
    .A2(_0581_),
    .A1(_0550_));
 sg13g2_nor2_1 _2289_ (.A(net483),
    .B(net674),
    .Y(_0201_));
 sg13g2_a22oi_1 _2290_ (.Y(_0592_),
    .B1(net418),
    .B2(net694),
    .A2(_0581_),
    .A1(_0552_));
 sg13g2_nor2_1 _2291_ (.A(net484),
    .B(net695),
    .Y(_0202_));
 sg13g2_a22oi_1 _2292_ (.Y(_0593_),
    .B1(net418),
    .B2(net649),
    .A2(_0581_),
    .A1(_0554_));
 sg13g2_nor2_1 _2293_ (.A(net484),
    .B(net650),
    .Y(_0203_));
 sg13g2_a22oi_1 _2294_ (.Y(_0594_),
    .B1(_0586_),
    .B2(net639),
    .A2(_0581_),
    .A1(_0556_));
 sg13g2_nor2_1 _2295_ (.A(net486),
    .B(net640),
    .Y(_0204_));
 sg13g2_nor2b_2 _2296_ (.A(_0314_),
    .B_N(_0333_),
    .Y(_0595_));
 sg13g2_nand2_2 _2297_ (.Y(_0596_),
    .A(_0319_),
    .B(net449));
 sg13g2_and2_1 _2298_ (.A(_0317_),
    .B(net449),
    .X(_0597_));
 sg13g2_a22oi_1 _2299_ (.Y(_0598_),
    .B1(net416),
    .B2(_0409_),
    .A2(_0596_),
    .A1(net742));
 sg13g2_nor2_1 _2300_ (.A(net472),
    .B(_0598_),
    .Y(_0205_));
 sg13g2_a22oi_1 _2301_ (.Y(_0599_),
    .B1(net416),
    .B2(_0411_),
    .A2(_0596_),
    .A1(net756));
 sg13g2_nor2_1 _2302_ (.A(net472),
    .B(_0599_),
    .Y(_0206_));
 sg13g2_a22oi_1 _2303_ (.Y(_0600_),
    .B1(net417),
    .B2(_0413_),
    .A2(_0596_),
    .A1(net726));
 sg13g2_nor2_1 _2304_ (.A(net475),
    .B(_0600_),
    .Y(_0207_));
 sg13g2_nand2_1 _2305_ (.Y(_0601_),
    .A(_0417_),
    .B(net449));
 sg13g2_a22oi_1 _2306_ (.Y(_0602_),
    .B1(_0601_),
    .B2(net623),
    .A2(net416),
    .A1(_0419_));
 sg13g2_nor2_1 _2307_ (.A(net471),
    .B(_0602_),
    .Y(_0208_));
 sg13g2_a22oi_1 _2308_ (.Y(_0603_),
    .B1(_0601_),
    .B2(net685),
    .A2(net416),
    .A1(_0421_));
 sg13g2_nor2_1 _2309_ (.A(net471),
    .B(_0603_),
    .Y(_0209_));
 sg13g2_a22oi_1 _2310_ (.Y(_0604_),
    .B1(_0601_),
    .B2(net608),
    .A2(net416),
    .A1(_0423_));
 sg13g2_nor2_1 _2311_ (.A(net471),
    .B(_0604_),
    .Y(_0210_));
 sg13g2_and2_1 _2312_ (.A(net456),
    .B(net449),
    .X(_0605_));
 sg13g2_nand2_1 _2313_ (.Y(_0606_),
    .A(net456),
    .B(net449));
 sg13g2_a21oi_1 _2314_ (.A1(net552),
    .A2(net458),
    .Y(_0607_),
    .B1(_0606_));
 sg13g2_o21ai_1 _2315_ (.B1(net494),
    .Y(_0608_),
    .A1(net1026),
    .A2(_0605_));
 sg13g2_nor2_1 _2316_ (.A(_0607_),
    .B(_0608_),
    .Y(_0211_));
 sg13g2_a21oi_1 _2317_ (.A1(net551),
    .A2(net458),
    .Y(_0609_),
    .B1(_0606_));
 sg13g2_o21ai_1 _2318_ (.B1(net496),
    .Y(_0610_),
    .A1(net978),
    .A2(_0605_));
 sg13g2_nor2_1 _2319_ (.A(_0609_),
    .B(_0610_),
    .Y(_0212_));
 sg13g2_a21oi_1 _2320_ (.A1(\model_byte[2] ),
    .A2(net458),
    .Y(_0611_),
    .B1(_0606_));
 sg13g2_o21ai_1 _2321_ (.B1(net496),
    .Y(_0612_),
    .A1(net960),
    .A2(_0605_));
 sg13g2_nor2_1 _2322_ (.A(_0611_),
    .B(_0612_),
    .Y(_0213_));
 sg13g2_nand2_1 _2323_ (.Y(_0613_),
    .A(_0438_),
    .B(net449));
 sg13g2_a22oi_1 _2324_ (.Y(_0614_),
    .B1(_0613_),
    .B2(net681),
    .A2(net450),
    .A1(_0440_));
 sg13g2_nor2_1 _2325_ (.A(net473),
    .B(net682),
    .Y(_0214_));
 sg13g2_a22oi_1 _2326_ (.Y(_0615_),
    .B1(_0613_),
    .B2(net665),
    .A2(net450),
    .A1(_0442_));
 sg13g2_nor2_1 _2327_ (.A(net474),
    .B(net666),
    .Y(_0215_));
 sg13g2_a22oi_1 _2328_ (.Y(_0616_),
    .B1(_0613_),
    .B2(net705),
    .A2(net450),
    .A1(_0444_));
 sg13g2_nor2_1 _2329_ (.A(net473),
    .B(net706),
    .Y(_0216_));
 sg13g2_nand2_1 _2330_ (.Y(_0617_),
    .A(_0449_),
    .B(net449));
 sg13g2_a22oi_1 _2331_ (.Y(_0618_),
    .B1(_0617_),
    .B2(net710),
    .A2(net416),
    .A1(_0451_));
 sg13g2_nor2_1 _2332_ (.A(net477),
    .B(_0618_),
    .Y(_0217_));
 sg13g2_a22oi_1 _2333_ (.Y(_0619_),
    .B1(_0617_),
    .B2(net683),
    .A2(net416),
    .A1(_0453_));
 sg13g2_nor2_1 _2334_ (.A(net478),
    .B(_0619_),
    .Y(_0218_));
 sg13g2_a22oi_1 _2335_ (.Y(_0620_),
    .B1(_0617_),
    .B2(net709),
    .A2(net416),
    .A1(_0455_));
 sg13g2_nor2_1 _2336_ (.A(net477),
    .B(_0620_),
    .Y(_0219_));
 sg13g2_nand2_1 _2337_ (.Y(_0621_),
    .A(_0458_),
    .B(net449));
 sg13g2_a22oi_1 _2338_ (.Y(_0622_),
    .B1(_0621_),
    .B2(net611),
    .A2(net417),
    .A1(_0460_));
 sg13g2_nor2_1 _2339_ (.A(net482),
    .B(_0622_),
    .Y(_0220_));
 sg13g2_a22oi_1 _2340_ (.Y(_0623_),
    .B1(_0621_),
    .B2(net624),
    .A2(net417),
    .A1(_0462_));
 sg13g2_nor2_1 _2341_ (.A(net477),
    .B(_0623_),
    .Y(_0221_));
 sg13g2_a22oi_1 _2342_ (.Y(_0624_),
    .B1(_0621_),
    .B2(net622),
    .A2(net417),
    .A1(_0464_));
 sg13g2_nor2_1 _2343_ (.A(net477),
    .B(_0624_),
    .Y(_0222_));
 sg13g2_nand2_1 _2344_ (.Y(_0625_),
    .A(_0467_),
    .B(net450));
 sg13g2_a22oi_1 _2345_ (.Y(_0626_),
    .B1(_0625_),
    .B2(net655),
    .A2(net417),
    .A1(_0469_));
 sg13g2_nor2_1 _2346_ (.A(net479),
    .B(_0626_),
    .Y(_0223_));
 sg13g2_a22oi_1 _2347_ (.Y(_0627_),
    .B1(_0625_),
    .B2(net696),
    .A2(net417),
    .A1(_0471_));
 sg13g2_nor2_1 _2348_ (.A(net479),
    .B(net697),
    .Y(_0224_));
 sg13g2_a22oi_1 _2349_ (.Y(_0628_),
    .B1(_0625_),
    .B2(net663),
    .A2(net417),
    .A1(_0473_));
 sg13g2_nor2_1 _2350_ (.A(net481),
    .B(_0628_),
    .Y(_0225_));
 sg13g2_a21oi_1 _2351_ (.A1(net920),
    .A2(_0596_),
    .Y(_0629_),
    .B1(net401));
 sg13g2_nor2_1 _2352_ (.A(net485),
    .B(_0629_),
    .Y(_0226_));
 sg13g2_o21ai_1 _2353_ (.B1(net514),
    .Y(_0630_),
    .A1(net586),
    .A2(\u_feature_loader.feature_idx_q[0] ));
 sg13g2_a21oi_1 _2354_ (.A1(net586),
    .A2(\u_feature_loader.feature_idx_q[0] ),
    .Y(_0227_),
    .B1(_0630_));
 sg13g2_a21oi_1 _2355_ (.A1(net586),
    .A2(\u_feature_loader.feature_idx_q[0] ),
    .Y(_0631_),
    .B1(net976));
 sg13g2_nor3_1 _2356_ (.A(net490),
    .B(_1145_),
    .C(net977),
    .Y(_0228_));
 sg13g2_o21ai_1 _2357_ (.B1(net513),
    .Y(_0632_),
    .A1(net544),
    .A2(_1145_));
 sg13g2_nor2b_1 _2358_ (.A(_0632_),
    .B_N(_1146_),
    .Y(_0229_));
 sg13g2_and3_1 _2359_ (.X(_0230_),
    .A(net643),
    .B(net513),
    .C(_1146_));
 sg13g2_o21ai_1 _2360_ (.B1(net497),
    .Y(_0633_),
    .A1(\feature_byte[0] ),
    .A2(net436));
 sg13g2_a21oi_1 _2361_ (.A1(_0836_),
    .A2(net436),
    .Y(_0231_),
    .B1(_0633_));
 sg13g2_o21ai_1 _2362_ (.B1(net497),
    .Y(_0634_),
    .A1(\feature_byte[1] ),
    .A2(net436));
 sg13g2_a21oi_1 _2363_ (.A1(_0835_),
    .A2(net436),
    .Y(_0232_),
    .B1(_0634_));
 sg13g2_o21ai_1 _2364_ (.B1(net497),
    .Y(_0635_),
    .A1(\feature_byte[2] ),
    .A2(net436));
 sg13g2_a21oi_1 _2365_ (.A1(_0834_),
    .A2(net436),
    .Y(_0233_),
    .B1(_0635_));
 sg13g2_o21ai_1 _2366_ (.B1(net497),
    .Y(_0636_),
    .A1(\feature_byte[3] ),
    .A2(net436));
 sg13g2_a21oi_1 _2367_ (.A1(_0833_),
    .A2(net436),
    .Y(_0234_),
    .B1(_0636_));
 sg13g2_o21ai_1 _2368_ (.B1(net513),
    .Y(_0637_),
    .A1(\feature_byte[4] ),
    .A2(net435));
 sg13g2_a21oi_1 _2369_ (.A1(_0832_),
    .A2(net435),
    .Y(_0235_),
    .B1(_0637_));
 sg13g2_o21ai_1 _2370_ (.B1(net513),
    .Y(_0638_),
    .A1(\feature_byte[5] ),
    .A2(net435));
 sg13g2_a21oi_1 _2371_ (.A1(_0831_),
    .A2(net435),
    .Y(_0236_),
    .B1(_0638_));
 sg13g2_o21ai_1 _2372_ (.B1(net511),
    .Y(_0639_),
    .A1(\feature_byte[6] ),
    .A2(net435));
 sg13g2_a21oi_1 _2373_ (.A1(_0830_),
    .A2(net435),
    .Y(_0237_),
    .B1(_0639_));
 sg13g2_o21ai_1 _2374_ (.B1(net513),
    .Y(_0640_),
    .A1(\feature_byte[7] ),
    .A2(net435));
 sg13g2_a21oi_1 _2375_ (.A1(_0829_),
    .A2(net435),
    .Y(_0238_),
    .B1(_0640_));
 sg13g2_nor2b_2 _2376_ (.A(\u_feature_loader.feature_idx_q[1] ),
    .B_N(\u_feature_loader.feature_idx_q[0] ),
    .Y(_0641_));
 sg13g2_nand3b_1 _2377_ (.B(_1149_),
    .C(net461),
    .Y(_0642_),
    .A_N(net543));
 sg13g2_and2_1 _2378_ (.A(\feature_byte[0] ),
    .B(net461),
    .X(_0643_));
 sg13g2_o21ai_1 _2379_ (.B1(net544),
    .Y(_0644_),
    .A1(\u_feature_loader.feature_idx_q[1] ),
    .A2(\u_feature_loader.feature_idx_q[0] ));
 sg13g2_nand2b_1 _2380_ (.Y(_0645_),
    .B(_0644_),
    .A_N(\u_feature_loader.feature_idx_q[3] ));
 sg13g2_nor3_2 _2381_ (.A(_0825_),
    .B(_1148_),
    .C(_0645_),
    .Y(_0646_));
 sg13g2_a22oi_1 _2382_ (.Y(_0647_),
    .B1(_0643_),
    .B2(net412),
    .A2(_0642_),
    .A1(net784));
 sg13g2_nor2_1 _2383_ (.A(net480),
    .B(net785),
    .Y(_0239_));
 sg13g2_and2_1 _2384_ (.A(\feature_byte[1] ),
    .B(net461),
    .X(_0648_));
 sg13g2_a22oi_1 _2385_ (.Y(_0649_),
    .B1(net412),
    .B2(_0648_),
    .A2(_0642_),
    .A1(net801));
 sg13g2_nor2_1 _2386_ (.A(net480),
    .B(net802),
    .Y(_0240_));
 sg13g2_and2_1 _2387_ (.A(\feature_byte[2] ),
    .B(net461),
    .X(_0650_));
 sg13g2_a22oi_1 _2388_ (.Y(_0651_),
    .B1(net412),
    .B2(_0650_),
    .A2(_0642_),
    .A1(net797));
 sg13g2_nor2_1 _2389_ (.A(net480),
    .B(net798),
    .Y(_0241_));
 sg13g2_and2_1 _2390_ (.A(\feature_byte[3] ),
    .B(net461),
    .X(_0652_));
 sg13g2_a22oi_1 _2391_ (.Y(_0653_),
    .B1(net413),
    .B2(_0652_),
    .A2(_0642_),
    .A1(net884));
 sg13g2_nor2_1 _2392_ (.A(net487),
    .B(net885),
    .Y(_0242_));
 sg13g2_and2_1 _2393_ (.A(\feature_byte[4] ),
    .B(net461),
    .X(_0654_));
 sg13g2_a22oi_1 _2394_ (.Y(_0655_),
    .B1(net414),
    .B2(_0654_),
    .A2(_0642_),
    .A1(net832));
 sg13g2_nor2_1 _2395_ (.A(net490),
    .B(net833),
    .Y(_0243_));
 sg13g2_and2_1 _2396_ (.A(\feature_byte[5] ),
    .B(net461),
    .X(_0656_));
 sg13g2_a22oi_1 _2397_ (.Y(_0657_),
    .B1(net414),
    .B2(_0656_),
    .A2(_0642_),
    .A1(net811));
 sg13g2_nor2_1 _2398_ (.A(net489),
    .B(net812),
    .Y(_0244_));
 sg13g2_and2_1 _2399_ (.A(\feature_byte[6] ),
    .B(_0641_),
    .X(_0658_));
 sg13g2_a22oi_1 _2400_ (.Y(_0659_),
    .B1(net415),
    .B2(_0658_),
    .A2(_0642_),
    .A1(net794));
 sg13g2_nor2_1 _2401_ (.A(net488),
    .B(net795),
    .Y(_0245_));
 sg13g2_and2_1 _2402_ (.A(\feature_byte[7] ),
    .B(_0641_),
    .X(_0660_));
 sg13g2_a22oi_1 _2403_ (.Y(_0661_),
    .B1(net414),
    .B2(_0660_),
    .A2(_0642_),
    .A1(net799));
 sg13g2_nor2_1 _2404_ (.A(net489),
    .B(net800),
    .Y(_0246_));
 sg13g2_nor2b_2 _2405_ (.A(\u_feature_loader.feature_idx_q[0] ),
    .B_N(\u_feature_loader.feature_idx_q[1] ),
    .Y(_0662_));
 sg13g2_and2_1 _2406_ (.A(net415),
    .B(_0662_),
    .X(_0663_));
 sg13g2_nand2_2 _2407_ (.Y(_0664_),
    .A(net414),
    .B(_0662_));
 sg13g2_a21oi_1 _2408_ (.A1(\feature_byte[0] ),
    .A2(net459),
    .Y(_0665_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2409_ (.B1(net497),
    .Y(_0666_),
    .A1(net974),
    .A2(_0663_));
 sg13g2_nor2_1 _2410_ (.A(_0665_),
    .B(_0666_),
    .Y(_0247_));
 sg13g2_a21oi_1 _2411_ (.A1(\feature_byte[1] ),
    .A2(net459),
    .Y(_0667_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2412_ (.B1(net497),
    .Y(_0668_),
    .A1(net899),
    .A2(_0663_));
 sg13g2_nor2_1 _2413_ (.A(_0667_),
    .B(_0668_),
    .Y(_0248_));
 sg13g2_a21oi_1 _2414_ (.A1(\feature_byte[2] ),
    .A2(net459),
    .Y(_0669_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2415_ (.B1(net497),
    .Y(_0670_),
    .A1(net1011),
    .A2(_0663_));
 sg13g2_nor2_1 _2416_ (.A(_0669_),
    .B(_0670_),
    .Y(_0249_));
 sg13g2_a21oi_1 _2417_ (.A1(\feature_byte[3] ),
    .A2(net459),
    .Y(_0671_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2418_ (.B1(net498),
    .Y(_0672_),
    .A1(net988),
    .A2(_0663_));
 sg13g2_nor2_1 _2419_ (.A(_0671_),
    .B(_0672_),
    .Y(_0250_));
 sg13g2_a21oi_1 _2420_ (.A1(\feature_byte[4] ),
    .A2(net460),
    .Y(_0673_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2421_ (.B1(net513),
    .Y(_0674_),
    .A1(net952),
    .A2(_0663_));
 sg13g2_nor2_1 _2422_ (.A(_0673_),
    .B(_0674_),
    .Y(_0251_));
 sg13g2_a21oi_1 _2423_ (.A1(\feature_byte[5] ),
    .A2(net460),
    .Y(_0675_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2424_ (.B1(net513),
    .Y(_0676_),
    .A1(net912),
    .A2(_0663_));
 sg13g2_nor2_1 _2425_ (.A(_0675_),
    .B(_0676_),
    .Y(_0252_));
 sg13g2_a21oi_1 _2426_ (.A1(\feature_byte[6] ),
    .A2(net460),
    .Y(_0677_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2427_ (.B1(net511),
    .Y(_0678_),
    .A1(net994),
    .A2(_0663_));
 sg13g2_nor2_1 _2428_ (.A(_0677_),
    .B(_0678_),
    .Y(_0253_));
 sg13g2_a21oi_1 _2429_ (.A1(\feature_byte[7] ),
    .A2(net460),
    .Y(_0679_),
    .B1(_0664_));
 sg13g2_o21ai_1 _2430_ (.B1(net513),
    .Y(_0680_),
    .A1(net950),
    .A2(_0663_));
 sg13g2_nor2_1 _2431_ (.A(_0679_),
    .B(_0680_),
    .Y(_0254_));
 sg13g2_nand2_2 _2432_ (.Y(_0681_),
    .A(net462),
    .B(net413));
 sg13g2_and2_1 _2433_ (.A(\feature_byte[0] ),
    .B(net462),
    .X(_0682_));
 sg13g2_a22oi_1 _2434_ (.Y(_0683_),
    .B1(_0682_),
    .B2(net412),
    .A2(_0681_),
    .A1(net869));
 sg13g2_nor2_1 _2435_ (.A(net480),
    .B(net870),
    .Y(_0255_));
 sg13g2_and2_1 _2436_ (.A(\feature_byte[1] ),
    .B(net462),
    .X(_0684_));
 sg13g2_a22oi_1 _2437_ (.Y(_0685_),
    .B1(_0684_),
    .B2(net412),
    .A2(_0681_),
    .A1(net892));
 sg13g2_nor2_1 _2438_ (.A(net480),
    .B(net893),
    .Y(_0256_));
 sg13g2_and2_1 _2439_ (.A(\feature_byte[2] ),
    .B(net462),
    .X(_0686_));
 sg13g2_a22oi_1 _2440_ (.Y(_0687_),
    .B1(_0686_),
    .B2(net412),
    .A2(_0681_),
    .A1(net808));
 sg13g2_nor2_1 _2441_ (.A(net479),
    .B(net809),
    .Y(_0257_));
 sg13g2_and2_1 _2442_ (.A(\feature_byte[3] ),
    .B(net462),
    .X(_0688_));
 sg13g2_a22oi_1 _2443_ (.Y(_0689_),
    .B1(_0688_),
    .B2(net413),
    .A2(_0681_),
    .A1(net791));
 sg13g2_nor2_1 _2444_ (.A(net487),
    .B(net792),
    .Y(_0258_));
 sg13g2_and2_1 _2445_ (.A(\feature_byte[4] ),
    .B(net462),
    .X(_0690_));
 sg13g2_a22oi_1 _2446_ (.Y(_0691_),
    .B1(_0690_),
    .B2(net414),
    .A2(_0681_),
    .A1(net743));
 sg13g2_nor2_1 _2447_ (.A(net491),
    .B(net744),
    .Y(_0259_));
 sg13g2_and2_1 _2448_ (.A(\feature_byte[5] ),
    .B(net462),
    .X(_0692_));
 sg13g2_a22oi_1 _2449_ (.Y(_0693_),
    .B1(_0692_),
    .B2(net414),
    .A2(_0681_),
    .A1(net814));
 sg13g2_nor2_1 _2450_ (.A(net489),
    .B(net815),
    .Y(_0260_));
 sg13g2_and2_1 _2451_ (.A(\feature_byte[6] ),
    .B(net462),
    .X(_0694_));
 sg13g2_a22oi_1 _2452_ (.Y(_0695_),
    .B1(_0694_),
    .B2(net415),
    .A2(_0681_),
    .A1(net734));
 sg13g2_nor2_1 _2453_ (.A(net488),
    .B(net735),
    .Y(_0261_));
 sg13g2_and2_1 _2454_ (.A(\feature_byte[7] ),
    .B(_1144_),
    .X(_0696_));
 sg13g2_a22oi_1 _2455_ (.Y(_0697_),
    .B1(_0696_),
    .B2(net414),
    .A2(_0681_),
    .A1(net874));
 sg13g2_nor2_1 _2456_ (.A(net490),
    .B(net875),
    .Y(_0262_));
 sg13g2_nand2_2 _2457_ (.Y(_0698_),
    .A(net543),
    .B(net413));
 sg13g2_nand2_1 _2458_ (.Y(_0699_),
    .A(net571),
    .B(_0698_));
 sg13g2_nand3_1 _2459_ (.B(\feature_byte[0] ),
    .C(net412),
    .A(net543),
    .Y(_0700_));
 sg13g2_a21oi_1 _2460_ (.A1(_0699_),
    .A2(_0700_),
    .Y(_0263_),
    .B1(net487));
 sg13g2_nand2_1 _2461_ (.Y(_0701_),
    .A(net364),
    .B(_0698_));
 sg13g2_nand3_1 _2462_ (.B(\feature_byte[1] ),
    .C(net412),
    .A(net543),
    .Y(_0702_));
 sg13g2_a21oi_1 _2463_ (.A1(_0701_),
    .A2(_0702_),
    .Y(_0264_),
    .B1(net480));
 sg13g2_nand2_1 _2464_ (.Y(_0703_),
    .A(net579),
    .B(_0698_));
 sg13g2_nand3_1 _2465_ (.B(\feature_byte[2] ),
    .C(net413),
    .A(net543),
    .Y(_0704_));
 sg13g2_a21oi_1 _2466_ (.A1(_0703_),
    .A2(_0704_),
    .Y(_0265_),
    .B1(net487));
 sg13g2_nand2_1 _2467_ (.Y(_0705_),
    .A(net573),
    .B(_0698_));
 sg13g2_nand3_1 _2468_ (.B(\feature_byte[3] ),
    .C(net413),
    .A(net543),
    .Y(_0706_));
 sg13g2_a21oi_1 _2469_ (.A1(_0705_),
    .A2(_0706_),
    .Y(_0266_),
    .B1(net487));
 sg13g2_nand2_1 _2470_ (.Y(_0707_),
    .A(net575),
    .B(_0698_));
 sg13g2_nand3_1 _2471_ (.B(\feature_byte[4] ),
    .C(net414),
    .A(net544),
    .Y(_0708_));
 sg13g2_a21oi_1 _2472_ (.A1(_0707_),
    .A2(_0708_),
    .Y(_0267_),
    .B1(net489));
 sg13g2_nand2_1 _2473_ (.Y(_0709_),
    .A(net361),
    .B(_0698_));
 sg13g2_nand3_1 _2474_ (.B(\feature_byte[5] ),
    .C(net415),
    .A(net543),
    .Y(_0710_));
 sg13g2_a21oi_1 _2475_ (.A1(_0709_),
    .A2(_0710_),
    .Y(_0268_),
    .B1(net488));
 sg13g2_nand2_1 _2476_ (.Y(_0711_),
    .A(net583),
    .B(_0698_));
 sg13g2_nand3_1 _2477_ (.B(\feature_byte[6] ),
    .C(net415),
    .A(net543),
    .Y(_0712_));
 sg13g2_a21oi_1 _2478_ (.A1(_0711_),
    .A2(_0712_),
    .Y(_0269_),
    .B1(net487));
 sg13g2_nand2_1 _2479_ (.Y(_0713_),
    .A(net557),
    .B(_0698_));
 sg13g2_nand3_1 _2480_ (.B(\feature_byte[7] ),
    .C(net415),
    .A(net544),
    .Y(_0714_));
 sg13g2_a21oi_1 _2481_ (.A1(_0713_),
    .A2(_0714_),
    .Y(_0270_),
    .B1(net489));
 sg13g2_nand2b_1 _2482_ (.Y(_0715_),
    .B(\u_feature_loader.feature_idx_q[3] ),
    .A_N(_1148_));
 sg13g2_and3_1 _2483_ (.X(_0716_),
    .A(net586),
    .B(_0645_),
    .C(_0715_));
 sg13g2_nand2_2 _2484_ (.Y(_0717_),
    .A(net461),
    .B(net411));
 sg13g2_a22oi_1 _2485_ (.Y(_0718_),
    .B1(_0717_),
    .B2(net652),
    .A2(net409),
    .A1(_0643_));
 sg13g2_nor2_1 _2486_ (.A(net481),
    .B(net653),
    .Y(_0271_));
 sg13g2_a22oi_1 _2487_ (.Y(_0719_),
    .B1(_0717_),
    .B2(net625),
    .A2(net409),
    .A1(_0648_));
 sg13g2_nor2_1 _2488_ (.A(net480),
    .B(net626),
    .Y(_0272_));
 sg13g2_a22oi_1 _2489_ (.Y(_0720_),
    .B1(_0717_),
    .B2(net703),
    .A2(net409),
    .A1(_0650_));
 sg13g2_nor2_1 _2490_ (.A(net479),
    .B(net704),
    .Y(_0273_));
 sg13g2_a22oi_1 _2491_ (.Y(_0721_),
    .B1(_0717_),
    .B2(net645),
    .A2(net411),
    .A1(_0652_));
 sg13g2_nor2_1 _2492_ (.A(net487),
    .B(net646),
    .Y(_0274_));
 sg13g2_a22oi_1 _2493_ (.Y(_0722_),
    .B1(_0717_),
    .B2(net676),
    .A2(net411),
    .A1(_0654_));
 sg13g2_nor2_1 _2494_ (.A(net489),
    .B(net677),
    .Y(_0275_));
 sg13g2_a22oi_1 _2495_ (.Y(_0723_),
    .B1(_0717_),
    .B2(net656),
    .A2(net410),
    .A1(_0656_));
 sg13g2_nor2_1 _2496_ (.A(net488),
    .B(net657),
    .Y(_0276_));
 sg13g2_a22oi_1 _2497_ (.Y(_0724_),
    .B1(_0717_),
    .B2(net619),
    .A2(net410),
    .A1(_0658_));
 sg13g2_nor2_1 _2498_ (.A(net488),
    .B(net620),
    .Y(_0277_));
 sg13g2_a22oi_1 _2499_ (.Y(_0725_),
    .B1(_0717_),
    .B2(net633),
    .A2(net410),
    .A1(_0660_));
 sg13g2_nor2_1 _2500_ (.A(net489),
    .B(net634),
    .Y(_0278_));
 sg13g2_and2_1 _2501_ (.A(_0662_),
    .B(net410),
    .X(_0726_));
 sg13g2_nand2_2 _2502_ (.Y(_0727_),
    .A(_0662_),
    .B(net410));
 sg13g2_a21oi_1 _2503_ (.A1(\feature_byte[0] ),
    .A2(net459),
    .Y(_0728_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2504_ (.B1(net511),
    .Y(_0729_),
    .A1(net1013),
    .A2(_0726_));
 sg13g2_nor2_1 _2505_ (.A(_0728_),
    .B(_0729_),
    .Y(_0279_));
 sg13g2_a21oi_1 _2506_ (.A1(\feature_byte[1] ),
    .A2(net459),
    .Y(_0730_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2507_ (.B1(net497),
    .Y(_0731_),
    .A1(net849),
    .A2(_0726_));
 sg13g2_nor2_1 _2508_ (.A(_0730_),
    .B(_0731_),
    .Y(_0280_));
 sg13g2_a21oi_1 _2509_ (.A1(\feature_byte[2] ),
    .A2(net459),
    .Y(_0732_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2510_ (.B1(net511),
    .Y(_0733_),
    .A1(net964),
    .A2(_0726_));
 sg13g2_nor2_1 _2511_ (.A(_0732_),
    .B(_0733_),
    .Y(_0281_));
 sg13g2_a21oi_1 _2512_ (.A1(\feature_byte[3] ),
    .A2(net459),
    .Y(_0734_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2513_ (.B1(net511),
    .Y(_0735_),
    .A1(net922),
    .A2(_0726_));
 sg13g2_nor2_1 _2514_ (.A(_0734_),
    .B(_0735_),
    .Y(_0282_));
 sg13g2_a21oi_1 _2515_ (.A1(\feature_byte[4] ),
    .A2(net460),
    .Y(_0736_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2516_ (.B1(net515),
    .Y(_0737_),
    .A1(net997),
    .A2(_0726_));
 sg13g2_nor2_1 _2517_ (.A(_0736_),
    .B(net998),
    .Y(_0283_));
 sg13g2_a21oi_1 _2518_ (.A1(\feature_byte[5] ),
    .A2(net460),
    .Y(_0738_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2519_ (.B1(net511),
    .Y(_0739_),
    .A1(net858),
    .A2(_0726_));
 sg13g2_nor2_1 _2520_ (.A(_0738_),
    .B(_0739_),
    .Y(_0284_));
 sg13g2_a21oi_1 _2521_ (.A1(\feature_byte[6] ),
    .A2(net460),
    .Y(_0740_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2522_ (.B1(net511),
    .Y(_0741_),
    .A1(net1028),
    .A2(_0726_));
 sg13g2_nor2_1 _2523_ (.A(_0740_),
    .B(_0741_),
    .Y(_0285_));
 sg13g2_a21oi_1 _2524_ (.A1(\feature_byte[7] ),
    .A2(net460),
    .Y(_0742_),
    .B1(_0727_));
 sg13g2_o21ai_1 _2525_ (.B1(net511),
    .Y(_0743_),
    .A1(net816),
    .A2(_0726_));
 sg13g2_nor2_1 _2526_ (.A(_0742_),
    .B(_0743_),
    .Y(_0286_));
 sg13g2_a22oi_1 _2527_ (.Y(_0744_),
    .B1(_0682_),
    .B2(net409),
    .A2(net406),
    .A1(net862));
 sg13g2_nor2_1 _2528_ (.A(net481),
    .B(net863),
    .Y(_0287_));
 sg13g2_a22oi_1 _2529_ (.Y(_0745_),
    .B1(_0684_),
    .B2(net409),
    .A2(net406),
    .A1(net916));
 sg13g2_nor2_1 _2530_ (.A(net480),
    .B(net917),
    .Y(_0288_));
 sg13g2_a22oi_1 _2531_ (.Y(_0746_),
    .B1(_0686_),
    .B2(net409),
    .A2(net406),
    .A1(net771));
 sg13g2_nor2_1 _2532_ (.A(net488),
    .B(net772),
    .Y(_0289_));
 sg13g2_a22oi_1 _2533_ (.Y(_0747_),
    .B1(_0688_),
    .B2(net409),
    .A2(net406),
    .A1(net763));
 sg13g2_nor2_1 _2534_ (.A(net487),
    .B(net764),
    .Y(_0290_));
 sg13g2_a22oi_1 _2535_ (.Y(_0748_),
    .B1(_0690_),
    .B2(net410),
    .A2(net406),
    .A1(net718));
 sg13g2_nor2_1 _2536_ (.A(net491),
    .B(net719),
    .Y(_0291_));
 sg13g2_a22oi_1 _2537_ (.Y(_0749_),
    .B1(_0692_),
    .B2(net410),
    .A2(net406),
    .A1(net750));
 sg13g2_nor2_1 _2538_ (.A(net489),
    .B(net751),
    .Y(_0292_));
 sg13g2_a22oi_1 _2539_ (.Y(_0750_),
    .B1(_0694_),
    .B2(net409),
    .A2(net406),
    .A1(net715));
 sg13g2_nor2_1 _2540_ (.A(net488),
    .B(net716),
    .Y(_0293_));
 sg13g2_a22oi_1 _2541_ (.Y(_0751_),
    .B1(_0696_),
    .B2(net410),
    .A2(_1147_),
    .A1(net754));
 sg13g2_nor2_1 _2542_ (.A(net490),
    .B(net755),
    .Y(_0294_));
 sg13g2_and4_1 _2543_ (.A(net3),
    .B(net554),
    .C(net12),
    .D(_1125_),
    .X(_0295_));
 sg13g2_nor2_1 _2544_ (.A(net688),
    .B(_1116_),
    .Y(_0752_));
 sg13g2_nor2b_1 _2545_ (.A(net689),
    .B_N(_0001_),
    .Y(_0296_));
 sg13g2_xnor2_1 _2546_ (.Y(_0753_),
    .A(_1088_),
    .B(_1112_));
 sg13g2_xnor2_1 _2547_ (.Y(_0754_),
    .A(_1087_),
    .B(_1112_));
 sg13g2_a21oi_1 _2548_ (.A1(_1095_),
    .A2(_1100_),
    .Y(_0755_),
    .B1(net380));
 sg13g2_mux4_1 _2549_ (.S0(net379),
    .A0(\leaf_value_flat[24] ),
    .A1(\leaf_value_flat[8] ),
    .A2(\leaf_value_flat[0] ),
    .A3(\leaf_value_flat[16] ),
    .S1(net382),
    .X(_0756_));
 sg13g2_or2_1 _2550_ (.X(_0757_),
    .B(_0756_),
    .A(_0753_));
 sg13g2_mux4_1 _2551_ (.S0(net379),
    .A0(\leaf_value_flat[56] ),
    .A1(\leaf_value_flat[40] ),
    .A2(\leaf_value_flat[32] ),
    .A3(\leaf_value_flat[48] ),
    .S1(net382),
    .X(_0758_));
 sg13g2_nand2b_1 _2552_ (.Y(_0759_),
    .B(_0753_),
    .A_N(_0758_));
 sg13g2_nand3_1 _2553_ (.B(_1087_),
    .C(_1112_),
    .A(_1075_),
    .Y(_0760_));
 sg13g2_and3_2 _2554_ (.X(_0761_),
    .A(_1113_),
    .B(_1114_),
    .C(_0760_));
 sg13g2_nand3_1 _2555_ (.B(_1114_),
    .C(_0760_),
    .A(_1113_),
    .Y(_0762_));
 sg13g2_nand3_1 _2556_ (.B(_0759_),
    .C(_0761_),
    .A(_0757_),
    .Y(_0763_));
 sg13g2_nand2_1 _2557_ (.Y(_0764_),
    .A(net845),
    .B(net508));
 sg13g2_a22oi_1 _2558_ (.Y(_0297_),
    .B1(_0764_),
    .B2(net376),
    .A2(_0763_),
    .A1(net377));
 sg13g2_mux4_1 _2559_ (.S0(net379),
    .A0(\leaf_value_flat[25] ),
    .A1(\leaf_value_flat[9] ),
    .A2(\leaf_value_flat[1] ),
    .A3(\leaf_value_flat[17] ),
    .S1(net380),
    .X(_0765_));
 sg13g2_mux4_1 _2560_ (.S0(net379),
    .A0(\leaf_value_flat[57] ),
    .A1(\leaf_value_flat[41] ),
    .A2(\leaf_value_flat[33] ),
    .A3(\leaf_value_flat[49] ),
    .S1(net380),
    .X(_0766_));
 sg13g2_mux2_1 _2561_ (.A0(_0765_),
    .A1(_0766_),
    .S(_0753_),
    .X(_0767_));
 sg13g2_nand2_1 _2562_ (.Y(_0768_),
    .A(_0761_),
    .B(_0767_));
 sg13g2_nand2_1 _2563_ (.Y(_0769_),
    .A(net729),
    .B(net508));
 sg13g2_a22oi_1 _2564_ (.Y(_0298_),
    .B1(_0769_),
    .B2(net376),
    .A2(_0768_),
    .A1(net377));
 sg13g2_mux4_1 _2565_ (.S0(net379),
    .A0(\leaf_value_flat[58] ),
    .A1(\leaf_value_flat[42] ),
    .A2(\leaf_value_flat[34] ),
    .A3(\leaf_value_flat[50] ),
    .S1(net380),
    .X(_0770_));
 sg13g2_mux4_1 _2566_ (.S0(net379),
    .A0(\leaf_value_flat[26] ),
    .A1(\leaf_value_flat[10] ),
    .A2(\leaf_value_flat[2] ),
    .A3(\leaf_value_flat[18] ),
    .S1(net380),
    .X(_0771_));
 sg13g2_mux2_1 _2567_ (.A0(_0770_),
    .A1(_0771_),
    .S(_0754_),
    .X(_0772_));
 sg13g2_nand2_1 _2568_ (.Y(_0773_),
    .A(_0761_),
    .B(_0772_));
 sg13g2_nand2_1 _2569_ (.Y(_0774_),
    .A(net748),
    .B(net508));
 sg13g2_a22oi_1 _2570_ (.Y(_0299_),
    .B1(_0774_),
    .B2(net376),
    .A2(_0773_),
    .A1(net377));
 sg13g2_mux2_1 _2571_ (.A0(\leaf_value_flat[59] ),
    .A1(\leaf_value_flat[51] ),
    .S(net380),
    .X(_0775_));
 sg13g2_or3_1 _2572_ (.A(_1112_),
    .B(_0755_),
    .C(_0775_),
    .X(_0776_));
 sg13g2_a22oi_1 _2573_ (.Y(_0777_),
    .B1(_0755_),
    .B2(_0883_),
    .A2(_1088_),
    .A1(_0884_));
 sg13g2_a21oi_1 _2574_ (.A1(_0776_),
    .A2(_0777_),
    .Y(_0778_),
    .B1(_0754_));
 sg13g2_mux4_1 _2575_ (.S0(net379),
    .A0(\leaf_value_flat[27] ),
    .A1(\leaf_value_flat[11] ),
    .A2(\leaf_value_flat[3] ),
    .A3(\leaf_value_flat[19] ),
    .S1(net380),
    .X(_0779_));
 sg13g2_nor2_1 _2576_ (.A(_0753_),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_or3_1 _2577_ (.A(_0762_),
    .B(_0778_),
    .C(_0780_),
    .X(_0781_));
 sg13g2_nand2_1 _2578_ (.Y(_0782_),
    .A(net818),
    .B(net508));
 sg13g2_a22oi_1 _2579_ (.Y(_0300_),
    .B1(_0782_),
    .B2(net376),
    .A2(_0781_),
    .A1(_1153_));
 sg13g2_mux4_1 _2580_ (.S0(net378),
    .A0(\leaf_value_flat[28] ),
    .A1(\leaf_value_flat[12] ),
    .A2(\leaf_value_flat[4] ),
    .A3(\leaf_value_flat[20] ),
    .S1(net381),
    .X(_0783_));
 sg13g2_mux4_1 _2581_ (.S0(net378),
    .A0(\leaf_value_flat[60] ),
    .A1(\leaf_value_flat[44] ),
    .A2(\leaf_value_flat[36] ),
    .A3(\leaf_value_flat[52] ),
    .S1(net381),
    .X(_0784_));
 sg13g2_mux2_1 _2582_ (.A0(_0783_),
    .A1(_0784_),
    .S(_0753_),
    .X(_0785_));
 sg13g2_nand2_1 _2583_ (.Y(_0786_),
    .A(_0761_),
    .B(_0785_));
 sg13g2_nand2_1 _2584_ (.Y(_0787_),
    .A(net698),
    .B(net508));
 sg13g2_a22oi_1 _2585_ (.Y(_0301_),
    .B1(_0787_),
    .B2(net376),
    .A2(_0786_),
    .A1(net377));
 sg13g2_mux4_1 _2586_ (.S0(_1101_),
    .A0(\leaf_value_flat[29] ),
    .A1(\leaf_value_flat[13] ),
    .A2(\leaf_value_flat[5] ),
    .A3(\leaf_value_flat[21] ),
    .S1(net381),
    .X(_0788_));
 sg13g2_mux4_1 _2587_ (.S0(net378),
    .A0(\leaf_value_flat[61] ),
    .A1(\leaf_value_flat[45] ),
    .A2(\leaf_value_flat[37] ),
    .A3(\leaf_value_flat[53] ),
    .S1(net381),
    .X(_0789_));
 sg13g2_mux2_1 _2588_ (.A0(_0788_),
    .A1(_0789_),
    .S(_0753_),
    .X(_0790_));
 sg13g2_nand2_1 _2589_ (.Y(_0791_),
    .A(_0761_),
    .B(_0790_));
 sg13g2_nand2_1 _2590_ (.Y(_0792_),
    .A(net723),
    .B(net509));
 sg13g2_a22oi_1 _2591_ (.Y(_0302_),
    .B1(_0792_),
    .B2(net376),
    .A2(_0791_),
    .A1(net377));
 sg13g2_mux4_1 _2592_ (.S0(net378),
    .A0(\leaf_value_flat[62] ),
    .A1(\leaf_value_flat[46] ),
    .A2(\leaf_value_flat[38] ),
    .A3(\leaf_value_flat[54] ),
    .S1(net382),
    .X(_0793_));
 sg13g2_mux4_1 _2593_ (.S0(net378),
    .A0(\leaf_value_flat[30] ),
    .A1(\leaf_value_flat[14] ),
    .A2(\leaf_value_flat[6] ),
    .A3(\leaf_value_flat[22] ),
    .S1(net381),
    .X(_0794_));
 sg13g2_mux2_1 _2594_ (.A0(_0793_),
    .A1(_0794_),
    .S(_0754_),
    .X(_0795_));
 sg13g2_nand2_1 _2595_ (.Y(_0796_),
    .A(_0761_),
    .B(_0795_));
 sg13g2_nand2_1 _2596_ (.Y(_0797_),
    .A(net761),
    .B(net508));
 sg13g2_a22oi_1 _2597_ (.Y(_0303_),
    .B1(_0797_),
    .B2(_1154_),
    .A2(_0796_),
    .A1(net377));
 sg13g2_mux4_1 _2598_ (.S0(net378),
    .A0(\leaf_value_flat[63] ),
    .A1(\leaf_value_flat[47] ),
    .A2(\leaf_value_flat[39] ),
    .A3(\leaf_value_flat[55] ),
    .S1(net381),
    .X(_0798_));
 sg13g2_mux4_1 _2599_ (.S0(net378),
    .A0(\leaf_value_flat[31] ),
    .A1(\leaf_value_flat[15] ),
    .A2(\leaf_value_flat[7] ),
    .A3(\leaf_value_flat[23] ),
    .S1(net381),
    .X(_0799_));
 sg13g2_mux2_1 _2600_ (.A0(_0798_),
    .A1(_0799_),
    .S(_0754_),
    .X(_0800_));
 sg13g2_nand2_1 _2601_ (.Y(_0801_),
    .A(_0761_),
    .B(_0800_));
 sg13g2_nand2_1 _2602_ (.Y(_0802_),
    .A(net691),
    .B(net508));
 sg13g2_a22oi_1 _2603_ (.Y(_0304_),
    .B1(_0802_),
    .B2(net376),
    .A2(_0801_),
    .A1(net377));
 sg13g2_o21ai_1 _2604_ (.B1(_1121_),
    .Y(_0803_),
    .A1(_1113_),
    .A2(_1115_));
 sg13g2_nand2_1 _2605_ (.Y(_0804_),
    .A(\u_tree_core.state_q[1] ),
    .B(_0902_));
 sg13g2_o21ai_1 _2606_ (.B1(_0804_),
    .Y(_0805_),
    .A1(_0902_),
    .A2(_1117_));
 sg13g2_a21oi_1 _2607_ (.A1(\u_tree_core.state_q[1] ),
    .A2(_0762_),
    .Y(_0806_),
    .B1(_0803_));
 sg13g2_a221oi_1 _2608_ (.B2(_0806_),
    .C1(net485),
    .B1(_0805_),
    .A1(_0823_),
    .Y(_0305_),
    .A2(_0803_));
 sg13g2_and2_1 _2609_ (.A(_1118_),
    .B(_0804_),
    .X(_0807_));
 sg13g2_a221oi_1 _2610_ (.B2(_0804_),
    .C1(_1120_),
    .B1(_1118_),
    .A1(\u_tree_core.state_q[1] ),
    .Y(_0808_),
    .A2(_1113_));
 sg13g2_nand2b_1 _2611_ (.Y(_0809_),
    .B(\u_tree_core.state_q[1] ),
    .A_N(net1041));
 sg13g2_o21ai_1 _2612_ (.B1(net509),
    .Y(_0810_),
    .A1(net1041),
    .A2(_0808_));
 sg13g2_a21oi_1 _2613_ (.A1(_0808_),
    .A2(_0809_),
    .Y(_0306_),
    .B1(_0810_));
 sg13g2_and3_1 _2614_ (.X(_0811_),
    .A(net593),
    .B(_0808_),
    .C(_0809_));
 sg13g2_nor3_2 _2615_ (.A(_1113_),
    .B(_1115_),
    .C(_0807_),
    .Y(_0812_));
 sg13g2_a21oi_1 _2616_ (.A1(\u_tree_core.depth_q[0] ),
    .A2(_0812_),
    .Y(_0813_),
    .B1(net593));
 sg13g2_nor3_1 _2617_ (.A(net485),
    .B(_0811_),
    .C(net594),
    .Y(_0307_));
 sg13g2_nand2b_1 _2618_ (.Y(_0814_),
    .B(net541),
    .A_N(_0808_));
 sg13g2_nand2_1 _2619_ (.Y(_0815_),
    .A(net381),
    .B(_0812_));
 sg13g2_a21oi_1 _2620_ (.A1(_0814_),
    .A2(_0815_),
    .Y(_0308_),
    .B1(net485));
 sg13g2_nand2b_1 _2621_ (.Y(_0816_),
    .B(net534),
    .A_N(_0808_));
 sg13g2_nand2b_1 _2622_ (.Y(_0817_),
    .B(_0812_),
    .A_N(net378));
 sg13g2_a21oi_1 _2623_ (.A1(_0816_),
    .A2(_0817_),
    .Y(_0309_),
    .B1(net485));
 sg13g2_nand2b_1 _2624_ (.Y(_0818_),
    .B(net533),
    .A_N(_0808_));
 sg13g2_nand2_1 _2625_ (.Y(_0819_),
    .A(_1087_),
    .B(_0812_));
 sg13g2_a21oi_1 _2626_ (.A1(_0818_),
    .A2(_0819_),
    .Y(_0310_),
    .B1(net485));
 sg13g2_dfrbpq_1 _2627_ (.RESET_B(net312),
    .D(_0002_),
    .Q(run_cmd),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _2628_ (.RESET_B(net201),
    .D(_0003_),
    .Q(feature_byte_valid),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2629_ (.RESET_B(net200),
    .D(_0004_),
    .Q(\feature_byte[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2630_ (.RESET_B(net198),
    .D(_0005_),
    .Q(\feature_byte[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2631_ (.RESET_B(net196),
    .D(_0006_),
    .Q(\feature_byte[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2632_ (.RESET_B(net194),
    .D(_0007_),
    .Q(\feature_byte[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _2633_ (.RESET_B(net192),
    .D(_0008_),
    .Q(\feature_byte[4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2634_ (.RESET_B(net190),
    .D(_0009_),
    .Q(\feature_byte[5] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _2635_ (.RESET_B(net188),
    .D(_0010_),
    .Q(\feature_byte[6] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2636_ (.RESET_B(net186),
    .D(_0011_),
    .Q(\feature_byte[7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2637_ (.RESET_B(net184),
    .D(_0012_),
    .Q(model_byte_valid),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _2638_ (.RESET_B(net183),
    .D(_0013_),
    .Q(\model_byte[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _2639_ (.RESET_B(net181),
    .D(_0014_),
    .Q(\model_byte[1] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2640_ (.RESET_B(net179),
    .D(_0015_),
    .Q(\model_byte[2] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2641_ (.RESET_B(net177),
    .D(_0016_),
    .Q(\model_byte[3] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _2642_ (.RESET_B(net175),
    .D(_0017_),
    .Q(\model_byte[4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _2643_ (.RESET_B(net173),
    .D(_0018_),
    .Q(\model_byte[5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _2644_ (.RESET_B(net171),
    .D(_0019_),
    .Q(\model_byte[6] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _2645_ (.RESET_B(net169),
    .D(_0020_),
    .Q(\model_byte[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _2646_ (.RESET_B(net167),
    .D(net1021),
    .Q(features_loaded),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2647_ (.RESET_B(net166),
    .D(_0022_),
    .Q(pred_valid),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2648_ (.RESET_B(net165),
    .D(net562),
    .Q(\u_model_loader.byte_idx_q[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _2649_ (.RESET_B(net163),
    .D(net882),
    .Q(\u_model_loader.byte_idx_q[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _2650_ (.RESET_B(net161),
    .D(_0025_),
    .Q(\u_model_loader.byte_idx_q[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _2651_ (.RESET_B(net159),
    .D(net1038),
    .Q(\u_model_loader.byte_idx_q[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _2652_ (.RESET_B(net157),
    .D(net1074),
    .Q(\u_model_loader.byte_idx_q[4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _2653_ (.RESET_B(net155),
    .D(_0028_),
    .Q(\u_model_loader.byte_idx_q[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2654_ (.RESET_B(net153),
    .D(net967),
    .Q(\leaf_value_flat[0] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2655_ (.RESET_B(net151),
    .D(net969),
    .Q(\leaf_value_flat[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2656_ (.RESET_B(net149),
    .D(net927),
    .Q(\leaf_value_flat[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2657_ (.RESET_B(net147),
    .D(_0032_),
    .Q(\leaf_value_flat[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2658_ (.RESET_B(net145),
    .D(net866),
    .Q(\leaf_value_flat[4] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2659_ (.RESET_B(net143),
    .D(net891),
    .Q(\leaf_value_flat[5] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2660_ (.RESET_B(net141),
    .D(net857),
    .Q(\leaf_value_flat[6] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2661_ (.RESET_B(net139),
    .D(net981),
    .Q(\leaf_value_flat[7] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2662_ (.RESET_B(net137),
    .D(net915),
    .Q(\leaf_value_flat[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2663_ (.RESET_B(net135),
    .D(net1016),
    .Q(\leaf_value_flat[9] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2664_ (.RESET_B(net133),
    .D(net853),
    .Q(\leaf_value_flat[10] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2665_ (.RESET_B(net131),
    .D(_0040_),
    .Q(\leaf_value_flat[11] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2666_ (.RESET_B(net129),
    .D(net1003),
    .Q(\leaf_value_flat[12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2667_ (.RESET_B(net127),
    .D(net1035),
    .Q(\leaf_value_flat[13] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2668_ (.RESET_B(net125),
    .D(net825),
    .Q(\leaf_value_flat[14] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2669_ (.RESET_B(net123),
    .D(net873),
    .Q(\leaf_value_flat[15] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2670_ (.RESET_B(net121),
    .D(net1010),
    .Q(\leaf_value_flat[16] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2671_ (.RESET_B(net119),
    .D(net935),
    .Q(\leaf_value_flat[17] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2672_ (.RESET_B(net117),
    .D(net861),
    .Q(\leaf_value_flat[18] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2673_ (.RESET_B(net115),
    .D(_0048_),
    .Q(\leaf_value_flat[19] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2674_ (.RESET_B(net113),
    .D(net957),
    .Q(\leaf_value_flat[20] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2675_ (.RESET_B(net111),
    .D(net902),
    .Q(\leaf_value_flat[21] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2676_ (.RESET_B(net109),
    .D(net939),
    .Q(\leaf_value_flat[22] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2677_ (.RESET_B(net107),
    .D(net1040),
    .Q(\leaf_value_flat[23] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2678_ (.RESET_B(net105),
    .D(net1025),
    .Q(\leaf_value_flat[24] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2679_ (.RESET_B(net103),
    .D(net1023),
    .Q(\leaf_value_flat[25] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2680_ (.RESET_B(net101),
    .D(net963),
    .Q(\leaf_value_flat[26] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2681_ (.RESET_B(net99),
    .D(_0056_),
    .Q(\leaf_value_flat[27] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2682_ (.RESET_B(net97),
    .D(net823),
    .Q(\leaf_value_flat[28] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2683_ (.RESET_B(net95),
    .D(net1018),
    .Q(\leaf_value_flat[29] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2684_ (.RESET_B(net93),
    .D(net959),
    .Q(\leaf_value_flat[30] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _2685_ (.RESET_B(net91),
    .D(net983),
    .Q(\leaf_value_flat[31] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2686_ (.RESET_B(net89),
    .D(net887),
    .Q(\leaf_value_flat[32] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2687_ (.RESET_B(net87),
    .D(net847),
    .Q(\leaf_value_flat[33] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2688_ (.RESET_B(net85),
    .D(net937),
    .Q(\leaf_value_flat[34] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2689_ (.RESET_B(net83),
    .D(_0064_),
    .Q(\leaf_value_flat[35] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2690_ (.RESET_B(net81),
    .D(net919),
    .Q(\leaf_value_flat[36] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2691_ (.RESET_B(net79),
    .D(net844),
    .Q(\leaf_value_flat[37] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2692_ (.RESET_B(net77),
    .D(net842),
    .Q(\leaf_value_flat[38] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2693_ (.RESET_B(net75),
    .D(net838),
    .Q(\leaf_value_flat[39] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2694_ (.RESET_B(net73),
    .D(net889),
    .Q(\leaf_value_flat[40] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2695_ (.RESET_B(net71),
    .D(net911),
    .Q(\leaf_value_flat[41] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2696_ (.RESET_B(net69),
    .D(net879),
    .Q(\leaf_value_flat[42] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2697_ (.RESET_B(net67),
    .D(_0072_),
    .Q(\leaf_value_flat[43] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2698_ (.RESET_B(net65),
    .D(net895),
    .Q(\leaf_value_flat[44] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2699_ (.RESET_B(net63),
    .D(net829),
    .Q(\leaf_value_flat[45] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2700_ (.RESET_B(net61),
    .D(net840),
    .Q(\leaf_value_flat[46] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2701_ (.RESET_B(net59),
    .D(net904),
    .Q(\leaf_value_flat[47] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2702_ (.RESET_B(net57),
    .D(net868),
    .Q(\leaf_value_flat[48] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2703_ (.RESET_B(net55),
    .D(net929),
    .Q(\leaf_value_flat[49] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2704_ (.RESET_B(net53),
    .D(net991),
    .Q(\leaf_value_flat[50] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2705_ (.RESET_B(net51),
    .D(_0080_),
    .Q(\leaf_value_flat[51] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _2706_ (.RESET_B(net49),
    .D(net985),
    .Q(\leaf_value_flat[52] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2707_ (.RESET_B(net47),
    .D(net943),
    .Q(\leaf_value_flat[53] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _2708_ (.RESET_B(net45),
    .D(net948),
    .Q(\leaf_value_flat[54] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2709_ (.RESET_B(net43),
    .D(net925),
    .Q(\leaf_value_flat[55] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2710_ (.RESET_B(net41),
    .D(net955),
    .Q(\leaf_value_flat[56] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2711_ (.RESET_B(net39),
    .D(net855),
    .Q(\leaf_value_flat[57] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _2712_ (.RESET_B(net37),
    .D(net1001),
    .Q(\leaf_value_flat[58] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _2713_ (.RESET_B(net35),
    .D(net877),
    .Q(\leaf_value_flat[59] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2714_ (.RESET_B(net33),
    .D(net831),
    .Q(\leaf_value_flat[60] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _2715_ (.RESET_B(net31),
    .D(net933),
    .Q(\leaf_value_flat[61] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2716_ (.RESET_B(net29),
    .D(net821),
    .Q(\leaf_value_flat[62] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _2717_ (.RESET_B(net27),
    .D(net931),
    .Q(\leaf_value_flat[63] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _2718_ (.RESET_B(net25),
    .D(_0093_),
    .Q(\node_right_flat[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2719_ (.RESET_B(net23),
    .D(_0094_),
    .Q(\node_right_flat[1] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2720_ (.RESET_B(net21),
    .D(_0095_),
    .Q(\node_right_flat[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2721_ (.RESET_B(net19),
    .D(net344),
    .Q(\node_right_flat[3] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2722_ (.RESET_B(net328),
    .D(_0097_),
    .Q(\node_right_flat[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2723_ (.RESET_B(net326),
    .D(_0098_),
    .Q(\node_right_flat[5] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2724_ (.RESET_B(net324),
    .D(_0099_),
    .Q(\node_right_flat[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2725_ (.RESET_B(net322),
    .D(net367),
    .Q(\node_right_flat[7] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2726_ (.RESET_B(net320),
    .D(net898),
    .Q(\node_right_flat[8] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2727_ (.RESET_B(net318),
    .D(net909),
    .Q(\node_right_flat[9] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2728_ (.RESET_B(net316),
    .D(net1006),
    .Q(\node_right_flat[10] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2729_ (.RESET_B(net314),
    .D(_0104_),
    .Q(\node_right_flat[11] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2730_ (.RESET_B(net310),
    .D(_0105_),
    .Q(\node_right_flat[12] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2731_ (.RESET_B(net308),
    .D(_0106_),
    .Q(\node_right_flat[13] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2732_ (.RESET_B(net306),
    .D(_0107_),
    .Q(\node_right_flat[14] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2733_ (.RESET_B(net304),
    .D(_0108_),
    .Q(\node_right_flat[15] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2734_ (.RESET_B(net302),
    .D(net768),
    .Q(\node_right_flat[16] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2735_ (.RESET_B(net300),
    .D(net783),
    .Q(\node_right_flat[17] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2736_ (.RESET_B(net298),
    .D(_0111_),
    .Q(\node_right_flat[18] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2737_ (.RESET_B(net296),
    .D(net353),
    .Q(\node_right_flat[19] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2738_ (.RESET_B(net294),
    .D(net766),
    .Q(\node_right_flat[20] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2739_ (.RESET_B(net292),
    .D(net827),
    .Q(\node_right_flat[21] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2740_ (.RESET_B(net290),
    .D(_0115_),
    .Q(\node_right_flat[22] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2741_ (.RESET_B(net288),
    .D(net560),
    .Q(\node_right_flat[23] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2742_ (.RESET_B(net286),
    .D(_0117_),
    .Q(\node_right_flat[24] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2743_ (.RESET_B(net284),
    .D(_0118_),
    .Q(\node_right_flat[25] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2744_ (.RESET_B(net282),
    .D(_0119_),
    .Q(\node_right_flat[26] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2745_ (.RESET_B(net280),
    .D(net342),
    .Q(\node_right_flat[27] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2746_ (.RESET_B(net278),
    .D(_0121_),
    .Q(\node_left_flat[0] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2747_ (.RESET_B(net276),
    .D(_0122_),
    .Q(\node_left_flat[1] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2748_ (.RESET_B(net274),
    .D(_0123_),
    .Q(\node_left_flat[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2749_ (.RESET_B(net272),
    .D(net369),
    .Q(\node_left_flat[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2750_ (.RESET_B(net270),
    .D(_0125_),
    .Q(\node_left_flat[4] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _2751_ (.RESET_B(net268),
    .D(_0126_),
    .Q(\node_left_flat[5] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2752_ (.RESET_B(net266),
    .D(_0127_),
    .Q(\node_left_flat[6] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2753_ (.RESET_B(net264),
    .D(net338),
    .Q(\node_left_flat[7] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2754_ (.RESET_B(net262),
    .D(net1031),
    .Q(\node_left_flat[8] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2755_ (.RESET_B(net260),
    .D(net971),
    .Q(\node_left_flat[9] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2756_ (.RESET_B(net258),
    .D(net906),
    .Q(\node_left_flat[10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2757_ (.RESET_B(net256),
    .D(_0132_),
    .Q(\node_left_flat[11] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2758_ (.RESET_B(net254),
    .D(_0133_),
    .Q(\node_left_flat[12] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _2759_ (.RESET_B(net252),
    .D(_0134_),
    .Q(\node_left_flat[13] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2760_ (.RESET_B(net250),
    .D(_0135_),
    .Q(\node_left_flat[14] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2761_ (.RESET_B(net248),
    .D(net604),
    .Q(\node_left_flat[15] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _2762_ (.RESET_B(net246),
    .D(net679),
    .Q(\node_left_flat[16] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2763_ (.RESET_B(net244),
    .D(net638),
    .Q(\node_left_flat[17] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2764_ (.RESET_B(net242),
    .D(_0139_),
    .Q(\node_left_flat[18] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2765_ (.RESET_B(net240),
    .D(net569),
    .Q(\node_left_flat[19] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2766_ (.RESET_B(net238),
    .D(_0141_),
    .Q(\node_left_flat[20] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2767_ (.RESET_B(net236),
    .D(_0142_),
    .Q(\node_left_flat[21] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2768_ (.RESET_B(net234),
    .D(_0143_),
    .Q(\node_left_flat[22] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2769_ (.RESET_B(net232),
    .D(net336),
    .Q(\node_left_flat[23] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2770_ (.RESET_B(net230),
    .D(net630),
    .Q(\node_left_flat[24] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2771_ (.RESET_B(net228),
    .D(net616),
    .Q(\node_left_flat[25] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2772_ (.RESET_B(net226),
    .D(_0147_),
    .Q(\node_left_flat[26] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2773_ (.RESET_B(net224),
    .D(net371),
    .Q(\node_left_flat[27] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2774_ (.RESET_B(net222),
    .D(_0149_),
    .Q(\node_threshold_flat[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2775_ (.RESET_B(net220),
    .D(_0150_),
    .Q(\node_threshold_flat[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2776_ (.RESET_B(net218),
    .D(_0151_),
    .Q(\node_threshold_flat[2] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2777_ (.RESET_B(net216),
    .D(_0152_),
    .Q(\node_threshold_flat[3] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2778_ (.RESET_B(net214),
    .D(net600),
    .Q(\node_threshold_flat[4] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2779_ (.RESET_B(net212),
    .D(net610),
    .Q(\node_threshold_flat[5] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2780_ (.RESET_B(net210),
    .D(net578),
    .Q(\node_threshold_flat[6] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2781_ (.RESET_B(net208),
    .D(net672),
    .Q(\node_threshold_flat[7] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2782_ (.RESET_B(net206),
    .D(_0157_),
    .Q(\node_threshold_flat[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2783_ (.RESET_B(net204),
    .D(_0158_),
    .Q(\node_threshold_flat[9] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2784_ (.RESET_B(net202),
    .D(net660),
    .Q(\node_threshold_flat[10] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2785_ (.RESET_B(net197),
    .D(net375),
    .Q(\node_threshold_flat[11] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2786_ (.RESET_B(net193),
    .D(_0161_),
    .Q(\node_threshold_flat[12] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2787_ (.RESET_B(net189),
    .D(_0162_),
    .Q(\node_threshold_flat[13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2788_ (.RESET_B(net185),
    .D(_0163_),
    .Q(\node_threshold_flat[14] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2789_ (.RESET_B(net180),
    .D(_0164_),
    .Q(\node_threshold_flat[15] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2790_ (.RESET_B(net176),
    .D(net358),
    .Q(\node_threshold_flat[16] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2791_ (.RESET_B(net172),
    .D(net373),
    .Q(\node_threshold_flat[17] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2792_ (.RESET_B(net168),
    .D(net582),
    .Q(\node_threshold_flat[18] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2793_ (.RESET_B(net162),
    .D(net602),
    .Q(\node_threshold_flat[19] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2794_ (.RESET_B(net158),
    .D(_0169_),
    .Q(\node_threshold_flat[20] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2795_ (.RESET_B(net154),
    .D(_0170_),
    .Q(\node_threshold_flat[21] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2796_ (.RESET_B(net150),
    .D(_0171_),
    .Q(\node_threshold_flat[22] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2797_ (.RESET_B(net146),
    .D(net733),
    .Q(\node_threshold_flat[23] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2798_ (.RESET_B(net142),
    .D(net941),
    .Q(\node_threshold_flat[24] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2799_ (.RESET_B(net138),
    .D(net987),
    .Q(\node_threshold_flat[25] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2800_ (.RESET_B(net134),
    .D(net1008),
    .Q(\node_threshold_flat[26] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2801_ (.RESET_B(net130),
    .D(_0176_),
    .Q(\node_threshold_flat[27] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _2802_ (.RESET_B(net126),
    .D(net1046),
    .Q(\node_threshold_flat[28] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2803_ (.RESET_B(net122),
    .D(net1044),
    .Q(\node_threshold_flat[29] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _2804_ (.RESET_B(net118),
    .D(net1033),
    .Q(\node_threshold_flat[30] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2805_ (.RESET_B(net114),
    .D(net993),
    .Q(\node_threshold_flat[31] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2806_ (.RESET_B(net110),
    .D(_0181_),
    .Q(\node_threshold_flat[32] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2807_ (.RESET_B(net106),
    .D(_0182_),
    .Q(\node_threshold_flat[33] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _2808_ (.RESET_B(net102),
    .D(_0183_),
    .Q(\node_threshold_flat[34] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2809_ (.RESET_B(net98),
    .D(_0184_),
    .Q(\node_threshold_flat[35] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2810_ (.RESET_B(net94),
    .D(net351),
    .Q(\node_threshold_flat[36] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2811_ (.RESET_B(net90),
    .D(net355),
    .Q(\node_threshold_flat[37] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2812_ (.RESET_B(net86),
    .D(net360),
    .Q(\node_threshold_flat[38] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2813_ (.RESET_B(net82),
    .D(net566),
    .Q(\node_threshold_flat[39] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2814_ (.RESET_B(net78),
    .D(_0189_),
    .Q(\node_threshold_flat[40] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2815_ (.RESET_B(net74),
    .D(_0190_),
    .Q(\node_threshold_flat[41] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2816_ (.RESET_B(net70),
    .D(_0191_),
    .Q(\node_threshold_flat[42] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _2817_ (.RESET_B(net66),
    .D(_0192_),
    .Q(\node_threshold_flat[43] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2818_ (.RESET_B(net62),
    .D(_0193_),
    .Q(\node_threshold_flat[44] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2819_ (.RESET_B(net58),
    .D(net789),
    .Q(\node_threshold_flat[45] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2820_ (.RESET_B(net54),
    .D(net702),
    .Q(\node_threshold_flat[46] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2821_ (.RESET_B(net50),
    .D(net779),
    .Q(\node_threshold_flat[47] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2822_ (.RESET_B(net46),
    .D(_0197_),
    .Q(\node_threshold_flat[48] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2823_ (.RESET_B(net42),
    .D(_0198_),
    .Q(\node_threshold_flat[49] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2824_ (.RESET_B(net38),
    .D(net607),
    .Q(\node_threshold_flat[50] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2825_ (.RESET_B(net34),
    .D(_0200_),
    .Q(\node_threshold_flat[51] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2826_ (.RESET_B(net30),
    .D(_0201_),
    .Q(\node_threshold_flat[52] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _2827_ (.RESET_B(net26),
    .D(_0202_),
    .Q(\node_threshold_flat[53] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2828_ (.RESET_B(net22),
    .D(_0203_),
    .Q(\node_threshold_flat[54] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _2829_ (.RESET_B(net329),
    .D(net641),
    .Q(\node_threshold_flat[55] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2830_ (.RESET_B(net325),
    .D(_0205_),
    .Q(\node_feature_flat[0] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2831_ (.RESET_B(net321),
    .D(_0206_),
    .Q(\node_feature_flat[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2832_ (.RESET_B(net317),
    .D(_0207_),
    .Q(\node_feature_flat[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2833_ (.RESET_B(net311),
    .D(_0208_),
    .Q(\node_feature_flat[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2834_ (.RESET_B(net307),
    .D(_0209_),
    .Q(\node_feature_flat[4] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2835_ (.RESET_B(net303),
    .D(_0210_),
    .Q(\node_feature_flat[5] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _2836_ (.RESET_B(net299),
    .D(net1027),
    .Q(\node_feature_flat[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2837_ (.RESET_B(net295),
    .D(net979),
    .Q(\node_feature_flat[7] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2838_ (.RESET_B(net291),
    .D(net961),
    .Q(\node_feature_flat[8] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _2839_ (.RESET_B(net287),
    .D(_0214_),
    .Q(\node_feature_flat[9] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2840_ (.RESET_B(net283),
    .D(_0215_),
    .Q(\node_feature_flat[10] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _2841_ (.RESET_B(net279),
    .D(_0216_),
    .Q(\node_feature_flat[11] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _2842_ (.RESET_B(net275),
    .D(_0217_),
    .Q(\node_feature_flat[12] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2843_ (.RESET_B(net271),
    .D(net684),
    .Q(\node_feature_flat[13] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _2844_ (.RESET_B(net267),
    .D(_0219_),
    .Q(\node_feature_flat[14] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2845_ (.RESET_B(net263),
    .D(net612),
    .Q(\node_feature_flat[15] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2846_ (.RESET_B(net259),
    .D(_0221_),
    .Q(\node_feature_flat[16] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2847_ (.RESET_B(net255),
    .D(_0222_),
    .Q(\node_feature_flat[17] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _2848_ (.RESET_B(net251),
    .D(_0223_),
    .Q(\node_feature_flat[18] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2849_ (.RESET_B(net247),
    .D(_0224_),
    .Q(\node_feature_flat[19] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2850_ (.RESET_B(net243),
    .D(net664),
    .Q(\node_feature_flat[20] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _2851_ (.RESET_B(net239),
    .D(net921),
    .Q(model_loaded),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _2852_ (.RESET_B(net235),
    .D(net587),
    .Q(\u_feature_loader.feature_idx_q[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2853_ (.RESET_B(net231),
    .D(_0228_),
    .Q(\u_feature_loader.feature_idx_q[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2854_ (.RESET_B(net227),
    .D(_0229_),
    .Q(\u_feature_loader.feature_idx_q[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _2855_ (.RESET_B(net223),
    .D(net644),
    .Q(\u_feature_loader.feature_idx_q[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2856_ (.RESET_B(net219),
    .D(net347),
    .Q(\feature_vector_flat[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2857_ (.RESET_B(net215),
    .D(net632),
    .Q(\feature_vector_flat[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2858_ (.RESET_B(net211),
    .D(net349),
    .Q(\feature_vector_flat[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2859_ (.RESET_B(net207),
    .D(net564),
    .Q(\feature_vector_flat[3] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2860_ (.RESET_B(net203),
    .D(net589),
    .Q(\feature_vector_flat[4] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2861_ (.RESET_B(net195),
    .D(net592),
    .Q(\feature_vector_flat[5] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2862_ (.RESET_B(net187),
    .D(net340),
    .Q(\feature_vector_flat[6] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2863_ (.RESET_B(net178),
    .D(net618),
    .Q(\feature_vector_flat[7] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2864_ (.RESET_B(net170),
    .D(_0239_),
    .Q(\feature_vector_flat[8] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2865_ (.RESET_B(net160),
    .D(_0240_),
    .Q(\feature_vector_flat[9] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2866_ (.RESET_B(net152),
    .D(_0241_),
    .Q(\feature_vector_flat[10] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2867_ (.RESET_B(net144),
    .D(_0242_),
    .Q(\feature_vector_flat[11] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2868_ (.RESET_B(net136),
    .D(_0243_),
    .Q(\feature_vector_flat[12] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2869_ (.RESET_B(net128),
    .D(_0244_),
    .Q(\feature_vector_flat[13] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2870_ (.RESET_B(net120),
    .D(net796),
    .Q(\feature_vector_flat[14] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2871_ (.RESET_B(net112),
    .D(_0246_),
    .Q(\feature_vector_flat[15] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2872_ (.RESET_B(net104),
    .D(net975),
    .Q(\feature_vector_flat[16] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2873_ (.RESET_B(net96),
    .D(net900),
    .Q(\feature_vector_flat[17] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2874_ (.RESET_B(net88),
    .D(net1012),
    .Q(\feature_vector_flat[18] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2875_ (.RESET_B(net80),
    .D(net989),
    .Q(\feature_vector_flat[19] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2876_ (.RESET_B(net72),
    .D(net953),
    .Q(\feature_vector_flat[20] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2877_ (.RESET_B(net64),
    .D(net913),
    .Q(\feature_vector_flat[21] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2878_ (.RESET_B(net56),
    .D(net995),
    .Q(\feature_vector_flat[22] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2879_ (.RESET_B(net48),
    .D(net951),
    .Q(\feature_vector_flat[23] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2880_ (.RESET_B(net40),
    .D(_0255_),
    .Q(\feature_vector_flat[24] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2881_ (.RESET_B(net32),
    .D(_0256_),
    .Q(\feature_vector_flat[25] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _2882_ (.RESET_B(net24),
    .D(_0257_),
    .Q(\feature_vector_flat[26] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2883_ (.RESET_B(net327),
    .D(_0258_),
    .Q(\feature_vector_flat[27] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2884_ (.RESET_B(net319),
    .D(net745),
    .Q(\feature_vector_flat[28] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _2885_ (.RESET_B(net309),
    .D(_0260_),
    .Q(\feature_vector_flat[29] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2886_ (.RESET_B(net301),
    .D(net736),
    .Q(\feature_vector_flat[30] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2887_ (.RESET_B(net293),
    .D(_0262_),
    .Q(\feature_vector_flat[31] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2888_ (.RESET_B(net285),
    .D(net572),
    .Q(\feature_vector_flat[32] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2889_ (.RESET_B(net277),
    .D(net365),
    .Q(\feature_vector_flat[33] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2890_ (.RESET_B(net269),
    .D(net580),
    .Q(\feature_vector_flat[34] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2891_ (.RESET_B(net261),
    .D(net574),
    .Q(\feature_vector_flat[35] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2892_ (.RESET_B(net253),
    .D(net576),
    .Q(\feature_vector_flat[36] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2893_ (.RESET_B(net245),
    .D(net362),
    .Q(\feature_vector_flat[37] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2894_ (.RESET_B(net237),
    .D(net584),
    .Q(\feature_vector_flat[38] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2895_ (.RESET_B(net229),
    .D(net558),
    .Q(\feature_vector_flat[39] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2896_ (.RESET_B(net221),
    .D(net654),
    .Q(\feature_vector_flat[40] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2897_ (.RESET_B(net213),
    .D(_0272_),
    .Q(\feature_vector_flat[41] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2898_ (.RESET_B(net205),
    .D(_0273_),
    .Q(\feature_vector_flat[42] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2899_ (.RESET_B(net191),
    .D(_0274_),
    .Q(\feature_vector_flat[43] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2900_ (.RESET_B(net174),
    .D(_0275_),
    .Q(\feature_vector_flat[44] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2901_ (.RESET_B(net156),
    .D(net658),
    .Q(\feature_vector_flat[45] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2902_ (.RESET_B(net140),
    .D(net621),
    .Q(\feature_vector_flat[46] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2903_ (.RESET_B(net124),
    .D(_0278_),
    .Q(\feature_vector_flat[47] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _2904_ (.RESET_B(net108),
    .D(net1014),
    .Q(\feature_vector_flat[48] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2905_ (.RESET_B(net92),
    .D(net850),
    .Q(\feature_vector_flat[49] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _2906_ (.RESET_B(net76),
    .D(net965),
    .Q(\feature_vector_flat[50] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2907_ (.RESET_B(net60),
    .D(net923),
    .Q(\feature_vector_flat[51] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2908_ (.RESET_B(net44),
    .D(net999),
    .Q(\feature_vector_flat[52] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _2909_ (.RESET_B(net28),
    .D(net859),
    .Q(\feature_vector_flat[53] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _2910_ (.RESET_B(net323),
    .D(net1029),
    .Q(\feature_vector_flat[54] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _2911_ (.RESET_B(net305),
    .D(net817),
    .Q(\feature_vector_flat[55] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2912_ (.RESET_B(net289),
    .D(net864),
    .Q(\feature_vector_flat[56] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2913_ (.RESET_B(net273),
    .D(_0288_),
    .Q(\feature_vector_flat[57] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _2914_ (.RESET_B(net257),
    .D(net773),
    .Q(\feature_vector_flat[58] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2915_ (.RESET_B(net241),
    .D(_0290_),
    .Q(\feature_vector_flat[59] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2916_ (.RESET_B(net225),
    .D(net720),
    .Q(\feature_vector_flat[60] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2917_ (.RESET_B(net209),
    .D(_0292_),
    .Q(\feature_vector_flat[61] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _2918_ (.RESET_B(net182),
    .D(net717),
    .Q(\feature_vector_flat[62] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _2919_ (.RESET_B(net313),
    .D(_0294_),
    .Q(\feature_vector_flat[63] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _2920_ (.RESET_B(net132),
    .D(net1055),
    .Q(\u_tree_core.state_q[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2921_ (.RESET_B(net148),
    .D(net1062),
    .Q(\u_tree_core.state_q[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2922_ (.RESET_B(net116),
    .D(_0295_),
    .Q(clear_cmd),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _2923_ (.RESET_B(net100),
    .D(net690),
    .Q(core_busy),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _2924_ (.RESET_B(net68),
    .D(_0297_),
    .Q(uo_out[0]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2925_ (.RESET_B(net36),
    .D(net730),
    .Q(uo_out[1]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _2926_ (.RESET_B(net315),
    .D(net749),
    .Q(uo_out[2]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2927_ (.RESET_B(net281),
    .D(net819),
    .Q(uo_out[3]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2928_ (.RESET_B(net249),
    .D(net699),
    .Q(uo_out[4]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2929_ (.RESET_B(net217),
    .D(net724),
    .Q(uo_out[5]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _2930_ (.RESET_B(net164),
    .D(net762),
    .Q(uo_out[6]),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _2931_ (.RESET_B(net84),
    .D(net692),
    .Q(uo_out[7]),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _2932_ (.RESET_B(net20),
    .D(net739),
    .Q(core_error),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _2933_ (.RESET_B(net265),
    .D(net1042),
    .Q(\u_tree_core.depth_q[0] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _2934_ (.RESET_B(net199),
    .D(net595),
    .Q(\u_tree_core.depth_q[1] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _2935_ (.RESET_B(net52),
    .D(net1079),
    .Q(\u_tree_core.current_node_q[0] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _2936_ (.RESET_B(net233),
    .D(net1077),
    .Q(\u_tree_core.current_node_q[1] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _2937_ (.RESET_B(net297),
    .D(net1068),
    .Q(\u_tree_core.current_node_q[2] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_tiehi _2932__20 (.L_HI(net20));
 sg13g2_tiehi _2720__21 (.L_HI(net21));
 sg13g2_tiehi _2828__22 (.L_HI(net22));
 sg13g2_tiehi _2719__23 (.L_HI(net23));
 sg13g2_tiehi _2882__24 (.L_HI(net24));
 sg13g2_tiehi _2718__25 (.L_HI(net25));
 sg13g2_tiehi _2827__26 (.L_HI(net26));
 sg13g2_tiehi _2717__27 (.L_HI(net27));
 sg13g2_tiehi _2909__28 (.L_HI(net28));
 sg13g2_tiehi _2716__29 (.L_HI(net29));
 sg13g2_tiehi _2826__30 (.L_HI(net30));
 sg13g2_tiehi _2715__31 (.L_HI(net31));
 sg13g2_tiehi _2881__32 (.L_HI(net32));
 sg13g2_tiehi _2714__33 (.L_HI(net33));
 sg13g2_tiehi _2825__34 (.L_HI(net34));
 sg13g2_tiehi _2713__35 (.L_HI(net35));
 sg13g2_tiehi _2925__36 (.L_HI(net36));
 sg13g2_tiehi _2712__37 (.L_HI(net37));
 sg13g2_tiehi _2824__38 (.L_HI(net38));
 sg13g2_tiehi _2711__39 (.L_HI(net39));
 sg13g2_tiehi _2880__40 (.L_HI(net40));
 sg13g2_tiehi _2710__41 (.L_HI(net41));
 sg13g2_tiehi _2823__42 (.L_HI(net42));
 sg13g2_tiehi _2709__43 (.L_HI(net43));
 sg13g2_tiehi _2908__44 (.L_HI(net44));
 sg13g2_tiehi _2708__45 (.L_HI(net45));
 sg13g2_tiehi _2822__46 (.L_HI(net46));
 sg13g2_tiehi _2707__47 (.L_HI(net47));
 sg13g2_tiehi _2879__48 (.L_HI(net48));
 sg13g2_tiehi _2706__49 (.L_HI(net49));
 sg13g2_tiehi _2821__50 (.L_HI(net50));
 sg13g2_tiehi _2705__51 (.L_HI(net51));
 sg13g2_tiehi _2935__52 (.L_HI(net52));
 sg13g2_tiehi _2704__53 (.L_HI(net53));
 sg13g2_tiehi _2820__54 (.L_HI(net54));
 sg13g2_tiehi _2703__55 (.L_HI(net55));
 sg13g2_tiehi _2878__56 (.L_HI(net56));
 sg13g2_tiehi _2702__57 (.L_HI(net57));
 sg13g2_tiehi _2819__58 (.L_HI(net58));
 sg13g2_tiehi _2701__59 (.L_HI(net59));
 sg13g2_tiehi _2907__60 (.L_HI(net60));
 sg13g2_tiehi _2700__61 (.L_HI(net61));
 sg13g2_tiehi _2818__62 (.L_HI(net62));
 sg13g2_tiehi _2699__63 (.L_HI(net63));
 sg13g2_tiehi _2877__64 (.L_HI(net64));
 sg13g2_tiehi _2698__65 (.L_HI(net65));
 sg13g2_tiehi _2817__66 (.L_HI(net66));
 sg13g2_tiehi _2697__67 (.L_HI(net67));
 sg13g2_tiehi _2924__68 (.L_HI(net68));
 sg13g2_tiehi _2696__69 (.L_HI(net69));
 sg13g2_tiehi _2816__70 (.L_HI(net70));
 sg13g2_tiehi _2695__71 (.L_HI(net71));
 sg13g2_tiehi _2876__72 (.L_HI(net72));
 sg13g2_tiehi _2694__73 (.L_HI(net73));
 sg13g2_tiehi _2815__74 (.L_HI(net74));
 sg13g2_tiehi _2693__75 (.L_HI(net75));
 sg13g2_tiehi _2906__76 (.L_HI(net76));
 sg13g2_tiehi _2692__77 (.L_HI(net77));
 sg13g2_tiehi _2814__78 (.L_HI(net78));
 sg13g2_tiehi _2691__79 (.L_HI(net79));
 sg13g2_tiehi _2875__80 (.L_HI(net80));
 sg13g2_tiehi _2690__81 (.L_HI(net81));
 sg13g2_tiehi _2813__82 (.L_HI(net82));
 sg13g2_tiehi _2689__83 (.L_HI(net83));
 sg13g2_tiehi _2931__84 (.L_HI(net84));
 sg13g2_tiehi _2688__85 (.L_HI(net85));
 sg13g2_tiehi _2812__86 (.L_HI(net86));
 sg13g2_tiehi _2687__87 (.L_HI(net87));
 sg13g2_tiehi _2874__88 (.L_HI(net88));
 sg13g2_tiehi _2686__89 (.L_HI(net89));
 sg13g2_tiehi _2811__90 (.L_HI(net90));
 sg13g2_tiehi _2685__91 (.L_HI(net91));
 sg13g2_tiehi _2905__92 (.L_HI(net92));
 sg13g2_tiehi _2684__93 (.L_HI(net93));
 sg13g2_tiehi _2810__94 (.L_HI(net94));
 sg13g2_tiehi _2683__95 (.L_HI(net95));
 sg13g2_tiehi _2873__96 (.L_HI(net96));
 sg13g2_tiehi _2682__97 (.L_HI(net97));
 sg13g2_tiehi _2809__98 (.L_HI(net98));
 sg13g2_tiehi _2681__99 (.L_HI(net99));
 sg13g2_tiehi _2923__100 (.L_HI(net100));
 sg13g2_tiehi _2680__101 (.L_HI(net101));
 sg13g2_tiehi _2808__102 (.L_HI(net102));
 sg13g2_tiehi _2679__103 (.L_HI(net103));
 sg13g2_tiehi _2872__104 (.L_HI(net104));
 sg13g2_tiehi _2678__105 (.L_HI(net105));
 sg13g2_tiehi _2807__106 (.L_HI(net106));
 sg13g2_tiehi _2677__107 (.L_HI(net107));
 sg13g2_tiehi _2904__108 (.L_HI(net108));
 sg13g2_tiehi _2676__109 (.L_HI(net109));
 sg13g2_tiehi _2806__110 (.L_HI(net110));
 sg13g2_tiehi _2675__111 (.L_HI(net111));
 sg13g2_tiehi _2871__112 (.L_HI(net112));
 sg13g2_tiehi _2674__113 (.L_HI(net113));
 sg13g2_tiehi _2805__114 (.L_HI(net114));
 sg13g2_tiehi _2673__115 (.L_HI(net115));
 sg13g2_tiehi _2922__116 (.L_HI(net116));
 sg13g2_tiehi _2672__117 (.L_HI(net117));
 sg13g2_tiehi _2804__118 (.L_HI(net118));
 sg13g2_tiehi _2671__119 (.L_HI(net119));
 sg13g2_tiehi _2870__120 (.L_HI(net120));
 sg13g2_tiehi _2670__121 (.L_HI(net121));
 sg13g2_tiehi _2803__122 (.L_HI(net122));
 sg13g2_tiehi _2669__123 (.L_HI(net123));
 sg13g2_tiehi _2903__124 (.L_HI(net124));
 sg13g2_tiehi _2668__125 (.L_HI(net125));
 sg13g2_tiehi _2802__126 (.L_HI(net126));
 sg13g2_tiehi _2667__127 (.L_HI(net127));
 sg13g2_tiehi _2869__128 (.L_HI(net128));
 sg13g2_tiehi _2666__129 (.L_HI(net129));
 sg13g2_tiehi _2801__130 (.L_HI(net130));
 sg13g2_tiehi _2665__131 (.L_HI(net131));
 sg13g2_tiehi _2920__132 (.L_HI(net132));
 sg13g2_tiehi _2664__133 (.L_HI(net133));
 sg13g2_tiehi _2800__134 (.L_HI(net134));
 sg13g2_tiehi _2663__135 (.L_HI(net135));
 sg13g2_tiehi _2868__136 (.L_HI(net136));
 sg13g2_tiehi _2662__137 (.L_HI(net137));
 sg13g2_tiehi _2799__138 (.L_HI(net138));
 sg13g2_tiehi _2661__139 (.L_HI(net139));
 sg13g2_tiehi _2902__140 (.L_HI(net140));
 sg13g2_tiehi _2660__141 (.L_HI(net141));
 sg13g2_tiehi _2798__142 (.L_HI(net142));
 sg13g2_tiehi _2659__143 (.L_HI(net143));
 sg13g2_tiehi _2867__144 (.L_HI(net144));
 sg13g2_tiehi _2658__145 (.L_HI(net145));
 sg13g2_tiehi _2797__146 (.L_HI(net146));
 sg13g2_tiehi _2657__147 (.L_HI(net147));
 sg13g2_tiehi _2921__148 (.L_HI(net148));
 sg13g2_tiehi _2656__149 (.L_HI(net149));
 sg13g2_tiehi _2796__150 (.L_HI(net150));
 sg13g2_tiehi _2655__151 (.L_HI(net151));
 sg13g2_tiehi _2866__152 (.L_HI(net152));
 sg13g2_tiehi _2654__153 (.L_HI(net153));
 sg13g2_tiehi _2795__154 (.L_HI(net154));
 sg13g2_tiehi _2653__155 (.L_HI(net155));
 sg13g2_tiehi _2901__156 (.L_HI(net156));
 sg13g2_tiehi _2652__157 (.L_HI(net157));
 sg13g2_tiehi _2794__158 (.L_HI(net158));
 sg13g2_tiehi _2651__159 (.L_HI(net159));
 sg13g2_tiehi _2865__160 (.L_HI(net160));
 sg13g2_tiehi _2650__161 (.L_HI(net161));
 sg13g2_tiehi _2793__162 (.L_HI(net162));
 sg13g2_tiehi _2649__163 (.L_HI(net163));
 sg13g2_tiehi _2930__164 (.L_HI(net164));
 sg13g2_tiehi _2648__165 (.L_HI(net165));
 sg13g2_tiehi _2647__166 (.L_HI(net166));
 sg13g2_tiehi _2646__167 (.L_HI(net167));
 sg13g2_tiehi _2792__168 (.L_HI(net168));
 sg13g2_tiehi _2645__169 (.L_HI(net169));
 sg13g2_tiehi _2864__170 (.L_HI(net170));
 sg13g2_tiehi _2644__171 (.L_HI(net171));
 sg13g2_tiehi _2791__172 (.L_HI(net172));
 sg13g2_tiehi _2643__173 (.L_HI(net173));
 sg13g2_tiehi _2900__174 (.L_HI(net174));
 sg13g2_tiehi _2642__175 (.L_HI(net175));
 sg13g2_tiehi _2790__176 (.L_HI(net176));
 sg13g2_tiehi _2641__177 (.L_HI(net177));
 sg13g2_tiehi _2863__178 (.L_HI(net178));
 sg13g2_tiehi _2640__179 (.L_HI(net179));
 sg13g2_tiehi _2789__180 (.L_HI(net180));
 sg13g2_tiehi _2639__181 (.L_HI(net181));
 sg13g2_tiehi _2918__182 (.L_HI(net182));
 sg13g2_tiehi _2638__183 (.L_HI(net183));
 sg13g2_tiehi _2637__184 (.L_HI(net184));
 sg13g2_tiehi _2788__185 (.L_HI(net185));
 sg13g2_tiehi _2636__186 (.L_HI(net186));
 sg13g2_tiehi _2862__187 (.L_HI(net187));
 sg13g2_tiehi _2635__188 (.L_HI(net188));
 sg13g2_tiehi _2787__189 (.L_HI(net189));
 sg13g2_tiehi _2634__190 (.L_HI(net190));
 sg13g2_tiehi _2899__191 (.L_HI(net191));
 sg13g2_tiehi _2633__192 (.L_HI(net192));
 sg13g2_tiehi _2786__193 (.L_HI(net193));
 sg13g2_tiehi _2632__194 (.L_HI(net194));
 sg13g2_tiehi _2861__195 (.L_HI(net195));
 sg13g2_tiehi _2631__196 (.L_HI(net196));
 sg13g2_tiehi _2785__197 (.L_HI(net197));
 sg13g2_tiehi _2630__198 (.L_HI(net198));
 sg13g2_tiehi _2934__199 (.L_HI(net199));
 sg13g2_tiehi _2629__200 (.L_HI(net200));
 sg13g2_tiehi _2628__201 (.L_HI(net201));
 sg13g2_tiehi _2784__202 (.L_HI(net202));
 sg13g2_tiehi _2860__203 (.L_HI(net203));
 sg13g2_tiehi _2783__204 (.L_HI(net204));
 sg13g2_tiehi _2898__205 (.L_HI(net205));
 sg13g2_tiehi _2782__206 (.L_HI(net206));
 sg13g2_tiehi _2859__207 (.L_HI(net207));
 sg13g2_tiehi _2781__208 (.L_HI(net208));
 sg13g2_tiehi _2917__209 (.L_HI(net209));
 sg13g2_tiehi _2780__210 (.L_HI(net210));
 sg13g2_tiehi _2858__211 (.L_HI(net211));
 sg13g2_tiehi _2779__212 (.L_HI(net212));
 sg13g2_tiehi _2897__213 (.L_HI(net213));
 sg13g2_tiehi _2778__214 (.L_HI(net214));
 sg13g2_tiehi _2857__215 (.L_HI(net215));
 sg13g2_tiehi _2777__216 (.L_HI(net216));
 sg13g2_tiehi _2929__217 (.L_HI(net217));
 sg13g2_tiehi _2776__218 (.L_HI(net218));
 sg13g2_tiehi _2856__219 (.L_HI(net219));
 sg13g2_tiehi _2775__220 (.L_HI(net220));
 sg13g2_tiehi _2896__221 (.L_HI(net221));
 sg13g2_tiehi _2774__222 (.L_HI(net222));
 sg13g2_tiehi _2855__223 (.L_HI(net223));
 sg13g2_tiehi _2773__224 (.L_HI(net224));
 sg13g2_tiehi _2916__225 (.L_HI(net225));
 sg13g2_tiehi _2772__226 (.L_HI(net226));
 sg13g2_tiehi _2854__227 (.L_HI(net227));
 sg13g2_tiehi _2771__228 (.L_HI(net228));
 sg13g2_tiehi _2895__229 (.L_HI(net229));
 sg13g2_tiehi _2770__230 (.L_HI(net230));
 sg13g2_tiehi _2853__231 (.L_HI(net231));
 sg13g2_tiehi _2769__232 (.L_HI(net232));
 sg13g2_tiehi _2936__233 (.L_HI(net233));
 sg13g2_tiehi _2768__234 (.L_HI(net234));
 sg13g2_tiehi _2852__235 (.L_HI(net235));
 sg13g2_tiehi _2767__236 (.L_HI(net236));
 sg13g2_tiehi _2894__237 (.L_HI(net237));
 sg13g2_tiehi _2766__238 (.L_HI(net238));
 sg13g2_tiehi _2851__239 (.L_HI(net239));
 sg13g2_tiehi _2765__240 (.L_HI(net240));
 sg13g2_tiehi _2915__241 (.L_HI(net241));
 sg13g2_tiehi _2764__242 (.L_HI(net242));
 sg13g2_tiehi _2850__243 (.L_HI(net243));
 sg13g2_tiehi _2763__244 (.L_HI(net244));
 sg13g2_tiehi _2893__245 (.L_HI(net245));
 sg13g2_tiehi _2762__246 (.L_HI(net246));
 sg13g2_tiehi _2849__247 (.L_HI(net247));
 sg13g2_tiehi _2761__248 (.L_HI(net248));
 sg13g2_tiehi _2928__249 (.L_HI(net249));
 sg13g2_tiehi _2760__250 (.L_HI(net250));
 sg13g2_tiehi _2848__251 (.L_HI(net251));
 sg13g2_tiehi _2759__252 (.L_HI(net252));
 sg13g2_tiehi _2892__253 (.L_HI(net253));
 sg13g2_tiehi _2758__254 (.L_HI(net254));
 sg13g2_tiehi _2847__255 (.L_HI(net255));
 sg13g2_tiehi _2757__256 (.L_HI(net256));
 sg13g2_tiehi _2914__257 (.L_HI(net257));
 sg13g2_tiehi _2756__258 (.L_HI(net258));
 sg13g2_tiehi _2846__259 (.L_HI(net259));
 sg13g2_tiehi _2755__260 (.L_HI(net260));
 sg13g2_tiehi _2891__261 (.L_HI(net261));
 sg13g2_tiehi _2754__262 (.L_HI(net262));
 sg13g2_tiehi _2845__263 (.L_HI(net263));
 sg13g2_tiehi _2753__264 (.L_HI(net264));
 sg13g2_tiehi _2933__265 (.L_HI(net265));
 sg13g2_tiehi _2752__266 (.L_HI(net266));
 sg13g2_tiehi _2844__267 (.L_HI(net267));
 sg13g2_tiehi _2751__268 (.L_HI(net268));
 sg13g2_tiehi _2890__269 (.L_HI(net269));
 sg13g2_tiehi _2750__270 (.L_HI(net270));
 sg13g2_tiehi _2843__271 (.L_HI(net271));
 sg13g2_tiehi _2749__272 (.L_HI(net272));
 sg13g2_tiehi _2913__273 (.L_HI(net273));
 sg13g2_tiehi _2748__274 (.L_HI(net274));
 sg13g2_tiehi _2842__275 (.L_HI(net275));
 sg13g2_tiehi _2747__276 (.L_HI(net276));
 sg13g2_tiehi _2889__277 (.L_HI(net277));
 sg13g2_tiehi _2746__278 (.L_HI(net278));
 sg13g2_tiehi _2841__279 (.L_HI(net279));
 sg13g2_tiehi _2745__280 (.L_HI(net280));
 sg13g2_tiehi _2927__281 (.L_HI(net281));
 sg13g2_tiehi _2744__282 (.L_HI(net282));
 sg13g2_tiehi _2840__283 (.L_HI(net283));
 sg13g2_tiehi _2743__284 (.L_HI(net284));
 sg13g2_tiehi _2888__285 (.L_HI(net285));
 sg13g2_tiehi _2742__286 (.L_HI(net286));
 sg13g2_tiehi _2839__287 (.L_HI(net287));
 sg13g2_tiehi _2741__288 (.L_HI(net288));
 sg13g2_tiehi _2912__289 (.L_HI(net289));
 sg13g2_tiehi _2740__290 (.L_HI(net290));
 sg13g2_tiehi _2838__291 (.L_HI(net291));
 sg13g2_tiehi _2739__292 (.L_HI(net292));
 sg13g2_tiehi _2887__293 (.L_HI(net293));
 sg13g2_tiehi _2738__294 (.L_HI(net294));
 sg13g2_tiehi _2837__295 (.L_HI(net295));
 sg13g2_tiehi _2737__296 (.L_HI(net296));
 sg13g2_tiehi _2937__297 (.L_HI(net297));
 sg13g2_tiehi _2736__298 (.L_HI(net298));
 sg13g2_tiehi _2836__299 (.L_HI(net299));
 sg13g2_tiehi _2735__300 (.L_HI(net300));
 sg13g2_tiehi _2886__301 (.L_HI(net301));
 sg13g2_tiehi _2734__302 (.L_HI(net302));
 sg13g2_tiehi _2835__303 (.L_HI(net303));
 sg13g2_tiehi _2733__304 (.L_HI(net304));
 sg13g2_tiehi _2911__305 (.L_HI(net305));
 sg13g2_tiehi _2732__306 (.L_HI(net306));
 sg13g2_tiehi _2834__307 (.L_HI(net307));
 sg13g2_tiehi _2731__308 (.L_HI(net308));
 sg13g2_tiehi _2885__309 (.L_HI(net309));
 sg13g2_tiehi _2730__310 (.L_HI(net310));
 sg13g2_tiehi _2833__311 (.L_HI(net311));
 sg13g2_tiehi _2627__312 (.L_HI(net312));
 sg13g2_tiehi _2919__313 (.L_HI(net313));
 sg13g2_tiehi _2729__314 (.L_HI(net314));
 sg13g2_tiehi _2926__315 (.L_HI(net315));
 sg13g2_tiehi _2728__316 (.L_HI(net316));
 sg13g2_tiehi _2832__317 (.L_HI(net317));
 sg13g2_tiehi _2727__318 (.L_HI(net318));
 sg13g2_tiehi _2884__319 (.L_HI(net319));
 sg13g2_tiehi _2726__320 (.L_HI(net320));
 sg13g2_tiehi _2831__321 (.L_HI(net321));
 sg13g2_tiehi _2725__322 (.L_HI(net322));
 sg13g2_tiehi _2910__323 (.L_HI(net323));
 sg13g2_tiehi _2724__324 (.L_HI(net324));
 sg13g2_tiehi _2830__325 (.L_HI(net325));
 sg13g2_tiehi _2723__326 (.L_HI(net326));
 sg13g2_tiehi _2883__327 (.L_HI(net327));
 sg13g2_tiehi _2722__328 (.L_HI(net328));
 sg13g2_tiehi _2829__329 (.L_HI(net329));
 sg13g2_tiehi tt_um_pgfarley_tophat_top_330 (.L_HI(net330));
 sg13g2_tiehi tt_um_pgfarley_tophat_top_331 (.L_HI(net331));
 sg13g2_tiehi tt_um_pgfarley_tophat_top_332 (.L_HI(net332));
 sg13g2_tiehi tt_um_pgfarley_tophat_top_333 (.L_HI(net333));
 sg13g2_tiehi tt_um_pgfarley_tophat_top_334 (.L_HI(net334));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tielo tt_um_pgfarley_tophat_top_14 (.L_LO(net14));
 sg13g2_tielo tt_um_pgfarley_tophat_top_15 (.L_LO(net15));
 sg13g2_tielo tt_um_pgfarley_tophat_top_16 (.L_LO(net16));
 sg13g2_tielo tt_um_pgfarley_tophat_top_17 (.L_LO(net17));
 sg13g2_tielo tt_um_pgfarley_tophat_top_18 (.L_LO(net18));
 sg13g2_tiehi _2721__19 (.L_HI(net19));
 sg13g2_buf_1 _3260_ (.A(io_ready),
    .X(uio_out[3]));
 sg13g2_buf_1 _3261_ (.A(core_busy),
    .X(uio_out[4]));
 sg13g2_buf_1 _3262_ (.A(pred_valid),
    .X(uio_out[5]));
 sg13g2_buf_1 _3263_ (.A(model_loaded),
    .X(uio_out[6]));
 sg13g2_buf_8 fanout376 (.A(_1154_),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(_1153_),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(net379),
    .X(net378));
 sg13g2_buf_8 fanout379 (.A(_1101_),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(net382),
    .X(net380));
 sg13g2_buf_8 fanout381 (.A(net382),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(_1111_),
    .X(net382));
 sg13g2_buf_8 fanout383 (.A(net386),
    .X(net383));
 sg13g2_buf_8 fanout384 (.A(net386),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(net386),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(_1064_),
    .X(net386));
 sg13g2_buf_8 fanout387 (.A(net388),
    .X(net387));
 sg13g2_buf_8 fanout388 (.A(_0390_),
    .X(net388));
 sg13g2_buf_8 fanout389 (.A(_0381_),
    .X(net389));
 sg13g2_buf_8 fanout390 (.A(_0381_),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(_0372_),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(_0372_),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(_0363_),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(_0363_),
    .X(net394));
 sg13g2_buf_8 fanout395 (.A(_0354_),
    .X(net395));
 sg13g2_buf_8 fanout396 (.A(_0354_),
    .X(net396));
 sg13g2_buf_8 fanout397 (.A(_0344_),
    .X(net397));
 sg13g2_buf_8 fanout398 (.A(_0344_),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(_0334_),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(_0334_),
    .X(net400));
 sg13g2_buf_8 fanout401 (.A(net403),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(_0325_),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(_0325_),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(_0576_),
    .X(net404));
 sg13g2_buf_8 fanout405 (.A(_0528_),
    .X(net405));
 sg13g2_buf_8 fanout406 (.A(_1147_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_0938_),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(_0938_),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(net411),
    .X(net409));
 sg13g2_buf_8 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_8 fanout411 (.A(_0716_),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(_0646_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_0646_),
    .X(net413));
 sg13g2_buf_8 fanout414 (.A(net415),
    .X(net414));
 sg13g2_buf_8 fanout415 (.A(_0646_),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(net417),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(_0597_),
    .X(net417));
 sg13g2_buf_8 fanout418 (.A(_0586_),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_8 fanout420 (.A(_0567_),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(net422),
    .X(net421));
 sg13g2_buf_8 fanout422 (.A(_0558_),
    .X(net422));
 sg13g2_buf_8 fanout423 (.A(net424),
    .X(net423));
 sg13g2_buf_1 fanout424 (.A(net425),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_0519_),
    .X(net425));
 sg13g2_buf_8 fanout426 (.A(_0518_),
    .X(net426));
 sg13g2_buf_1 fanout427 (.A(_0518_),
    .X(net427));
 sg13g2_buf_8 fanout428 (.A(net430),
    .X(net428));
 sg13g2_buf_1 fanout429 (.A(net430),
    .X(net429));
 sg13g2_buf_8 fanout430 (.A(_0478_),
    .X(net430));
 sg13g2_buf_8 fanout431 (.A(net434),
    .X(net431));
 sg13g2_buf_8 fanout432 (.A(net434),
    .X(net432));
 sg13g2_buf_8 fanout433 (.A(net434),
    .X(net433));
 sg13g2_buf_8 fanout434 (.A(_0407_),
    .X(net434));
 sg13g2_buf_8 fanout435 (.A(_1151_),
    .X(net435));
 sg13g2_buf_8 fanout436 (.A(_1151_),
    .X(net436));
 sg13g2_buf_8 fanout437 (.A(net438),
    .X(net437));
 sg13g2_buf_8 fanout438 (.A(_1135_),
    .X(net438));
 sg13g2_buf_8 fanout439 (.A(net440),
    .X(net439));
 sg13g2_buf_8 fanout440 (.A(_1126_),
    .X(net440));
 sg13g2_buf_8 fanout441 (.A(net443),
    .X(net441));
 sg13g2_buf_8 fanout442 (.A(net443),
    .X(net442));
 sg13g2_buf_8 fanout443 (.A(_0930_),
    .X(net443));
 sg13g2_buf_8 fanout444 (.A(net448),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(net448),
    .X(net445));
 sg13g2_buf_8 fanout446 (.A(net447),
    .X(net446));
 sg13g2_buf_8 fanout447 (.A(net448),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(_0921_),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(_0595_),
    .X(net449));
 sg13g2_buf_1 fanout450 (.A(_0595_),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(_0517_),
    .X(net451));
 sg13g2_buf_1 fanout452 (.A(_0517_),
    .X(net452));
 sg13g2_buf_8 fanout453 (.A(_0476_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_0476_),
    .X(net454));
 sg13g2_buf_8 fanout455 (.A(_0446_),
    .X(net455));
 sg13g2_buf_8 fanout456 (.A(_0427_),
    .X(net456));
 sg13g2_buf_8 fanout457 (.A(net458),
    .X(net457));
 sg13g2_buf_8 fanout458 (.A(_0320_),
    .X(net458));
 sg13g2_buf_8 fanout459 (.A(_1150_),
    .X(net459));
 sg13g2_buf_8 fanout460 (.A(_1150_),
    .X(net460));
 sg13g2_buf_8 fanout461 (.A(_0641_),
    .X(net461));
 sg13g2_buf_8 fanout462 (.A(_1144_),
    .X(net462));
 sg13g2_buf_8 fanout463 (.A(net464),
    .X(net463));
 sg13g2_buf_8 fanout464 (.A(_0910_),
    .X(net464));
 sg13g2_buf_8 fanout465 (.A(net468),
    .X(net465));
 sg13g2_buf_1 fanout466 (.A(net468),
    .X(net466));
 sg13g2_buf_8 fanout467 (.A(net468),
    .X(net467));
 sg13g2_buf_8 fanout468 (.A(_0908_),
    .X(net468));
 sg13g2_buf_8 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_8 fanout470 (.A(net476),
    .X(net470));
 sg13g2_buf_8 fanout471 (.A(net472),
    .X(net471));
 sg13g2_buf_8 fanout472 (.A(net476),
    .X(net472));
 sg13g2_buf_8 fanout473 (.A(net475),
    .X(net473));
 sg13g2_buf_8 fanout474 (.A(net475),
    .X(net474));
 sg13g2_buf_8 fanout475 (.A(net476),
    .X(net475));
 sg13g2_buf_8 fanout476 (.A(net482),
    .X(net476));
 sg13g2_buf_8 fanout477 (.A(net478),
    .X(net477));
 sg13g2_buf_8 fanout478 (.A(net482),
    .X(net478));
 sg13g2_buf_8 fanout479 (.A(net481),
    .X(net479));
 sg13g2_buf_8 fanout480 (.A(net481),
    .X(net480));
 sg13g2_buf_8 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_8 fanout482 (.A(_0905_),
    .X(net482));
 sg13g2_buf_8 fanout483 (.A(net484),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(net492),
    .X(net484));
 sg13g2_buf_8 fanout485 (.A(net492),
    .X(net485));
 sg13g2_buf_8 fanout486 (.A(net492),
    .X(net486));
 sg13g2_buf_8 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_8 fanout488 (.A(net492),
    .X(net488));
 sg13g2_buf_8 fanout489 (.A(net491),
    .X(net489));
 sg13g2_buf_1 fanout490 (.A(net491),
    .X(net490));
 sg13g2_buf_8 fanout491 (.A(net492),
    .X(net491));
 sg13g2_buf_8 fanout492 (.A(_0905_),
    .X(net492));
 sg13g2_buf_8 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_8 fanout494 (.A(net496),
    .X(net494));
 sg13g2_buf_8 fanout495 (.A(net516),
    .X(net495));
 sg13g2_buf_1 fanout496 (.A(net516),
    .X(net496));
 sg13g2_buf_8 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_8 fanout498 (.A(net499),
    .X(net498));
 sg13g2_buf_8 fanout499 (.A(net516),
    .X(net499));
 sg13g2_buf_8 fanout500 (.A(net501),
    .X(net500));
 sg13g2_buf_8 fanout501 (.A(net504),
    .X(net501));
 sg13g2_buf_8 fanout502 (.A(net503),
    .X(net502));
 sg13g2_buf_8 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_8 fanout504 (.A(net515),
    .X(net504));
 sg13g2_buf_8 fanout505 (.A(net506),
    .X(net505));
 sg13g2_buf_8 fanout506 (.A(net510),
    .X(net506));
 sg13g2_buf_8 fanout507 (.A(net510),
    .X(net507));
 sg13g2_buf_8 fanout508 (.A(net509),
    .X(net508));
 sg13g2_buf_8 fanout509 (.A(net510),
    .X(net509));
 sg13g2_buf_8 fanout510 (.A(net515),
    .X(net510));
 sg13g2_buf_8 fanout511 (.A(net512),
    .X(net511));
 sg13g2_buf_8 fanout512 (.A(net515),
    .X(net512));
 sg13g2_buf_8 fanout513 (.A(net514),
    .X(net513));
 sg13g2_buf_8 fanout514 (.A(net515),
    .X(net514));
 sg13g2_buf_8 fanout515 (.A(net516),
    .X(net515));
 sg13g2_buf_8 fanout516 (.A(_0904_),
    .X(net516));
 sg13g2_buf_8 fanout517 (.A(net518),
    .X(net517));
 sg13g2_buf_8 fanout518 (.A(_0900_),
    .X(net518));
 sg13g2_buf_8 fanout519 (.A(_0898_),
    .X(net519));
 sg13g2_buf_8 fanout520 (.A(_0896_),
    .X(net520));
 sg13g2_buf_8 fanout521 (.A(_0894_),
    .X(net521));
 sg13g2_buf_8 fanout522 (.A(_0892_),
    .X(net522));
 sg13g2_buf_8 fanout523 (.A(_0890_),
    .X(net523));
 sg13g2_buf_8 fanout524 (.A(_0888_),
    .X(net524));
 sg13g2_buf_8 fanout525 (.A(_0886_),
    .X(net525));
 sg13g2_buf_8 fanout526 (.A(_0822_),
    .X(net526));
 sg13g2_buf_8 fanout527 (.A(net529),
    .X(net527));
 sg13g2_buf_1 fanout528 (.A(net529),
    .X(net528));
 sg13g2_buf_8 fanout529 (.A(_0821_),
    .X(net529));
 sg13g2_buf_8 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_8 fanout531 (.A(_0820_),
    .X(net531));
 sg13g2_buf_8 fanout532 (.A(net533),
    .X(net532));
 sg13g2_buf_8 fanout533 (.A(net1067),
    .X(net533));
 sg13g2_buf_8 fanout534 (.A(net1076),
    .X(net534));
 sg13g2_buf_8 fanout535 (.A(\u_tree_core.current_node_q[1] ),
    .X(net535));
 sg13g2_buf_8 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_8 fanout537 (.A(net538),
    .X(net537));
 sg13g2_buf_8 fanout538 (.A(\u_tree_core.current_node_q[0] ),
    .X(net538));
 sg13g2_buf_8 fanout539 (.A(net540),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(net541),
    .X(net540));
 sg13g2_buf_1 fanout541 (.A(net542),
    .X(net541));
 sg13g2_buf_1 fanout542 (.A(\u_tree_core.current_node_q[0] ),
    .X(net542));
 sg13g2_buf_8 fanout543 (.A(\u_feature_loader.feature_idx_q[2] ),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(net1075),
    .X(net544));
 sg13g2_buf_8 fanout545 (.A(net1072),
    .X(net545));
 sg13g2_buf_8 fanout546 (.A(\u_model_loader.byte_idx_q[4] ),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(net561),
    .X(net547));
 sg13g2_buf_8 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(net1070),
    .X(net549));
 sg13g2_buf_8 fanout550 (.A(\model_byte[2] ),
    .X(net550));
 sg13g2_buf_8 fanout551 (.A(\model_byte[1] ),
    .X(net551));
 sg13g2_buf_8 fanout552 (.A(\model_byte[0] ),
    .X(net552));
 sg13g2_buf_8 fanout553 (.A(net556),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(net556),
    .X(net554));
 sg13g2_buf_1 fanout555 (.A(net556),
    .X(net555));
 sg13g2_buf_8 fanout556 (.A(rst_n),
    .X(net556));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[2]),
    .X(net12));
 sg13g2_tielo tt_um_pgfarley_tophat_top_13 (.L_LO(net13));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_leaf_38_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\node_left_flat[23] ),
    .X(net335));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0144_),
    .X(net336));
 sg13g2_dlygate4sd3_1 hold3 (.A(\node_left_flat[7] ),
    .X(net337));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0128_),
    .X(net338));
 sg13g2_dlygate4sd3_1 hold5 (.A(\feature_vector_flat[6] ),
    .X(net339));
 sg13g2_dlygate4sd3_1 hold6 (.A(_0237_),
    .X(net340));
 sg13g2_dlygate4sd3_1 hold7 (.A(\node_right_flat[27] ),
    .X(net341));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0120_),
    .X(net342));
 sg13g2_dlygate4sd3_1 hold9 (.A(\node_right_flat[3] ),
    .X(net343));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0096_),
    .X(net344));
 sg13g2_dlygate4sd3_1 hold11 (.A(\node_threshold_flat[35] ),
    .X(net345));
 sg13g2_dlygate4sd3_1 hold12 (.A(\feature_vector_flat[0] ),
    .X(net346));
 sg13g2_dlygate4sd3_1 hold13 (.A(_0231_),
    .X(net347));
 sg13g2_dlygate4sd3_1 hold14 (.A(\feature_vector_flat[2] ),
    .X(net348));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0233_),
    .X(net349));
 sg13g2_dlygate4sd3_1 hold16 (.A(\node_threshold_flat[36] ),
    .X(net350));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0185_),
    .X(net351));
 sg13g2_dlygate4sd3_1 hold18 (.A(\node_right_flat[19] ),
    .X(net352));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0112_),
    .X(net353));
 sg13g2_dlygate4sd3_1 hold20 (.A(\node_threshold_flat[37] ),
    .X(net354));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0186_),
    .X(net355));
 sg13g2_dlygate4sd3_1 hold22 (.A(\node_threshold_flat[16] ),
    .X(net356));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0543_),
    .X(net357));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0165_),
    .X(net358));
 sg13g2_dlygate4sd3_1 hold25 (.A(\node_threshold_flat[38] ),
    .X(net359));
 sg13g2_dlygate4sd3_1 hold26 (.A(_0187_),
    .X(net360));
 sg13g2_dlygate4sd3_1 hold27 (.A(\feature_vector_flat[37] ),
    .X(net361));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0268_),
    .X(net362));
 sg13g2_dlygate4sd3_1 hold29 (.A(\node_threshold_flat[3] ),
    .X(net363));
 sg13g2_dlygate4sd3_1 hold30 (.A(\feature_vector_flat[33] ),
    .X(net364));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0264_),
    .X(net365));
 sg13g2_dlygate4sd3_1 hold32 (.A(\node_right_flat[7] ),
    .X(net366));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0100_),
    .X(net367));
 sg13g2_dlygate4sd3_1 hold34 (.A(\node_left_flat[3] ),
    .X(net368));
 sg13g2_dlygate4sd3_1 hold35 (.A(_0124_),
    .X(net369));
 sg13g2_dlygate4sd3_1 hold36 (.A(\node_left_flat[27] ),
    .X(net370));
 sg13g2_dlygate4sd3_1 hold37 (.A(_0148_),
    .X(net371));
 sg13g2_dlygate4sd3_1 hold38 (.A(\node_threshold_flat[17] ),
    .X(net372));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0166_),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold40 (.A(\node_threshold_flat[11] ),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold41 (.A(_0160_),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold42 (.A(\feature_vector_flat[39] ),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold43 (.A(_0270_),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold44 (.A(\node_right_flat[23] ),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0116_),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u_model_loader.byte_idx_q[0] ),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0023_),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold48 (.A(\feature_vector_flat[3] ),
    .X(net563));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0234_),
    .X(net564));
 sg13g2_dlygate4sd3_1 hold50 (.A(\node_threshold_flat[39] ),
    .X(net565));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0188_),
    .X(net566));
 sg13g2_dlygate4sd3_1 hold52 (.A(\node_threshold_flat[51] ),
    .X(net567));
 sg13g2_dlygate4sd3_1 hold53 (.A(\node_left_flat[19] ),
    .X(net568));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0140_),
    .X(net569));
 sg13g2_dlygate4sd3_1 hold55 (.A(\node_threshold_flat[43] ),
    .X(net570));
 sg13g2_dlygate4sd3_1 hold56 (.A(\feature_vector_flat[32] ),
    .X(net571));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0263_),
    .X(net572));
 sg13g2_dlygate4sd3_1 hold58 (.A(\feature_vector_flat[35] ),
    .X(net573));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0266_),
    .X(net574));
 sg13g2_dlygate4sd3_1 hold60 (.A(\feature_vector_flat[36] ),
    .X(net575));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0267_),
    .X(net576));
 sg13g2_dlygate4sd3_1 hold62 (.A(\node_threshold_flat[6] ),
    .X(net577));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0155_),
    .X(net578));
 sg13g2_dlygate4sd3_1 hold64 (.A(\feature_vector_flat[34] ),
    .X(net579));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0265_),
    .X(net580));
 sg13g2_dlygate4sd3_1 hold66 (.A(\node_threshold_flat[18] ),
    .X(net581));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0167_),
    .X(net582));
 sg13g2_dlygate4sd3_1 hold68 (.A(\feature_vector_flat[38] ),
    .X(net583));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0269_),
    .X(net584));
 sg13g2_dlygate4sd3_1 hold70 (.A(\node_threshold_flat[8] ),
    .X(net585));
 sg13g2_dlygate4sd3_1 hold71 (.A(feature_byte_valid),
    .X(net586));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0227_),
    .X(net587));
 sg13g2_dlygate4sd3_1 hold73 (.A(\feature_vector_flat[4] ),
    .X(net588));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0235_),
    .X(net589));
 sg13g2_dlygate4sd3_1 hold75 (.A(\node_left_flat[5] ),
    .X(net590));
 sg13g2_dlygate4sd3_1 hold76 (.A(\feature_vector_flat[5] ),
    .X(net591));
 sg13g2_dlygate4sd3_1 hold77 (.A(_0236_),
    .X(net592));
 sg13g2_dlygate4sd3_1 hold78 (.A(\u_tree_core.depth_q[1] ),
    .X(net593));
 sg13g2_dlygate4sd3_1 hold79 (.A(_0813_),
    .X(net594));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0307_),
    .X(net595));
 sg13g2_dlygate4sd3_1 hold81 (.A(\node_left_flat[26] ),
    .X(net596));
 sg13g2_dlygate4sd3_1 hold82 (.A(\node_left_flat[14] ),
    .X(net597));
 sg13g2_dlygate4sd3_1 hold83 (.A(_0500_),
    .X(net598));
 sg13g2_dlygate4sd3_1 hold84 (.A(\node_threshold_flat[4] ),
    .X(net599));
 sg13g2_dlygate4sd3_1 hold85 (.A(_0153_),
    .X(net600));
 sg13g2_dlygate4sd3_1 hold86 (.A(\node_threshold_flat[19] ),
    .X(net601));
 sg13g2_dlygate4sd3_1 hold87 (.A(_0168_),
    .X(net602));
 sg13g2_dlygate4sd3_1 hold88 (.A(\node_left_flat[15] ),
    .X(net603));
 sg13g2_dlygate4sd3_1 hold89 (.A(_0136_),
    .X(net604));
 sg13g2_dlygate4sd3_1 hold90 (.A(\node_threshold_flat[40] ),
    .X(net605));
 sg13g2_dlygate4sd3_1 hold91 (.A(\node_threshold_flat[50] ),
    .X(net606));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0199_),
    .X(net607));
 sg13g2_dlygate4sd3_1 hold93 (.A(\node_feature_flat[5] ),
    .X(net608));
 sg13g2_dlygate4sd3_1 hold94 (.A(\node_threshold_flat[5] ),
    .X(net609));
 sg13g2_dlygate4sd3_1 hold95 (.A(_0154_),
    .X(net610));
 sg13g2_dlygate4sd3_1 hold96 (.A(\node_feature_flat[15] ),
    .X(net611));
 sg13g2_dlygate4sd3_1 hold97 (.A(_0220_),
    .X(net612));
 sg13g2_dlygate4sd3_1 hold98 (.A(\node_threshold_flat[42] ),
    .X(net613));
 sg13g2_dlygate4sd3_1 hold99 (.A(\node_left_flat[25] ),
    .X(net614));
 sg13g2_dlygate4sd3_1 hold100 (.A(_0514_),
    .X(net615));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0146_),
    .X(net616));
 sg13g2_dlygate4sd3_1 hold102 (.A(\feature_vector_flat[7] ),
    .X(net617));
 sg13g2_dlygate4sd3_1 hold103 (.A(_0238_),
    .X(net618));
 sg13g2_dlygate4sd3_1 hold104 (.A(\feature_vector_flat[46] ),
    .X(net619));
 sg13g2_dlygate4sd3_1 hold105 (.A(_0724_),
    .X(net620));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0277_),
    .X(net621));
 sg13g2_dlygate4sd3_1 hold107 (.A(\node_feature_flat[17] ),
    .X(net622));
 sg13g2_dlygate4sd3_1 hold108 (.A(\node_feature_flat[3] ),
    .X(net623));
 sg13g2_dlygate4sd3_1 hold109 (.A(\node_feature_flat[16] ),
    .X(net624));
 sg13g2_dlygate4sd3_1 hold110 (.A(\feature_vector_flat[41] ),
    .X(net625));
 sg13g2_dlygate4sd3_1 hold111 (.A(_0719_),
    .X(net626));
 sg13g2_dlygate4sd3_1 hold112 (.A(\node_left_flat[21] ),
    .X(net627));
 sg13g2_dlygate4sd3_1 hold113 (.A(\node_left_flat[4] ),
    .X(net628));
 sg13g2_dlygate4sd3_1 hold114 (.A(\node_left_flat[24] ),
    .X(net629));
 sg13g2_dlygate4sd3_1 hold115 (.A(_0145_),
    .X(net630));
 sg13g2_dlygate4sd3_1 hold116 (.A(\feature_vector_flat[1] ),
    .X(net631));
 sg13g2_dlygate4sd3_1 hold117 (.A(_0232_),
    .X(net632));
 sg13g2_dlygate4sd3_1 hold118 (.A(\feature_vector_flat[47] ),
    .X(net633));
 sg13g2_dlygate4sd3_1 hold119 (.A(_0725_),
    .X(net634));
 sg13g2_dlygate4sd3_1 hold120 (.A(\node_threshold_flat[49] ),
    .X(net635));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0588_),
    .X(net636));
 sg13g2_dlygate4sd3_1 hold122 (.A(\node_left_flat[17] ),
    .X(net637));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0138_),
    .X(net638));
 sg13g2_dlygate4sd3_1 hold124 (.A(\node_threshold_flat[55] ),
    .X(net639));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0594_),
    .X(net640));
 sg13g2_dlygate4sd3_1 hold126 (.A(_0204_),
    .X(net641));
 sg13g2_dlygate4sd3_1 hold127 (.A(\node_left_flat[11] ),
    .X(net642));
 sg13g2_dlygate4sd3_1 hold128 (.A(\u_feature_loader.feature_idx_q[3] ),
    .X(net643));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0230_),
    .X(net644));
 sg13g2_dlygate4sd3_1 hold130 (.A(\feature_vector_flat[43] ),
    .X(net645));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0721_),
    .X(net646));
 sg13g2_dlygate4sd3_1 hold132 (.A(\node_threshold_flat[9] ),
    .X(net647));
 sg13g2_dlygate4sd3_1 hold133 (.A(\node_left_flat[6] ),
    .X(net648));
 sg13g2_dlygate4sd3_1 hold134 (.A(\node_threshold_flat[54] ),
    .X(net649));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0593_),
    .X(net650));
 sg13g2_dlygate4sd3_1 hold136 (.A(\node_left_flat[20] ),
    .X(net651));
 sg13g2_dlygate4sd3_1 hold137 (.A(\feature_vector_flat[40] ),
    .X(net652));
 sg13g2_dlygate4sd3_1 hold138 (.A(_0718_),
    .X(net653));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0271_),
    .X(net654));
 sg13g2_dlygate4sd3_1 hold140 (.A(\node_feature_flat[18] ),
    .X(net655));
 sg13g2_dlygate4sd3_1 hold141 (.A(\feature_vector_flat[45] ),
    .X(net656));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0723_),
    .X(net657));
 sg13g2_dlygate4sd3_1 hold143 (.A(_0276_),
    .X(net658));
 sg13g2_dlygate4sd3_1 hold144 (.A(\node_threshold_flat[10] ),
    .X(net659));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0159_),
    .X(net660));
 sg13g2_dlygate4sd3_1 hold146 (.A(\node_threshold_flat[34] ),
    .X(net661));
 sg13g2_dlygate4sd3_1 hold147 (.A(\node_threshold_flat[32] ),
    .X(net662));
 sg13g2_dlygate4sd3_1 hold148 (.A(\node_feature_flat[20] ),
    .X(net663));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0225_),
    .X(net664));
 sg13g2_dlygate4sd3_1 hold150 (.A(\node_feature_flat[10] ),
    .X(net665));
 sg13g2_dlygate4sd3_1 hold151 (.A(_0615_),
    .X(net666));
 sg13g2_dlygate4sd3_1 hold152 (.A(\node_threshold_flat[41] ),
    .X(net667));
 sg13g2_dlygate4sd3_1 hold153 (.A(\node_left_flat[13] ),
    .X(net668));
 sg13g2_dlygate4sd3_1 hold154 (.A(_0499_),
    .X(net669));
 sg13g2_dlygate4sd3_1 hold155 (.A(\node_left_flat[22] ),
    .X(net670));
 sg13g2_dlygate4sd3_1 hold156 (.A(\node_threshold_flat[7] ),
    .X(net671));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0156_),
    .X(net672));
 sg13g2_dlygate4sd3_1 hold158 (.A(\node_threshold_flat[52] ),
    .X(net673));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0591_),
    .X(net674));
 sg13g2_dlygate4sd3_1 hold160 (.A(\node_threshold_flat[48] ),
    .X(net675));
 sg13g2_dlygate4sd3_1 hold161 (.A(\feature_vector_flat[44] ),
    .X(net676));
 sg13g2_dlygate4sd3_1 hold162 (.A(_0722_),
    .X(net677));
 sg13g2_dlygate4sd3_1 hold163 (.A(\node_left_flat[16] ),
    .X(net678));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0137_),
    .X(net679));
 sg13g2_dlygate4sd3_1 hold165 (.A(\node_left_flat[18] ),
    .X(net680));
 sg13g2_dlygate4sd3_1 hold166 (.A(\node_feature_flat[9] ),
    .X(net681));
 sg13g2_dlygate4sd3_1 hold167 (.A(_0614_),
    .X(net682));
 sg13g2_dlygate4sd3_1 hold168 (.A(\node_feature_flat[13] ),
    .X(net683));
 sg13g2_dlygate4sd3_1 hold169 (.A(_0218_),
    .X(net684));
 sg13g2_dlygate4sd3_1 hold170 (.A(\node_feature_flat[4] ),
    .X(net685));
 sg13g2_dlygate4sd3_1 hold171 (.A(\node_left_flat[12] ),
    .X(net686));
 sg13g2_dlygate4sd3_1 hold172 (.A(_0498_),
    .X(net687));
 sg13g2_dlygate4sd3_1 hold173 (.A(core_busy),
    .X(net688));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0752_),
    .X(net689));
 sg13g2_dlygate4sd3_1 hold175 (.A(_0296_),
    .X(net690));
 sg13g2_dlygate4sd3_1 hold176 (.A(uo_out[7]),
    .X(net691));
 sg13g2_dlygate4sd3_1 hold177 (.A(_0304_),
    .X(net692));
 sg13g2_dlygate4sd3_1 hold178 (.A(\node_threshold_flat[33] ),
    .X(net693));
 sg13g2_dlygate4sd3_1 hold179 (.A(\node_threshold_flat[53] ),
    .X(net694));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0592_),
    .X(net695));
 sg13g2_dlygate4sd3_1 hold181 (.A(\node_feature_flat[19] ),
    .X(net696));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0627_),
    .X(net697));
 sg13g2_dlygate4sd3_1 hold183 (.A(uo_out[4]),
    .X(net698));
 sg13g2_dlygate4sd3_1 hold184 (.A(_0301_),
    .X(net699));
 sg13g2_dlygate4sd3_1 hold185 (.A(\node_threshold_flat[46] ),
    .X(net700));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0584_),
    .X(net701));
 sg13g2_dlygate4sd3_1 hold187 (.A(_0195_),
    .X(net702));
 sg13g2_dlygate4sd3_1 hold188 (.A(\feature_vector_flat[42] ),
    .X(net703));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0720_),
    .X(net704));
 sg13g2_dlygate4sd3_1 hold190 (.A(\node_feature_flat[11] ),
    .X(net705));
 sg13g2_dlygate4sd3_1 hold191 (.A(_0616_),
    .X(net706));
 sg13g2_dlygate4sd3_1 hold192 (.A(\node_right_flat[26] ),
    .X(net707));
 sg13g2_dlygate4sd3_1 hold193 (.A(\node_threshold_flat[1] ),
    .X(net708));
 sg13g2_dlygate4sd3_1 hold194 (.A(\node_feature_flat[14] ),
    .X(net709));
 sg13g2_dlygate4sd3_1 hold195 (.A(\node_feature_flat[12] ),
    .X(net710));
 sg13g2_dlygate4sd3_1 hold196 (.A(\node_threshold_flat[15] ),
    .X(net711));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0541_),
    .X(net712));
 sg13g2_dlygate4sd3_1 hold198 (.A(\node_right_flat[25] ),
    .X(net713));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0472_),
    .X(net714));
 sg13g2_dlygate4sd3_1 hold200 (.A(\feature_vector_flat[62] ),
    .X(net715));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0750_),
    .X(net716));
 sg13g2_dlygate4sd3_1 hold202 (.A(_0293_),
    .X(net717));
 sg13g2_dlygate4sd3_1 hold203 (.A(\feature_vector_flat[60] ),
    .X(net718));
 sg13g2_dlygate4sd3_1 hold204 (.A(_0748_),
    .X(net719));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0291_),
    .X(net720));
 sg13g2_dlygate4sd3_1 hold206 (.A(\node_right_flat[14] ),
    .X(net721));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0445_),
    .X(net722));
 sg13g2_dlygate4sd3_1 hold208 (.A(uo_out[5]),
    .X(net723));
 sg13g2_dlygate4sd3_1 hold209 (.A(_0302_),
    .X(net724));
 sg13g2_dlygate4sd3_1 hold210 (.A(\node_right_flat[1] ),
    .X(net725));
 sg13g2_dlygate4sd3_1 hold211 (.A(\node_feature_flat[2] ),
    .X(net726));
 sg13g2_dlygate4sd3_1 hold212 (.A(\node_right_flat[15] ),
    .X(net727));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0448_),
    .X(net728));
 sg13g2_dlygate4sd3_1 hold214 (.A(uo_out[1]),
    .X(net729));
 sg13g2_dlygate4sd3_1 hold215 (.A(_0298_),
    .X(net730));
 sg13g2_dlygate4sd3_1 hold216 (.A(\node_threshold_flat[23] ),
    .X(net731));
 sg13g2_dlygate4sd3_1 hold217 (.A(_0557_),
    .X(net732));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0172_),
    .X(net733));
 sg13g2_dlygate4sd3_1 hold219 (.A(\feature_vector_flat[30] ),
    .X(net734));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0695_),
    .X(net735));
 sg13g2_dlygate4sd3_1 hold221 (.A(_0261_),
    .X(net736));
 sg13g2_dlygate4sd3_1 hold222 (.A(\node_right_flat[11] ),
    .X(net737));
 sg13g2_dlygate4sd3_1 hold223 (.A(core_error),
    .X(net738));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0305_),
    .X(net739));
 sg13g2_dlygate4sd3_1 hold225 (.A(\node_right_flat[12] ),
    .X(net740));
 sg13g2_dlygate4sd3_1 hold226 (.A(_0441_),
    .X(net741));
 sg13g2_dlygate4sd3_1 hold227 (.A(\node_feature_flat[0] ),
    .X(net742));
 sg13g2_dlygate4sd3_1 hold228 (.A(\feature_vector_flat[28] ),
    .X(net743));
 sg13g2_dlygate4sd3_1 hold229 (.A(_0691_),
    .X(net744));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0259_),
    .X(net745));
 sg13g2_dlygate4sd3_1 hold231 (.A(\node_threshold_flat[14] ),
    .X(net746));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0539_),
    .X(net747));
 sg13g2_dlygate4sd3_1 hold233 (.A(uo_out[2]),
    .X(net748));
 sg13g2_dlygate4sd3_1 hold234 (.A(_0299_),
    .X(net749));
 sg13g2_dlygate4sd3_1 hold235 (.A(\feature_vector_flat[61] ),
    .X(net750));
 sg13g2_dlygate4sd3_1 hold236 (.A(_0749_),
    .X(net751));
 sg13g2_dlygate4sd3_1 hold237 (.A(\node_threshold_flat[21] ),
    .X(net752));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0553_),
    .X(net753));
 sg13g2_dlygate4sd3_1 hold239 (.A(\feature_vector_flat[63] ),
    .X(net754));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0751_),
    .X(net755));
 sg13g2_dlygate4sd3_1 hold241 (.A(\node_feature_flat[1] ),
    .X(net756));
 sg13g2_dlygate4sd3_1 hold242 (.A(\node_right_flat[13] ),
    .X(net757));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0443_),
    .X(net758));
 sg13g2_dlygate4sd3_1 hold244 (.A(\node_threshold_flat[44] ),
    .X(net759));
 sg13g2_dlygate4sd3_1 hold245 (.A(_0582_),
    .X(net760));
 sg13g2_dlygate4sd3_1 hold246 (.A(uo_out[6]),
    .X(net761));
 sg13g2_dlygate4sd3_1 hold247 (.A(_0303_),
    .X(net762));
 sg13g2_dlygate4sd3_1 hold248 (.A(\feature_vector_flat[59] ),
    .X(net763));
 sg13g2_dlygate4sd3_1 hold249 (.A(_0747_),
    .X(net764));
 sg13g2_dlygate4sd3_1 hold250 (.A(\node_right_flat[20] ),
    .X(net765));
 sg13g2_dlygate4sd3_1 hold251 (.A(_0113_),
    .X(net766));
 sg13g2_dlygate4sd3_1 hold252 (.A(\node_right_flat[16] ),
    .X(net767));
 sg13g2_dlygate4sd3_1 hold253 (.A(_0109_),
    .X(net768));
 sg13g2_dlygate4sd3_1 hold254 (.A(\node_threshold_flat[2] ),
    .X(net769));
 sg13g2_dlygate4sd3_1 hold255 (.A(\node_left_flat[2] ),
    .X(net770));
 sg13g2_dlygate4sd3_1 hold256 (.A(\feature_vector_flat[58] ),
    .X(net771));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0746_),
    .X(net772));
 sg13g2_dlygate4sd3_1 hold258 (.A(_0289_),
    .X(net773));
 sg13g2_dlygate4sd3_1 hold259 (.A(\node_right_flat[2] ),
    .X(net774));
 sg13g2_dlygate4sd3_1 hold260 (.A(\node_right_flat[5] ),
    .X(net775));
 sg13g2_dlygate4sd3_1 hold261 (.A(\node_threshold_flat[0] ),
    .X(net776));
 sg13g2_dlygate4sd3_1 hold262 (.A(\node_threshold_flat[47] ),
    .X(net777));
 sg13g2_dlygate4sd3_1 hold263 (.A(_0585_),
    .X(net778));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0196_),
    .X(net779));
 sg13g2_dlygate4sd3_1 hold265 (.A(\node_threshold_flat[20] ),
    .X(net780));
 sg13g2_dlygate4sd3_1 hold266 (.A(_0551_),
    .X(net781));
 sg13g2_dlygate4sd3_1 hold267 (.A(\node_right_flat[17] ),
    .X(net782));
 sg13g2_dlygate4sd3_1 hold268 (.A(_0110_),
    .X(net783));
 sg13g2_dlygate4sd3_1 hold269 (.A(\feature_vector_flat[8] ),
    .X(net784));
 sg13g2_dlygate4sd3_1 hold270 (.A(_0647_),
    .X(net785));
 sg13g2_dlygate4sd3_1 hold271 (.A(\node_right_flat[22] ),
    .X(net786));
 sg13g2_dlygate4sd3_1 hold272 (.A(\node_threshold_flat[45] ),
    .X(net787));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0583_),
    .X(net788));
 sg13g2_dlygate4sd3_1 hold274 (.A(_0194_),
    .X(net789));
 sg13g2_dlygate4sd3_1 hold275 (.A(\node_right_flat[24] ),
    .X(net790));
 sg13g2_dlygate4sd3_1 hold276 (.A(\feature_vector_flat[27] ),
    .X(net791));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0689_),
    .X(net792));
 sg13g2_dlygate4sd3_1 hold278 (.A(\node_right_flat[0] ),
    .X(net793));
 sg13g2_dlygate4sd3_1 hold279 (.A(\feature_vector_flat[14] ),
    .X(net794));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0659_),
    .X(net795));
 sg13g2_dlygate4sd3_1 hold281 (.A(_0245_),
    .X(net796));
 sg13g2_dlygate4sd3_1 hold282 (.A(\feature_vector_flat[10] ),
    .X(net797));
 sg13g2_dlygate4sd3_1 hold283 (.A(_0651_),
    .X(net798));
 sg13g2_dlygate4sd3_1 hold284 (.A(\feature_vector_flat[15] ),
    .X(net799));
 sg13g2_dlygate4sd3_1 hold285 (.A(_0661_),
    .X(net800));
 sg13g2_dlygate4sd3_1 hold286 (.A(\feature_vector_flat[9] ),
    .X(net801));
 sg13g2_dlygate4sd3_1 hold287 (.A(_0649_),
    .X(net802));
 sg13g2_dlygate4sd3_1 hold288 (.A(\node_threshold_flat[22] ),
    .X(net803));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0555_),
    .X(net804));
 sg13g2_dlygate4sd3_1 hold290 (.A(\node_threshold_flat[12] ),
    .X(net805));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0535_),
    .X(net806));
 sg13g2_dlygate4sd3_1 hold292 (.A(\node_left_flat[1] ),
    .X(net807));
 sg13g2_dlygate4sd3_1 hold293 (.A(\feature_vector_flat[26] ),
    .X(net808));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0687_),
    .X(net809));
 sg13g2_dlygate4sd3_1 hold295 (.A(\node_right_flat[6] ),
    .X(net810));
 sg13g2_dlygate4sd3_1 hold296 (.A(\feature_vector_flat[13] ),
    .X(net811));
 sg13g2_dlygate4sd3_1 hold297 (.A(_0657_),
    .X(net812));
 sg13g2_dlygate4sd3_1 hold298 (.A(\node_right_flat[18] ),
    .X(net813));
 sg13g2_dlygate4sd3_1 hold299 (.A(\feature_vector_flat[29] ),
    .X(net814));
 sg13g2_dlygate4sd3_1 hold300 (.A(_0693_),
    .X(net815));
 sg13g2_dlygate4sd3_1 hold301 (.A(\feature_vector_flat[55] ),
    .X(net816));
 sg13g2_dlygate4sd3_1 hold302 (.A(_0286_),
    .X(net817));
 sg13g2_dlygate4sd3_1 hold303 (.A(uo_out[3]),
    .X(net818));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0300_),
    .X(net819));
 sg13g2_dlygate4sd3_1 hold305 (.A(\leaf_value_flat[62] ),
    .X(net820));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0091_),
    .X(net821));
 sg13g2_dlygate4sd3_1 hold307 (.A(\leaf_value_flat[28] ),
    .X(net822));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0057_),
    .X(net823));
 sg13g2_dlygate4sd3_1 hold309 (.A(\leaf_value_flat[14] ),
    .X(net824));
 sg13g2_dlygate4sd3_1 hold310 (.A(_0043_),
    .X(net825));
 sg13g2_dlygate4sd3_1 hold311 (.A(\node_right_flat[21] ),
    .X(net826));
 sg13g2_dlygate4sd3_1 hold312 (.A(_0114_),
    .X(net827));
 sg13g2_dlygate4sd3_1 hold313 (.A(\leaf_value_flat[45] ),
    .X(net828));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0074_),
    .X(net829));
 sg13g2_dlygate4sd3_1 hold315 (.A(\leaf_value_flat[60] ),
    .X(net830));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0089_),
    .X(net831));
 sg13g2_dlygate4sd3_1 hold317 (.A(\feature_vector_flat[12] ),
    .X(net832));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0655_),
    .X(net833));
 sg13g2_dlygate4sd3_1 hold319 (.A(\leaf_value_flat[35] ),
    .X(net834));
 sg13g2_dlygate4sd3_1 hold320 (.A(\node_threshold_flat[13] ),
    .X(net835));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0537_),
    .X(net836));
 sg13g2_dlygate4sd3_1 hold322 (.A(\leaf_value_flat[39] ),
    .X(net837));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0068_),
    .X(net838));
 sg13g2_dlygate4sd3_1 hold324 (.A(\leaf_value_flat[46] ),
    .X(net839));
 sg13g2_dlygate4sd3_1 hold325 (.A(_0075_),
    .X(net840));
 sg13g2_dlygate4sd3_1 hold326 (.A(\leaf_value_flat[38] ),
    .X(net841));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0067_),
    .X(net842));
 sg13g2_dlygate4sd3_1 hold328 (.A(\leaf_value_flat[37] ),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold329 (.A(_0066_),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold330 (.A(uo_out[0]),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold331 (.A(\leaf_value_flat[33] ),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0062_),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold333 (.A(\node_left_flat[0] ),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold334 (.A(\feature_vector_flat[49] ),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0280_),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold336 (.A(\node_right_flat[4] ),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold337 (.A(\leaf_value_flat[10] ),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0039_),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold339 (.A(\leaf_value_flat[57] ),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold340 (.A(_0086_),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold341 (.A(\leaf_value_flat[6] ),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold342 (.A(_0035_),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold343 (.A(\feature_vector_flat[53] ),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold344 (.A(_0284_),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold345 (.A(\leaf_value_flat[18] ),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0047_),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold347 (.A(\feature_vector_flat[56] ),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0744_),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold349 (.A(_0287_),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold350 (.A(\leaf_value_flat[4] ),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold351 (.A(_0033_),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold352 (.A(\leaf_value_flat[48] ),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold353 (.A(_0077_),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold354 (.A(\feature_vector_flat[24] ),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0683_),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold356 (.A(\leaf_value_flat[51] ),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold357 (.A(\leaf_value_flat[15] ),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold358 (.A(_0044_),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold359 (.A(\feature_vector_flat[31] ),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0697_),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold361 (.A(\leaf_value_flat[59] ),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold362 (.A(_0088_),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold363 (.A(\leaf_value_flat[42] ),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold364 (.A(_0071_),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold365 (.A(\u_model_loader.byte_idx_q[1] ),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold366 (.A(_1156_),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0024_),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold368 (.A(\leaf_value_flat[27] ),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold369 (.A(\feature_vector_flat[11] ),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold370 (.A(_0653_),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold371 (.A(\leaf_value_flat[32] ),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold372 (.A(_0061_),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold373 (.A(\leaf_value_flat[40] ),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold374 (.A(_0069_),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold375 (.A(\leaf_value_flat[5] ),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold376 (.A(_0034_),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold377 (.A(\feature_vector_flat[25] ),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0685_),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold379 (.A(\leaf_value_flat[44] ),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0073_),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold381 (.A(\node_right_flat[8] ),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0431_),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold383 (.A(_0101_),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold384 (.A(\feature_vector_flat[17] ),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold385 (.A(_0248_),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold386 (.A(\leaf_value_flat[21] ),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold387 (.A(_0050_),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold388 (.A(\leaf_value_flat[47] ),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold389 (.A(_0076_),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold390 (.A(\node_left_flat[10] ),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold391 (.A(_0131_),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold392 (.A(\node_right_flat[9] ),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold393 (.A(_0433_),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0102_),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold395 (.A(\leaf_value_flat[41] ),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0070_),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold397 (.A(\feature_vector_flat[21] ),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0252_),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold399 (.A(\leaf_value_flat[8] ),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold400 (.A(_0037_),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold401 (.A(\feature_vector_flat[57] ),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold402 (.A(_0745_),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold403 (.A(\leaf_value_flat[36] ),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold404 (.A(_0065_),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold405 (.A(model_loaded),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0226_),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold407 (.A(\feature_vector_flat[51] ),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold408 (.A(_0282_),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold409 (.A(\leaf_value_flat[55] ),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold410 (.A(_0084_),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold411 (.A(\leaf_value_flat[2] ),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold412 (.A(_0031_),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold413 (.A(\leaf_value_flat[49] ),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold414 (.A(_0078_),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold415 (.A(\leaf_value_flat[63] ),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0092_),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold417 (.A(\leaf_value_flat[61] ),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold418 (.A(_0090_),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold419 (.A(\leaf_value_flat[17] ),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0046_),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold421 (.A(\leaf_value_flat[34] ),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold422 (.A(_0063_),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold423 (.A(\leaf_value_flat[22] ),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold424 (.A(_0051_),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold425 (.A(\node_threshold_flat[24] ),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold426 (.A(_0173_),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold427 (.A(\leaf_value_flat[53] ),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold428 (.A(_0082_),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold429 (.A(\leaf_value_flat[3] ),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold430 (.A(\leaf_value_flat[11] ),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold431 (.A(\node_threshold_flat[27] ),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold432 (.A(\leaf_value_flat[54] ),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold433 (.A(_0083_),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold434 (.A(\leaf_value_flat[19] ),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold435 (.A(\feature_vector_flat[23] ),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold436 (.A(_0254_),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold437 (.A(\feature_vector_flat[20] ),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold438 (.A(_0251_),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold439 (.A(\leaf_value_flat[56] ),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold440 (.A(_0085_),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold441 (.A(\leaf_value_flat[20] ),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold442 (.A(_0049_),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold443 (.A(\leaf_value_flat[30] ),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold444 (.A(_0059_),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold445 (.A(\node_feature_flat[8] ),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold446 (.A(_0213_),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold447 (.A(\leaf_value_flat[26] ),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold448 (.A(_0055_),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold449 (.A(\feature_vector_flat[50] ),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0281_),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold451 (.A(\leaf_value_flat[0] ),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0029_),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold453 (.A(\leaf_value_flat[1] ),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold454 (.A(_0030_),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold455 (.A(\node_left_flat[9] ),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0130_),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold457 (.A(\u_model_loader.byte_idx_q[5] ),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold458 (.A(_0331_),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold459 (.A(\feature_vector_flat[16] ),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0247_),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold461 (.A(\u_feature_loader.feature_idx_q[1] ),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold462 (.A(_0631_),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold463 (.A(\node_feature_flat[7] ),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold464 (.A(_0212_),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold465 (.A(\leaf_value_flat[7] ),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0036_),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold467 (.A(\leaf_value_flat[31] ),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold468 (.A(_0060_),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold469 (.A(\leaf_value_flat[52] ),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold470 (.A(_0081_),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold471 (.A(\node_threshold_flat[25] ),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold472 (.A(_0174_),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold473 (.A(\feature_vector_flat[19] ),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0250_),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold475 (.A(\leaf_value_flat[50] ),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0079_),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold477 (.A(\node_threshold_flat[31] ),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0180_),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold479 (.A(\feature_vector_flat[22] ),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold480 (.A(_0253_),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold481 (.A(\leaf_value_flat[43] ),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold482 (.A(\feature_vector_flat[52] ),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold483 (.A(_0737_),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0283_),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold485 (.A(\leaf_value_flat[58] ),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0087_),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold487 (.A(\leaf_value_flat[12] ),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0041_),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold489 (.A(\node_right_flat[10] ),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0435_),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold491 (.A(_0103_),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold492 (.A(\node_threshold_flat[26] ),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold493 (.A(_0175_),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold494 (.A(\leaf_value_flat[16] ),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0045_),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold496 (.A(\feature_vector_flat[18] ),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0249_),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold498 (.A(\feature_vector_flat[48] ),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold499 (.A(_0279_),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold500 (.A(\leaf_value_flat[9] ),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold501 (.A(_0038_),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold502 (.A(\leaf_value_flat[29] ),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold503 (.A(_0058_),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold504 (.A(features_loaded),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold505 (.A(_1152_),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold506 (.A(_0021_),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold507 (.A(\leaf_value_flat[25] ),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold508 (.A(_0054_),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold509 (.A(\leaf_value_flat[24] ),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold510 (.A(_0053_),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold511 (.A(\node_feature_flat[6] ),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold512 (.A(_0211_),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold513 (.A(\feature_vector_flat[54] ),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold514 (.A(_0285_),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold515 (.A(\node_left_flat[8] ),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold516 (.A(_0129_),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold517 (.A(\node_threshold_flat[30] ),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0179_),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold519 (.A(\leaf_value_flat[13] ),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold520 (.A(_0042_),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold521 (.A(\u_model_loader.byte_idx_q[3] ),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold522 (.A(_0327_),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0026_),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold524 (.A(\leaf_value_flat[23] ),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold525 (.A(_0052_),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold526 (.A(\u_tree_core.depth_q[0] ),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0306_),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold528 (.A(\node_threshold_flat[29] ),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold529 (.A(_0178_),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold530 (.A(\node_threshold_flat[28] ),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold531 (.A(_0177_),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold532 (.A(\model_byte[0] ),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold533 (.A(\model_byte[1] ),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold534 (.A(\model_byte[2] ),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold535 (.A(\feature_byte[7] ),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold536 (.A(\model_byte[4] ),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold537 (.A(\feature_byte[6] ),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold538 (.A(\u_tree_core.state_q[0] ),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold539 (.A(_1123_),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold540 (.A(_0000_),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold541 (.A(\u_model_loader.byte_idx_q[2] ),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold542 (.A(_0326_),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold543 (.A(\feature_byte[4] ),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold544 (.A(\model_byte[5] ),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold545 (.A(\model_byte[6] ),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold546 (.A(run_cmd),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold547 (.A(_0001_),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold548 (.A(\model_byte[7] ),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold549 (.A(\feature_byte[5] ),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold550 (.A(\feature_byte[0] ),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold551 (.A(\feature_byte[2] ),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold552 (.A(\u_tree_core.current_node_q[2] ),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold553 (.A(_0310_),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold554 (.A(\feature_byte[3] ),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold555 (.A(\model_byte[3] ),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold556 (.A(\feature_byte[1] ),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold557 (.A(\u_model_loader.byte_idx_q[4] ),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold558 (.A(_0329_),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold559 (.A(_0027_),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold560 (.A(\u_feature_loader.feature_idx_q[2] ),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold561 (.A(\u_tree_core.current_node_q[1] ),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold562 (.A(_0309_),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold563 (.A(\u_tree_core.state_q[1] ),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold564 (.A(_0308_),
    .X(net1079));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_4 FILLER_0_175 ();
 sg13g2_fill_1 FILLER_0_179 ();
 sg13g2_fill_1 FILLER_0_185 ();
 sg13g2_fill_1 FILLER_0_194 ();
 sg13g2_fill_2 FILLER_0_200 ();
 sg13g2_fill_1 FILLER_0_202 ();
 sg13g2_fill_1 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_211 ();
 sg13g2_decap_8 FILLER_0_218 ();
 sg13g2_decap_8 FILLER_0_225 ();
 sg13g2_decap_8 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_239 ();
 sg13g2_decap_8 FILLER_0_246 ();
 sg13g2_decap_8 FILLER_0_253 ();
 sg13g2_fill_2 FILLER_0_260 ();
 sg13g2_fill_1 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_279 ();
 sg13g2_decap_8 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_293 ();
 sg13g2_decap_8 FILLER_0_300 ();
 sg13g2_decap_8 FILLER_0_307 ();
 sg13g2_decap_8 FILLER_0_314 ();
 sg13g2_decap_8 FILLER_0_321 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_4 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_fill_2 FILLER_1_140 ();
 sg13g2_fill_2 FILLER_1_169 ();
 sg13g2_fill_2 FILLER_1_225 ();
 sg13g2_fill_2 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_295 ();
 sg13g2_decap_8 FILLER_1_302 ();
 sg13g2_decap_8 FILLER_1_309 ();
 sg13g2_decap_8 FILLER_1_316 ();
 sg13g2_decap_8 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_330 ();
 sg13g2_decap_8 FILLER_1_337 ();
 sg13g2_decap_8 FILLER_1_344 ();
 sg13g2_decap_8 FILLER_1_351 ();
 sg13g2_decap_8 FILLER_1_358 ();
 sg13g2_decap_8 FILLER_1_365 ();
 sg13g2_decap_8 FILLER_1_372 ();
 sg13g2_decap_8 FILLER_1_379 ();
 sg13g2_decap_8 FILLER_1_386 ();
 sg13g2_decap_8 FILLER_1_393 ();
 sg13g2_decap_8 FILLER_1_400 ();
 sg13g2_fill_2 FILLER_1_407 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_153 ();
 sg13g2_fill_1 FILLER_2_160 ();
 sg13g2_decap_4 FILLER_2_226 ();
 sg13g2_fill_2 FILLER_2_230 ();
 sg13g2_fill_1 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_fill_2 FILLER_3_133 ();
 sg13g2_decap_4 FILLER_3_221 ();
 sg13g2_fill_2 FILLER_3_242 ();
 sg13g2_fill_1 FILLER_3_244 ();
 sg13g2_decap_8 FILLER_3_313 ();
 sg13g2_decap_8 FILLER_3_320 ();
 sg13g2_decap_8 FILLER_3_327 ();
 sg13g2_decap_8 FILLER_3_334 ();
 sg13g2_decap_8 FILLER_3_341 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_8 FILLER_3_355 ();
 sg13g2_decap_8 FILLER_3_362 ();
 sg13g2_decap_8 FILLER_3_369 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_4 FILLER_3_404 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_fill_2 FILLER_4_133 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_4 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_137 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_320 ();
 sg13g2_decap_8 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_334 ();
 sg13g2_decap_8 FILLER_5_341 ();
 sg13g2_decap_8 FILLER_5_348 ();
 sg13g2_decap_8 FILLER_5_355 ();
 sg13g2_decap_8 FILLER_5_362 ();
 sg13g2_decap_8 FILLER_5_369 ();
 sg13g2_decap_8 FILLER_5_376 ();
 sg13g2_decap_8 FILLER_5_383 ();
 sg13g2_decap_8 FILLER_5_390 ();
 sg13g2_decap_8 FILLER_5_397 ();
 sg13g2_decap_4 FILLER_5_404 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_fill_2 FILLER_6_176 ();
 sg13g2_fill_2 FILLER_6_201 ();
 sg13g2_fill_2 FILLER_6_210 ();
 sg13g2_fill_1 FILLER_6_212 ();
 sg13g2_decap_4 FILLER_6_243 ();
 sg13g2_fill_2 FILLER_6_247 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_4 FILLER_6_403 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_4 FILLER_7_140 ();
 sg13g2_fill_1 FILLER_7_148 ();
 sg13g2_decap_4 FILLER_7_153 ();
 sg13g2_decap_4 FILLER_7_193 ();
 sg13g2_fill_2 FILLER_7_197 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_decap_8 FILLER_7_215 ();
 sg13g2_decap_8 FILLER_7_222 ();
 sg13g2_decap_4 FILLER_7_229 ();
 sg13g2_fill_2 FILLER_7_233 ();
 sg13g2_decap_8 FILLER_7_239 ();
 sg13g2_decap_4 FILLER_7_246 ();
 sg13g2_fill_2 FILLER_7_250 ();
 sg13g2_fill_2 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_330 ();
 sg13g2_decap_8 FILLER_7_337 ();
 sg13g2_decap_8 FILLER_7_344 ();
 sg13g2_decap_8 FILLER_7_351 ();
 sg13g2_decap_8 FILLER_7_358 ();
 sg13g2_decap_8 FILLER_7_365 ();
 sg13g2_decap_8 FILLER_7_372 ();
 sg13g2_decap_8 FILLER_7_379 ();
 sg13g2_decap_8 FILLER_7_386 ();
 sg13g2_decap_8 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_400 ();
 sg13g2_fill_2 FILLER_7_407 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_4 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_208 ();
 sg13g2_decap_4 FILLER_8_215 ();
 sg13g2_fill_1 FILLER_8_219 ();
 sg13g2_decap_4 FILLER_8_247 ();
 sg13g2_fill_2 FILLER_8_265 ();
 sg13g2_fill_1 FILLER_8_267 ();
 sg13g2_decap_8 FILLER_8_328 ();
 sg13g2_decap_8 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_342 ();
 sg13g2_decap_8 FILLER_8_349 ();
 sg13g2_decap_8 FILLER_8_356 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_4 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_149 ();
 sg13g2_fill_2 FILLER_9_244 ();
 sg13g2_fill_1 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_331 ();
 sg13g2_decap_8 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_345 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_decap_8 FILLER_9_359 ();
 sg13g2_decap_8 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_9_373 ();
 sg13g2_decap_8 FILLER_9_380 ();
 sg13g2_decap_8 FILLER_9_387 ();
 sg13g2_decap_8 FILLER_9_394 ();
 sg13g2_decap_8 FILLER_9_401 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_fill_2 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_128 ();
 sg13g2_fill_2 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_decap_8 FILLER_10_248 ();
 sg13g2_decap_4 FILLER_10_255 ();
 sg13g2_decap_4 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_269 ();
 sg13g2_decap_8 FILLER_10_328 ();
 sg13g2_decap_8 FILLER_10_335 ();
 sg13g2_decap_8 FILLER_10_342 ();
 sg13g2_decap_8 FILLER_10_349 ();
 sg13g2_decap_8 FILLER_10_356 ();
 sg13g2_decap_8 FILLER_10_363 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_fill_2 FILLER_11_184 ();
 sg13g2_fill_1 FILLER_11_186 ();
 sg13g2_fill_2 FILLER_11_211 ();
 sg13g2_fill_2 FILLER_11_223 ();
 sg13g2_fill_1 FILLER_11_225 ();
 sg13g2_fill_2 FILLER_11_244 ();
 sg13g2_fill_1 FILLER_11_288 ();
 sg13g2_fill_2 FILLER_11_306 ();
 sg13g2_fill_1 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_fill_2 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_144 ();
 sg13g2_fill_1 FILLER_12_158 ();
 sg13g2_fill_1 FILLER_12_172 ();
 sg13g2_fill_2 FILLER_12_192 ();
 sg13g2_decap_8 FILLER_12_206 ();
 sg13g2_fill_2 FILLER_12_213 ();
 sg13g2_decap_4 FILLER_12_219 ();
 sg13g2_decap_4 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_328 ();
 sg13g2_decap_8 FILLER_12_335 ();
 sg13g2_decap_8 FILLER_12_342 ();
 sg13g2_decap_8 FILLER_12_349 ();
 sg13g2_decap_8 FILLER_12_356 ();
 sg13g2_decap_8 FILLER_12_363 ();
 sg13g2_decap_8 FILLER_12_370 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_fill_2 FILLER_13_133 ();
 sg13g2_fill_1 FILLER_13_135 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_fill_2 FILLER_13_147 ();
 sg13g2_fill_1 FILLER_13_176 ();
 sg13g2_decap_8 FILLER_13_205 ();
 sg13g2_decap_8 FILLER_13_212 ();
 sg13g2_decap_8 FILLER_13_219 ();
 sg13g2_decap_8 FILLER_13_226 ();
 sg13g2_decap_8 FILLER_13_233 ();
 sg13g2_decap_4 FILLER_13_240 ();
 sg13g2_fill_1 FILLER_13_244 ();
 sg13g2_fill_2 FILLER_13_262 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_fill_2 FILLER_14_133 ();
 sg13g2_fill_1 FILLER_14_135 ();
 sg13g2_fill_2 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_194 ();
 sg13g2_fill_1 FILLER_14_214 ();
 sg13g2_decap_4 FILLER_14_252 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_265 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_fill_2 FILLER_14_279 ();
 sg13g2_fill_1 FILLER_14_281 ();
 sg13g2_fill_1 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_4 FILLER_15_105 ();
 sg13g2_fill_2 FILLER_15_109 ();
 sg13g2_fill_1 FILLER_15_138 ();
 sg13g2_decap_8 FILLER_15_159 ();
 sg13g2_decap_4 FILLER_15_166 ();
 sg13g2_fill_2 FILLER_15_170 ();
 sg13g2_fill_1 FILLER_15_178 ();
 sg13g2_decap_4 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_4 FILLER_15_200 ();
 sg13g2_fill_1 FILLER_15_204 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_2 FILLER_15_262 ();
 sg13g2_fill_1 FILLER_15_264 ();
 sg13g2_fill_1 FILLER_15_271 ();
 sg13g2_fill_2 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_fill_2 FILLER_16_152 ();
 sg13g2_fill_2 FILLER_16_166 ();
 sg13g2_fill_1 FILLER_16_168 ();
 sg13g2_fill_2 FILLER_16_173 ();
 sg13g2_fill_1 FILLER_16_175 ();
 sg13g2_fill_2 FILLER_16_214 ();
 sg13g2_fill_2 FILLER_16_228 ();
 sg13g2_decap_4 FILLER_16_239 ();
 sg13g2_fill_1 FILLER_16_256 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_4 FILLER_17_105 ();
 sg13g2_decap_4 FILLER_17_215 ();
 sg13g2_fill_1 FILLER_17_219 ();
 sg13g2_decap_4 FILLER_17_224 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_234 ();
 sg13g2_fill_1 FILLER_17_266 ();
 sg13g2_fill_1 FILLER_17_293 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_1 FILLER_18_163 ();
 sg13g2_decap_4 FILLER_18_209 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_decap_4 FILLER_18_219 ();
 sg13g2_fill_2 FILLER_18_223 ();
 sg13g2_decap_4 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_242 ();
 sg13g2_decap_4 FILLER_18_257 ();
 sg13g2_decap_4 FILLER_18_271 ();
 sg13g2_decap_4 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_324 ();
 sg13g2_decap_8 FILLER_18_331 ();
 sg13g2_decap_8 FILLER_18_338 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_119 ();
 sg13g2_fill_2 FILLER_19_123 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_271 ();
 sg13g2_fill_1 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_324 ();
 sg13g2_decap_8 FILLER_19_331 ();
 sg13g2_decap_8 FILLER_19_338 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_decap_8 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_4 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_decap_4 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_1 FILLER_20_219 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_fill_1 FILLER_20_297 ();
 sg13g2_decap_8 FILLER_20_329 ();
 sg13g2_decap_8 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_decap_8 FILLER_20_350 ();
 sg13g2_decap_8 FILLER_20_357 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_4 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_102 ();
 sg13g2_fill_2 FILLER_21_223 ();
 sg13g2_fill_2 FILLER_21_235 ();
 sg13g2_fill_2 FILLER_21_241 ();
 sg13g2_fill_2 FILLER_21_272 ();
 sg13g2_fill_1 FILLER_21_274 ();
 sg13g2_fill_2 FILLER_21_290 ();
 sg13g2_fill_1 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_4 FILLER_22_63 ();
 sg13g2_fill_1 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_76 ();
 sg13g2_decap_8 FILLER_22_83 ();
 sg13g2_decap_8 FILLER_22_90 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_decap_4 FILLER_22_158 ();
 sg13g2_fill_2 FILLER_22_173 ();
 sg13g2_fill_2 FILLER_22_181 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_decap_4 FILLER_22_266 ();
 sg13g2_fill_2 FILLER_22_270 ();
 sg13g2_fill_2 FILLER_22_292 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_4 FILLER_22_349 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_decap_8 FILLER_22_362 ();
 sg13g2_decap_8 FILLER_22_369 ();
 sg13g2_decap_8 FILLER_22_376 ();
 sg13g2_decap_8 FILLER_22_383 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_8 FILLER_22_397 ();
 sg13g2_decap_4 FILLER_22_404 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_21 ();
 sg13g2_fill_2 FILLER_23_25 ();
 sg13g2_fill_2 FILLER_23_54 ();
 sg13g2_fill_1 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_89 ();
 sg13g2_decap_8 FILLER_23_96 ();
 sg13g2_decap_4 FILLER_23_103 ();
 sg13g2_fill_1 FILLER_23_134 ();
 sg13g2_decap_4 FILLER_23_187 ();
 sg13g2_fill_2 FILLER_23_191 ();
 sg13g2_fill_2 FILLER_23_205 ();
 sg13g2_fill_1 FILLER_23_211 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_decap_4 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_270 ();
 sg13g2_decap_4 FILLER_23_322 ();
 sg13g2_fill_2 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_4 FILLER_23_403 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_4 FILLER_24_28 ();
 sg13g2_fill_2 FILLER_24_68 ();
 sg13g2_decap_8 FILLER_24_93 ();
 sg13g2_decap_8 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_107 ();
 sg13g2_decap_8 FILLER_24_155 ();
 sg13g2_fill_2 FILLER_24_162 ();
 sg13g2_fill_1 FILLER_24_164 ();
 sg13g2_decap_8 FILLER_24_189 ();
 sg13g2_decap_8 FILLER_24_196 ();
 sg13g2_decap_8 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_210 ();
 sg13g2_fill_2 FILLER_24_217 ();
 sg13g2_fill_1 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_fill_2 FILLER_24_295 ();
 sg13g2_fill_1 FILLER_24_297 ();
 sg13g2_decap_8 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_323 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_24_387 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_fill_2 FILLER_25_60 ();
 sg13g2_decap_4 FILLER_25_98 ();
 sg13g2_fill_1 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_155 ();
 sg13g2_fill_2 FILLER_25_162 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_decap_4 FILLER_25_221 ();
 sg13g2_decap_4 FILLER_25_234 ();
 sg13g2_fill_1 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_4 FILLER_25_273 ();
 sg13g2_fill_1 FILLER_25_277 ();
 sg13g2_fill_2 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_4 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_73 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_fill_2 FILLER_26_116 ();
 sg13g2_fill_2 FILLER_26_147 ();
 sg13g2_fill_2 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_211 ();
 sg13g2_decap_8 FILLER_26_218 ();
 sg13g2_fill_2 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_decap_4 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_decap_8 FILLER_26_304 ();
 sg13g2_decap_4 FILLER_26_311 ();
 sg13g2_fill_2 FILLER_26_315 ();
 sg13g2_fill_2 FILLER_26_348 ();
 sg13g2_fill_2 FILLER_26_359 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_393 ();
 sg13g2_decap_8 FILLER_26_400 ();
 sg13g2_fill_2 FILLER_26_407 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_18 ();
 sg13g2_fill_2 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_fill_2 FILLER_27_262 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_306 ();
 sg13g2_decap_4 FILLER_27_313 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_fill_1 FILLER_28_57 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_fill_1 FILLER_28_87 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_fill_1 FILLER_28_196 ();
 sg13g2_fill_2 FILLER_28_206 ();
 sg13g2_fill_1 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_241 ();
 sg13g2_decap_4 FILLER_28_280 ();
 sg13g2_fill_2 FILLER_28_311 ();
 sg13g2_fill_1 FILLER_28_313 ();
 sg13g2_fill_1 FILLER_28_339 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_fill_2 FILLER_28_407 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_14 ();
 sg13g2_fill_2 FILLER_29_64 ();
 sg13g2_fill_1 FILLER_29_66 ();
 sg13g2_fill_2 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_178 ();
 sg13g2_fill_1 FILLER_29_188 ();
 sg13g2_fill_2 FILLER_29_202 ();
 sg13g2_fill_1 FILLER_29_204 ();
 sg13g2_fill_2 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_265 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_fill_2 FILLER_30_85 ();
 sg13g2_fill_1 FILLER_30_87 ();
 sg13g2_fill_1 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_138 ();
 sg13g2_fill_2 FILLER_30_160 ();
 sg13g2_fill_2 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_177 ();
 sg13g2_decap_4 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_226 ();
 sg13g2_fill_1 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_decap_4 FILLER_30_254 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_332 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_fill_1 FILLER_31_30 ();
 sg13g2_fill_1 FILLER_31_104 ();
 sg13g2_fill_2 FILLER_31_140 ();
 sg13g2_fill_1 FILLER_31_142 ();
 sg13g2_fill_1 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_fill_1 FILLER_31_168 ();
 sg13g2_decap_4 FILLER_31_175 ();
 sg13g2_fill_2 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_fill_1 FILLER_31_278 ();
 sg13g2_fill_2 FILLER_31_315 ();
 sg13g2_fill_1 FILLER_31_317 ();
 sg13g2_fill_2 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_fill_1 FILLER_31_389 ();
 sg13g2_fill_2 FILLER_31_407 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_4 FILLER_32_14 ();
 sg13g2_fill_2 FILLER_32_18 ();
 sg13g2_fill_2 FILLER_32_62 ();
 sg13g2_fill_2 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_146 ();
 sg13g2_decap_8 FILLER_32_153 ();
 sg13g2_decap_4 FILLER_32_160 ();
 sg13g2_fill_2 FILLER_32_174 ();
 sg13g2_fill_1 FILLER_32_182 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_decap_8 FILLER_32_215 ();
 sg13g2_decap_8 FILLER_32_222 ();
 sg13g2_decap_4 FILLER_32_234 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_257 ();
 sg13g2_fill_2 FILLER_32_305 ();
 sg13g2_fill_2 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_359 ();
 sg13g2_fill_2 FILLER_32_365 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_46 ();
 sg13g2_fill_2 FILLER_33_125 ();
 sg13g2_fill_2 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_172 ();
 sg13g2_fill_2 FILLER_33_190 ();
 sg13g2_fill_2 FILLER_33_201 ();
 sg13g2_fill_1 FILLER_33_203 ();
 sg13g2_fill_1 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_fill_2 FILLER_33_379 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_4 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_4 ();
 sg13g2_fill_2 FILLER_34_46 ();
 sg13g2_fill_1 FILLER_34_48 ();
 sg13g2_fill_2 FILLER_34_123 ();
 sg13g2_fill_1 FILLER_34_188 ();
 sg13g2_fill_1 FILLER_34_208 ();
 sg13g2_fill_1 FILLER_34_218 ();
 sg13g2_fill_2 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_fill_2 FILLER_34_303 ();
 sg13g2_fill_2 FILLER_34_328 ();
 sg13g2_fill_1 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_364 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_fill_2 FILLER_34_406 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_41 ();
 sg13g2_fill_2 FILLER_35_64 ();
 sg13g2_fill_1 FILLER_35_66 ();
 sg13g2_decap_4 FILLER_35_72 ();
 sg13g2_fill_2 FILLER_35_76 ();
 sg13g2_fill_2 FILLER_35_87 ();
 sg13g2_fill_1 FILLER_35_89 ();
 sg13g2_fill_2 FILLER_35_148 ();
 sg13g2_fill_1 FILLER_35_150 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_2 FILLER_35_264 ();
 sg13g2_fill_1 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_fill_1 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_299 ();
 sg13g2_decap_8 FILLER_35_306 ();
 sg13g2_decap_4 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_21 ();
 sg13g2_fill_1 FILLER_36_23 ();
 sg13g2_decap_8 FILLER_36_74 ();
 sg13g2_decap_4 FILLER_36_81 ();
 sg13g2_decap_8 FILLER_36_89 ();
 sg13g2_decap_8 FILLER_36_96 ();
 sg13g2_decap_4 FILLER_36_103 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_139 ();
 sg13g2_decap_4 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_2 FILLER_36_178 ();
 sg13g2_fill_1 FILLER_36_180 ();
 sg13g2_fill_2 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_2 FILLER_36_244 ();
 sg13g2_fill_1 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_decap_4 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_318 ();
 sg13g2_decap_4 FILLER_36_324 ();
 sg13g2_decap_8 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_349 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_fill_1 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_63 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_93 ();
 sg13g2_fill_1 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_167 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_decap_8 FILLER_37_181 ();
 sg13g2_fill_1 FILLER_37_197 ();
 sg13g2_decap_8 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_216 ();
 sg13g2_decap_8 FILLER_37_222 ();
 sg13g2_decap_8 FILLER_37_229 ();
 sg13g2_decap_4 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_265 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_fill_2 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_299 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_fill_2 FILLER_37_362 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_4 FILLER_38_28 ();
 sg13g2_fill_2 FILLER_38_68 ();
 sg13g2_fill_2 FILLER_38_97 ();
 sg13g2_fill_2 FILLER_38_138 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_4 FILLER_38_179 ();
 sg13g2_fill_1 FILLER_38_183 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_4 FILLER_38_207 ();
 sg13g2_fill_2 FILLER_38_211 ();
 sg13g2_decap_4 FILLER_38_247 ();
 sg13g2_fill_2 FILLER_38_262 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_fill_1 FILLER_38_296 ();
 sg13g2_fill_1 FILLER_38_310 ();
 sg13g2_fill_2 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_347 ();
 sg13g2_fill_2 FILLER_38_387 ();
 sg13g2_decap_8 FILLER_38_402 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_4 FILLER_39_14 ();
 sg13g2_fill_1 FILLER_39_18 ();
 sg13g2_fill_1 FILLER_39_110 ();
 sg13g2_fill_2 FILLER_39_140 ();
 sg13g2_fill_2 FILLER_39_227 ();
 sg13g2_fill_1 FILLER_39_244 ();
 sg13g2_fill_2 FILLER_39_274 ();
 sg13g2_fill_1 FILLER_39_276 ();
 sg13g2_fill_1 FILLER_39_288 ();
 sg13g2_decap_4 FILLER_39_300 ();
 sg13g2_fill_1 FILLER_39_316 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_324 ();
 sg13g2_fill_2 FILLER_39_335 ();
 sg13g2_fill_1 FILLER_39_337 ();
 sg13g2_fill_2 FILLER_39_379 ();
 sg13g2_fill_1 FILLER_39_381 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_fill_1 FILLER_40_21 ();
 sg13g2_fill_2 FILLER_40_79 ();
 sg13g2_fill_2 FILLER_40_86 ();
 sg13g2_fill_1 FILLER_40_100 ();
 sg13g2_fill_2 FILLER_40_121 ();
 sg13g2_fill_1 FILLER_40_153 ();
 sg13g2_fill_2 FILLER_40_195 ();
 sg13g2_fill_1 FILLER_40_197 ();
 sg13g2_fill_2 FILLER_40_211 ();
 sg13g2_fill_1 FILLER_40_277 ();
 sg13g2_decap_4 FILLER_40_360 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_4 FILLER_41_62 ();
 sg13g2_decap_4 FILLER_41_75 ();
 sg13g2_fill_2 FILLER_41_83 ();
 sg13g2_fill_1 FILLER_41_90 ();
 sg13g2_fill_1 FILLER_41_117 ();
 sg13g2_fill_1 FILLER_41_138 ();
 sg13g2_fill_1 FILLER_41_180 ();
 sg13g2_fill_2 FILLER_41_211 ();
 sg13g2_fill_2 FILLER_41_258 ();
 sg13g2_fill_1 FILLER_41_273 ();
 sg13g2_fill_2 FILLER_41_342 ();
 sg13g2_decap_8 FILLER_41_349 ();
 sg13g2_decap_8 FILLER_41_356 ();
 sg13g2_fill_1 FILLER_41_363 ();
 sg13g2_fill_1 FILLER_41_390 ();
 sg13g2_decap_4 FILLER_41_404 ();
 sg13g2_fill_1 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_4 FILLER_42_35 ();
 sg13g2_fill_1 FILLER_42_44 ();
 sg13g2_fill_2 FILLER_42_72 ();
 sg13g2_fill_2 FILLER_42_110 ();
 sg13g2_fill_2 FILLER_42_140 ();
 sg13g2_decap_4 FILLER_42_169 ();
 sg13g2_fill_2 FILLER_42_205 ();
 sg13g2_fill_1 FILLER_42_207 ();
 sg13g2_fill_2 FILLER_42_211 ();
 sg13g2_fill_1 FILLER_42_213 ();
 sg13g2_fill_2 FILLER_42_227 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_fill_2 FILLER_42_263 ();
 sg13g2_fill_1 FILLER_42_265 ();
 sg13g2_fill_1 FILLER_42_271 ();
 sg13g2_fill_2 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_288 ();
 sg13g2_decap_4 FILLER_42_292 ();
 sg13g2_fill_2 FILLER_42_296 ();
 sg13g2_fill_2 FILLER_42_330 ();
 sg13g2_decap_4 FILLER_42_353 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_4 FILLER_43_28 ();
 sg13g2_fill_2 FILLER_43_32 ();
 sg13g2_decap_4 FILLER_43_44 ();
 sg13g2_decap_4 FILLER_43_57 ();
 sg13g2_fill_2 FILLER_43_61 ();
 sg13g2_fill_2 FILLER_43_153 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_decap_4 FILLER_43_190 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_fill_2 FILLER_43_235 ();
 sg13g2_fill_1 FILLER_43_355 ();
 sg13g2_decap_4 FILLER_43_404 ();
 sg13g2_fill_1 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_4 FILLER_44_14 ();
 sg13g2_fill_1 FILLER_44_18 ();
 sg13g2_fill_1 FILLER_44_51 ();
 sg13g2_fill_1 FILLER_44_65 ();
 sg13g2_fill_2 FILLER_44_82 ();
 sg13g2_fill_1 FILLER_44_84 ();
 sg13g2_decap_4 FILLER_44_162 ();
 sg13g2_fill_2 FILLER_44_175 ();
 sg13g2_fill_2 FILLER_44_205 ();
 sg13g2_decap_8 FILLER_44_220 ();
 sg13g2_fill_2 FILLER_44_266 ();
 sg13g2_fill_2 FILLER_44_295 ();
 sg13g2_fill_1 FILLER_44_297 ();
 sg13g2_fill_2 FILLER_44_316 ();
 sg13g2_fill_1 FILLER_44_318 ();
 sg13g2_fill_2 FILLER_44_328 ();
 sg13g2_fill_2 FILLER_44_333 ();
 sg13g2_fill_1 FILLER_44_335 ();
 sg13g2_fill_1 FILLER_44_381 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_4 FILLER_45_14 ();
 sg13g2_fill_2 FILLER_45_18 ();
 sg13g2_decap_4 FILLER_45_69 ();
 sg13g2_fill_1 FILLER_45_110 ();
 sg13g2_fill_2 FILLER_45_205 ();
 sg13g2_fill_2 FILLER_45_212 ();
 sg13g2_fill_1 FILLER_45_214 ();
 sg13g2_decap_8 FILLER_45_243 ();
 sg13g2_decap_8 FILLER_45_250 ();
 sg13g2_fill_2 FILLER_45_257 ();
 sg13g2_fill_1 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_291 ();
 sg13g2_decap_4 FILLER_45_298 ();
 sg13g2_decap_8 FILLER_45_311 ();
 sg13g2_fill_2 FILLER_45_322 ();
 sg13g2_fill_2 FILLER_45_333 ();
 sg13g2_fill_1 FILLER_45_335 ();
 sg13g2_fill_2 FILLER_45_340 ();
 sg13g2_decap_4 FILLER_45_346 ();
 sg13g2_fill_2 FILLER_45_365 ();
 sg13g2_fill_2 FILLER_45_386 ();
 sg13g2_fill_1 FILLER_45_388 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_7 ();
 sg13g2_fill_1 FILLER_46_11 ();
 sg13g2_decap_4 FILLER_46_39 ();
 sg13g2_fill_1 FILLER_46_71 ();
 sg13g2_fill_2 FILLER_46_92 ();
 sg13g2_fill_1 FILLER_46_94 ();
 sg13g2_fill_1 FILLER_46_132 ();
 sg13g2_fill_1 FILLER_46_141 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_fill_1 FILLER_46_223 ();
 sg13g2_decap_8 FILLER_46_237 ();
 sg13g2_decap_8 FILLER_46_244 ();
 sg13g2_fill_1 FILLER_46_251 ();
 sg13g2_fill_2 FILLER_46_278 ();
 sg13g2_fill_2 FILLER_46_339 ();
 sg13g2_fill_1 FILLER_46_341 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_fill_2 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_16 ();
 sg13g2_fill_1 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_53 ();
 sg13g2_fill_1 FILLER_47_64 ();
 sg13g2_fill_1 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_152 ();
 sg13g2_fill_1 FILLER_47_154 ();
 sg13g2_fill_2 FILLER_47_168 ();
 sg13g2_fill_2 FILLER_47_176 ();
 sg13g2_fill_1 FILLER_47_178 ();
 sg13g2_decap_8 FILLER_47_185 ();
 sg13g2_decap_8 FILLER_47_192 ();
 sg13g2_decap_4 FILLER_47_199 ();
 sg13g2_decap_4 FILLER_47_216 ();
 sg13g2_decap_4 FILLER_47_224 ();
 sg13g2_fill_1 FILLER_47_228 ();
 sg13g2_decap_4 FILLER_47_265 ();
 sg13g2_decap_4 FILLER_47_276 ();
 sg13g2_fill_2 FILLER_47_280 ();
 sg13g2_fill_2 FILLER_47_345 ();
 sg13g2_fill_1 FILLER_47_347 ();
 sg13g2_fill_2 FILLER_47_361 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_fill_2 FILLER_48_46 ();
 sg13g2_fill_2 FILLER_48_74 ();
 sg13g2_fill_1 FILLER_48_89 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_decap_8 FILLER_48_151 ();
 sg13g2_fill_2 FILLER_48_158 ();
 sg13g2_fill_1 FILLER_48_183 ();
 sg13g2_fill_2 FILLER_48_197 ();
 sg13g2_fill_1 FILLER_48_199 ();
 sg13g2_decap_4 FILLER_48_213 ();
 sg13g2_fill_2 FILLER_48_231 ();
 sg13g2_fill_1 FILLER_48_233 ();
 sg13g2_fill_2 FILLER_48_278 ();
 sg13g2_fill_1 FILLER_48_280 ();
 sg13g2_fill_1 FILLER_48_284 ();
 sg13g2_fill_1 FILLER_48_298 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_fill_1 FILLER_48_368 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_4 FILLER_49_14 ();
 sg13g2_fill_2 FILLER_49_18 ();
 sg13g2_fill_2 FILLER_49_47 ();
 sg13g2_fill_1 FILLER_49_49 ();
 sg13g2_decap_4 FILLER_49_68 ();
 sg13g2_fill_1 FILLER_49_102 ();
 sg13g2_fill_1 FILLER_49_143 ();
 sg13g2_decap_8 FILLER_49_149 ();
 sg13g2_decap_8 FILLER_49_156 ();
 sg13g2_fill_1 FILLER_49_163 ();
 sg13g2_fill_1 FILLER_49_204 ();
 sg13g2_fill_2 FILLER_49_253 ();
 sg13g2_fill_2 FILLER_49_310 ();
 sg13g2_fill_1 FILLER_49_312 ();
 sg13g2_fill_2 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_328 ();
 sg13g2_fill_1 FILLER_49_381 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_fill_2 FILLER_50_28 ();
 sg13g2_fill_2 FILLER_50_39 ();
 sg13g2_fill_1 FILLER_50_41 ();
 sg13g2_fill_2 FILLER_50_56 ();
 sg13g2_fill_1 FILLER_50_58 ();
 sg13g2_fill_1 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_4 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_120 ();
 sg13g2_fill_2 FILLER_50_131 ();
 sg13g2_fill_1 FILLER_50_133 ();
 sg13g2_fill_2 FILLER_50_175 ();
 sg13g2_fill_1 FILLER_50_233 ();
 sg13g2_fill_1 FILLER_50_286 ();
 sg13g2_decap_4 FILLER_50_296 ();
 sg13g2_fill_2 FILLER_50_336 ();
 sg13g2_fill_2 FILLER_50_362 ();
 sg13g2_fill_1 FILLER_50_364 ();
 sg13g2_fill_2 FILLER_50_370 ();
 sg13g2_fill_2 FILLER_50_390 ();
 sg13g2_fill_1 FILLER_50_392 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_fill_2 FILLER_51_35 ();
 sg13g2_fill_1 FILLER_51_37 ();
 sg13g2_decap_4 FILLER_51_43 ();
 sg13g2_fill_2 FILLER_51_47 ();
 sg13g2_fill_2 FILLER_51_89 ();
 sg13g2_fill_1 FILLER_51_91 ();
 sg13g2_fill_2 FILLER_51_119 ();
 sg13g2_fill_1 FILLER_51_121 ();
 sg13g2_decap_8 FILLER_51_135 ();
 sg13g2_fill_1 FILLER_51_142 ();
 sg13g2_fill_2 FILLER_51_188 ();
 sg13g2_fill_1 FILLER_51_190 ();
 sg13g2_fill_2 FILLER_51_197 ();
 sg13g2_decap_8 FILLER_51_222 ();
 sg13g2_decap_8 FILLER_51_229 ();
 sg13g2_decap_8 FILLER_51_236 ();
 sg13g2_fill_1 FILLER_51_243 ();
 sg13g2_fill_2 FILLER_51_247 ();
 sg13g2_fill_1 FILLER_51_249 ();
 sg13g2_fill_1 FILLER_51_255 ();
 sg13g2_fill_1 FILLER_51_270 ();
 sg13g2_decap_8 FILLER_51_284 ();
 sg13g2_fill_1 FILLER_51_291 ();
 sg13g2_decap_8 FILLER_51_296 ();
 sg13g2_decap_4 FILLER_51_303 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_fill_2 FILLER_51_368 ();
 sg13g2_fill_2 FILLER_51_406 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_4 FILLER_52_14 ();
 sg13g2_fill_2 FILLER_52_18 ();
 sg13g2_fill_2 FILLER_52_24 ();
 sg13g2_decap_4 FILLER_52_40 ();
 sg13g2_fill_1 FILLER_52_84 ();
 sg13g2_fill_1 FILLER_52_94 ();
 sg13g2_decap_8 FILLER_52_131 ();
 sg13g2_fill_2 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_158 ();
 sg13g2_fill_1 FILLER_52_160 ();
 sg13g2_decap_8 FILLER_52_227 ();
 sg13g2_fill_2 FILLER_52_234 ();
 sg13g2_fill_1 FILLER_52_236 ();
 sg13g2_decap_4 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_277 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_fill_1 FILLER_53_14 ();
 sg13g2_fill_2 FILLER_53_47 ();
 sg13g2_fill_2 FILLER_53_200 ();
 sg13g2_fill_2 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_223 ();
 sg13g2_fill_2 FILLER_53_348 ();
 sg13g2_fill_1 FILLER_53_350 ();
 sg13g2_fill_1 FILLER_53_381 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_4 FILLER_54_14 ();
 sg13g2_fill_1 FILLER_54_68 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_fill_1 FILLER_54_107 ();
 sg13g2_decap_8 FILLER_54_121 ();
 sg13g2_fill_2 FILLER_54_128 ();
 sg13g2_fill_1 FILLER_54_130 ();
 sg13g2_fill_2 FILLER_54_186 ();
 sg13g2_fill_1 FILLER_54_188 ();
 sg13g2_decap_4 FILLER_54_277 ();
 sg13g2_fill_1 FILLER_54_344 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_fill_2 FILLER_54_380 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_fill_1 FILLER_55_14 ();
 sg13g2_fill_1 FILLER_55_64 ();
 sg13g2_fill_2 FILLER_55_87 ();
 sg13g2_fill_1 FILLER_55_112 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_fill_2 FILLER_55_198 ();
 sg13g2_decap_8 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_269 ();
 sg13g2_fill_2 FILLER_55_297 ();
 sg13g2_fill_1 FILLER_55_334 ();
 sg13g2_fill_1 FILLER_55_355 ();
 sg13g2_fill_1 FILLER_55_366 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_fill_1 FILLER_56_14 ();
 sg13g2_fill_1 FILLER_56_64 ();
 sg13g2_fill_2 FILLER_56_92 ();
 sg13g2_fill_1 FILLER_56_94 ();
 sg13g2_fill_2 FILLER_56_120 ();
 sg13g2_fill_2 FILLER_56_135 ();
 sg13g2_fill_1 FILLER_56_137 ();
 sg13g2_fill_2 FILLER_56_147 ();
 sg13g2_fill_1 FILLER_56_149 ();
 sg13g2_fill_2 FILLER_56_216 ();
 sg13g2_fill_2 FILLER_56_245 ();
 sg13g2_decap_8 FILLER_56_259 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_decap_4 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_275 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_fill_1 FILLER_56_290 ();
 sg13g2_fill_2 FILLER_56_308 ();
 sg13g2_fill_1 FILLER_56_310 ();
 sg13g2_fill_2 FILLER_56_329 ();
 sg13g2_fill_2 FILLER_56_370 ();
 sg13g2_fill_1 FILLER_56_372 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_fill_1 FILLER_57_21 ();
 sg13g2_fill_2 FILLER_57_76 ();
 sg13g2_fill_1 FILLER_57_104 ();
 sg13g2_fill_1 FILLER_57_110 ();
 sg13g2_fill_2 FILLER_57_140 ();
 sg13g2_fill_1 FILLER_57_142 ();
 sg13g2_fill_2 FILLER_57_167 ();
 sg13g2_fill_1 FILLER_57_173 ();
 sg13g2_fill_1 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_244 ();
 sg13g2_fill_2 FILLER_57_260 ();
 sg13g2_fill_1 FILLER_57_302 ();
 sg13g2_decap_4 FILLER_57_325 ();
 sg13g2_fill_1 FILLER_57_329 ();
 sg13g2_fill_2 FILLER_57_406 ();
 sg13g2_fill_1 FILLER_57_408 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_31 ();
 sg13g2_fill_2 FILLER_58_67 ();
 sg13g2_fill_2 FILLER_58_78 ();
 sg13g2_fill_1 FILLER_58_80 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_8 FILLER_58_133 ();
 sg13g2_fill_2 FILLER_58_140 ();
 sg13g2_fill_1 FILLER_58_146 ();
 sg13g2_fill_2 FILLER_58_161 ();
 sg13g2_fill_1 FILLER_58_215 ();
 sg13g2_fill_2 FILLER_58_224 ();
 sg13g2_decap_8 FILLER_58_274 ();
 sg13g2_fill_2 FILLER_58_281 ();
 sg13g2_fill_2 FILLER_58_331 ();
 sg13g2_fill_2 FILLER_58_390 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_4 FILLER_59_21 ();
 sg13g2_fill_2 FILLER_59_93 ();
 sg13g2_decap_4 FILLER_59_105 ();
 sg13g2_fill_2 FILLER_59_109 ();
 sg13g2_fill_2 FILLER_59_154 ();
 sg13g2_fill_1 FILLER_59_188 ();
 sg13g2_fill_1 FILLER_59_243 ();
 sg13g2_fill_1 FILLER_59_262 ();
 sg13g2_decap_4 FILLER_59_272 ();
 sg13g2_fill_2 FILLER_59_276 ();
 sg13g2_fill_2 FILLER_59_319 ();
 sg13g2_fill_1 FILLER_59_393 ();
 sg13g2_fill_2 FILLER_59_407 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_4 FILLER_60_35 ();
 sg13g2_fill_1 FILLER_60_76 ();
 sg13g2_decap_8 FILLER_60_100 ();
 sg13g2_decap_4 FILLER_60_107 ();
 sg13g2_fill_1 FILLER_60_161 ();
 sg13g2_decap_8 FILLER_60_175 ();
 sg13g2_fill_2 FILLER_60_206 ();
 sg13g2_fill_2 FILLER_60_259 ();
 sg13g2_fill_2 FILLER_60_268 ();
 sg13g2_fill_2 FILLER_60_355 ();
 sg13g2_fill_1 FILLER_60_357 ();
 sg13g2_fill_2 FILLER_60_371 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_4 FILLER_61_14 ();
 sg13g2_fill_2 FILLER_61_55 ();
 sg13g2_decap_8 FILLER_61_96 ();
 sg13g2_fill_1 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_180 ();
 sg13g2_fill_2 FILLER_61_200 ();
 sg13g2_fill_1 FILLER_61_208 ();
 sg13g2_fill_2 FILLER_61_226 ();
 sg13g2_fill_1 FILLER_61_228 ();
 sg13g2_fill_1 FILLER_61_251 ();
 sg13g2_fill_1 FILLER_61_279 ();
 sg13g2_fill_2 FILLER_61_322 ();
 sg13g2_fill_2 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_365 ();
 sg13g2_fill_1 FILLER_61_381 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_4 FILLER_62_7 ();
 sg13g2_fill_2 FILLER_62_11 ();
 sg13g2_fill_2 FILLER_62_40 ();
 sg13g2_fill_1 FILLER_62_137 ();
 sg13g2_fill_2 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_242 ();
 sg13g2_fill_1 FILLER_62_252 ();
 sg13g2_fill_1 FILLER_62_272 ();
 sg13g2_fill_1 FILLER_62_282 ();
 sg13g2_fill_2 FILLER_62_288 ();
 sg13g2_fill_1 FILLER_62_290 ();
 sg13g2_fill_2 FILLER_62_324 ();
 sg13g2_fill_2 FILLER_62_339 ();
 sg13g2_fill_1 FILLER_62_341 ();
 sg13g2_fill_2 FILLER_62_373 ();
 sg13g2_fill_1 FILLER_62_375 ();
 sg13g2_fill_1 FILLER_62_381 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_4 ();
 sg13g2_fill_2 FILLER_63_125 ();
 sg13g2_fill_1 FILLER_63_127 ();
 sg13g2_decap_8 FILLER_63_145 ();
 sg13g2_fill_2 FILLER_63_152 ();
 sg13g2_fill_1 FILLER_63_154 ();
 sg13g2_fill_2 FILLER_63_159 ();
 sg13g2_fill_2 FILLER_63_188 ();
 sg13g2_fill_1 FILLER_63_190 ();
 sg13g2_fill_1 FILLER_63_217 ();
 sg13g2_fill_1 FILLER_63_230 ();
 sg13g2_decap_4 FILLER_63_296 ();
 sg13g2_decap_8 FILLER_63_309 ();
 sg13g2_decap_8 FILLER_63_316 ();
 sg13g2_fill_2 FILLER_63_323 ();
 sg13g2_fill_1 FILLER_63_325 ();
 sg13g2_fill_2 FILLER_63_378 ();
 sg13g2_fill_2 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_7 ();
 sg13g2_fill_2 FILLER_64_47 ();
 sg13g2_fill_1 FILLER_64_86 ();
 sg13g2_fill_2 FILLER_64_100 ();
 sg13g2_fill_1 FILLER_64_102 ();
 sg13g2_decap_8 FILLER_64_148 ();
 sg13g2_decap_4 FILLER_64_155 ();
 sg13g2_fill_2 FILLER_64_159 ();
 sg13g2_decap_8 FILLER_64_223 ();
 sg13g2_decap_8 FILLER_64_234 ();
 sg13g2_fill_2 FILLER_64_241 ();
 sg13g2_decap_4 FILLER_64_246 ();
 sg13g2_fill_1 FILLER_64_250 ();
 sg13g2_fill_1 FILLER_64_287 ();
 sg13g2_fill_1 FILLER_64_326 ();
 sg13g2_fill_2 FILLER_64_357 ();
 sg13g2_fill_2 FILLER_64_406 ();
 sg13g2_fill_1 FILLER_64_408 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_4 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_11 ();
 sg13g2_fill_1 FILLER_65_57 ();
 sg13g2_fill_2 FILLER_65_90 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_fill_2 FILLER_65_130 ();
 sg13g2_fill_2 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_162 ();
 sg13g2_decap_8 FILLER_65_169 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_fill_2 FILLER_65_242 ();
 sg13g2_fill_2 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_255 ();
 sg13g2_fill_2 FILLER_65_367 ();
 sg13g2_fill_1 FILLER_65_369 ();
 sg13g2_fill_2 FILLER_65_379 ();
 sg13g2_fill_1 FILLER_65_381 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_fill_1 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_47 ();
 sg13g2_fill_1 FILLER_66_62 ();
 sg13g2_fill_2 FILLER_66_99 ();
 sg13g2_decap_4 FILLER_66_173 ();
 sg13g2_decap_8 FILLER_66_258 ();
 sg13g2_decap_8 FILLER_66_269 ();
 sg13g2_decap_4 FILLER_66_285 ();
 sg13g2_fill_1 FILLER_66_349 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_4 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_18 ();
 sg13g2_fill_1 FILLER_67_24 ();
 sg13g2_fill_2 FILLER_67_43 ();
 sg13g2_fill_2 FILLER_67_55 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_decap_4 FILLER_67_85 ();
 sg13g2_fill_1 FILLER_67_124 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_fill_1 FILLER_67_174 ();
 sg13g2_fill_2 FILLER_67_184 ();
 sg13g2_fill_1 FILLER_67_190 ();
 sg13g2_decap_4 FILLER_67_261 ();
 sg13g2_fill_2 FILLER_67_265 ();
 sg13g2_fill_1 FILLER_67_335 ();
 sg13g2_fill_2 FILLER_67_357 ();
 sg13g2_fill_1 FILLER_67_359 ();
 sg13g2_fill_2 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_4 FILLER_68_7 ();
 sg13g2_fill_2 FILLER_68_11 ();
 sg13g2_decap_4 FILLER_68_36 ();
 sg13g2_fill_2 FILLER_68_45 ();
 sg13g2_fill_1 FILLER_68_83 ();
 sg13g2_fill_1 FILLER_68_179 ();
 sg13g2_fill_1 FILLER_68_230 ();
 sg13g2_fill_2 FILLER_68_240 ();
 sg13g2_fill_1 FILLER_68_242 ();
 sg13g2_fill_1 FILLER_68_329 ();
 sg13g2_fill_2 FILLER_68_351 ();
 sg13g2_fill_1 FILLER_68_353 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_4 FILLER_69_7 ();
 sg13g2_fill_2 FILLER_69_42 ();
 sg13g2_fill_2 FILLER_69_53 ();
 sg13g2_fill_1 FILLER_69_55 ();
 sg13g2_fill_2 FILLER_69_97 ();
 sg13g2_fill_2 FILLER_69_114 ();
 sg13g2_fill_1 FILLER_69_134 ();
 sg13g2_decap_8 FILLER_69_166 ();
 sg13g2_decap_4 FILLER_69_173 ();
 sg13g2_fill_1 FILLER_69_204 ();
 sg13g2_fill_2 FILLER_69_223 ();
 sg13g2_fill_2 FILLER_69_261 ();
 sg13g2_fill_1 FILLER_69_272 ();
 sg13g2_fill_2 FILLER_69_278 ();
 sg13g2_fill_2 FILLER_69_347 ();
 sg13g2_fill_1 FILLER_69_349 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_fill_1 FILLER_70_59 ();
 sg13g2_fill_2 FILLER_70_87 ();
 sg13g2_fill_2 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_135 ();
 sg13g2_fill_2 FILLER_70_162 ();
 sg13g2_decap_4 FILLER_70_169 ();
 sg13g2_fill_1 FILLER_70_177 ();
 sg13g2_fill_2 FILLER_70_186 ();
 sg13g2_fill_1 FILLER_70_188 ();
 sg13g2_decap_8 FILLER_70_272 ();
 sg13g2_decap_4 FILLER_70_279 ();
 sg13g2_fill_2 FILLER_70_283 ();
 sg13g2_fill_1 FILLER_70_302 ();
 sg13g2_fill_2 FILLER_70_316 ();
 sg13g2_fill_2 FILLER_70_323 ();
 sg13g2_fill_2 FILLER_70_334 ();
 sg13g2_fill_2 FILLER_70_356 ();
 sg13g2_decap_4 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_71 ();
 sg13g2_fill_1 FILLER_71_73 ();
 sg13g2_fill_2 FILLER_71_100 ();
 sg13g2_fill_1 FILLER_71_167 ();
 sg13g2_decap_8 FILLER_71_199 ();
 sg13g2_fill_1 FILLER_71_206 ();
 sg13g2_fill_2 FILLER_71_252 ();
 sg13g2_fill_1 FILLER_71_272 ();
 sg13g2_fill_1 FILLER_71_290 ();
 sg13g2_fill_2 FILLER_71_300 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_fill_2 FILLER_71_312 ();
 sg13g2_fill_1 FILLER_71_361 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_fill_1 FILLER_71_408 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_4 FILLER_72_7 ();
 sg13g2_fill_2 FILLER_72_11 ();
 sg13g2_fill_1 FILLER_72_17 ();
 sg13g2_fill_2 FILLER_72_45 ();
 sg13g2_fill_1 FILLER_72_83 ();
 sg13g2_fill_1 FILLER_72_94 ();
 sg13g2_fill_1 FILLER_72_142 ();
 sg13g2_fill_2 FILLER_72_206 ();
 sg13g2_fill_1 FILLER_72_208 ();
 sg13g2_decap_8 FILLER_72_218 ();
 sg13g2_fill_1 FILLER_72_225 ();
 sg13g2_fill_2 FILLER_72_274 ();
 sg13g2_fill_1 FILLER_72_276 ();
 sg13g2_decap_4 FILLER_72_282 ();
 sg13g2_fill_2 FILLER_72_335 ();
 sg13g2_fill_1 FILLER_72_346 ();
 sg13g2_fill_1 FILLER_72_381 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_fill_1 FILLER_73_56 ();
 sg13g2_fill_2 FILLER_73_71 ();
 sg13g2_fill_2 FILLER_73_118 ();
 sg13g2_fill_1 FILLER_73_120 ();
 sg13g2_fill_2 FILLER_73_171 ();
 sg13g2_fill_1 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_374 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_fill_2 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_9 ();
 sg13g2_fill_2 FILLER_74_37 ();
 sg13g2_fill_1 FILLER_74_39 ();
 sg13g2_fill_2 FILLER_74_55 ();
 sg13g2_fill_1 FILLER_74_57 ();
 sg13g2_fill_1 FILLER_74_95 ();
 sg13g2_fill_1 FILLER_74_115 ();
 sg13g2_fill_1 FILLER_74_137 ();
 sg13g2_decap_4 FILLER_74_214 ();
 sg13g2_fill_1 FILLER_74_342 ();
 sg13g2_fill_2 FILLER_74_389 ();
 sg13g2_decap_4 FILLER_75_0 ();
 sg13g2_fill_1 FILLER_75_4 ();
 sg13g2_fill_2 FILLER_75_28 ();
 sg13g2_fill_1 FILLER_75_30 ();
 sg13g2_fill_1 FILLER_75_71 ();
 sg13g2_fill_2 FILLER_75_85 ();
 sg13g2_fill_1 FILLER_75_92 ();
 sg13g2_decap_8 FILLER_75_155 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_173 ();
 sg13g2_decap_4 FILLER_75_180 ();
 sg13g2_fill_2 FILLER_75_184 ();
 sg13g2_fill_1 FILLER_75_222 ();
 sg13g2_decap_4 FILLER_75_236 ();
 sg13g2_decap_4 FILLER_75_262 ();
 sg13g2_decap_4 FILLER_75_279 ();
 sg13g2_fill_2 FILLER_75_296 ();
 sg13g2_fill_2 FILLER_75_311 ();
 sg13g2_fill_1 FILLER_75_313 ();
 sg13g2_fill_2 FILLER_75_345 ();
 sg13g2_fill_1 FILLER_76_0 ();
 sg13g2_fill_2 FILLER_76_33 ();
 sg13g2_fill_1 FILLER_76_35 ();
 sg13g2_fill_1 FILLER_76_107 ();
 sg13g2_fill_1 FILLER_76_148 ();
 sg13g2_fill_1 FILLER_76_172 ();
 sg13g2_fill_1 FILLER_76_176 ();
 sg13g2_fill_1 FILLER_76_181 ();
 sg13g2_fill_1 FILLER_76_196 ();
 sg13g2_decap_8 FILLER_76_206 ();
 sg13g2_decap_8 FILLER_76_213 ();
 sg13g2_decap_8 FILLER_76_220 ();
 sg13g2_decap_8 FILLER_76_227 ();
 sg13g2_decap_8 FILLER_76_234 ();
 sg13g2_decap_8 FILLER_76_241 ();
 sg13g2_decap_8 FILLER_76_248 ();
 sg13g2_fill_2 FILLER_76_255 ();
 sg13g2_fill_1 FILLER_76_257 ();
 sg13g2_decap_8 FILLER_76_261 ();
 sg13g2_fill_1 FILLER_76_367 ();
 sg13g2_fill_2 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_394 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_49 ();
 sg13g2_fill_1 FILLER_77_64 ();
 sg13g2_fill_1 FILLER_77_74 ();
 sg13g2_fill_2 FILLER_77_130 ();
 sg13g2_fill_2 FILLER_77_247 ();
 sg13g2_fill_1 FILLER_77_262 ();
 sg13g2_fill_2 FILLER_77_314 ();
 sg13g2_fill_1 FILLER_77_316 ();
 sg13g2_fill_1 FILLER_77_344 ();
 sg13g2_fill_1 FILLER_77_363 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_fill_2 FILLER_78_81 ();
 sg13g2_fill_1 FILLER_78_83 ();
 sg13g2_fill_2 FILLER_78_93 ();
 sg13g2_fill_1 FILLER_78_95 ();
 sg13g2_fill_2 FILLER_78_137 ();
 sg13g2_fill_1 FILLER_78_139 ();
 sg13g2_fill_2 FILLER_78_212 ();
 sg13g2_fill_1 FILLER_78_371 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_4 FILLER_79_14 ();
 sg13g2_fill_1 FILLER_79_59 ();
 sg13g2_fill_1 FILLER_79_92 ();
 sg13g2_fill_2 FILLER_79_195 ();
 sg13g2_fill_2 FILLER_79_296 ();
 sg13g2_fill_1 FILLER_79_311 ();
 sg13g2_fill_2 FILLER_79_317 ();
 sg13g2_fill_2 FILLER_79_383 ();
 sg13g2_fill_2 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_fill_1 FILLER_80_52 ();
 sg13g2_fill_2 FILLER_80_97 ();
 sg13g2_fill_2 FILLER_80_113 ();
 sg13g2_fill_2 FILLER_80_127 ();
 sg13g2_fill_1 FILLER_80_129 ();
 sg13g2_fill_2 FILLER_80_134 ();
 sg13g2_fill_1 FILLER_80_136 ();
 sg13g2_decap_8 FILLER_80_141 ();
 sg13g2_fill_2 FILLER_80_148 ();
 sg13g2_fill_1 FILLER_80_150 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_4 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_188 ();
 sg13g2_decap_4 FILLER_80_195 ();
 sg13g2_fill_2 FILLER_80_199 ();
 sg13g2_decap_8 FILLER_80_210 ();
 sg13g2_fill_2 FILLER_80_217 ();
 sg13g2_fill_1 FILLER_80_223 ();
 sg13g2_fill_2 FILLER_80_228 ();
 sg13g2_fill_2 FILLER_80_239 ();
 sg13g2_fill_2 FILLER_80_266 ();
 sg13g2_fill_1 FILLER_80_289 ();
 sg13g2_fill_2 FILLER_80_312 ();
 sg13g2_fill_1 FILLER_80_314 ();
 sg13g2_fill_1 FILLER_80_363 ();
 sg13g2_fill_1 FILLER_80_373 ();
 sg13g2_fill_2 FILLER_80_392 ();
 sg13g2_fill_1 FILLER_80_394 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net330;
 assign uio_oe[4] = net331;
 assign uio_oe[5] = net332;
 assign uio_oe[6] = net333;
 assign uio_oe[7] = net334;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
endmodule
