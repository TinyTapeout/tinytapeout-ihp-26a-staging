module tt_um_vga_example (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire clknet_0_clk;
 wire horz_dir;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \square_x_pos[0] ;
 wire \square_x_pos[1] ;
 wire \square_x_pos[2] ;
 wire \square_x_pos[3] ;
 wire \square_x_pos[4] ;
 wire \square_x_pos[5] ;
 wire \square_x_pos[6] ;
 wire \square_x_pos[7] ;
 wire \square_x_pos[8] ;
 wire \square_x_pos[9] ;
 wire \square_y_pos[0] ;
 wire \square_y_pos[1] ;
 wire \square_y_pos[2] ;
 wire \square_y_pos[3] ;
 wire \square_y_pos[4] ;
 wire \square_y_pos[5] ;
 wire \square_y_pos[6] ;
 wire \square_y_pos[7] ;
 wire \square_y_pos[8] ;
 wire \square_y_pos[9] ;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire vert_dir;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;

 sg13g2_inv_1 _427_ (.Y(_403_),
    .A(net8));
 sg13g2_inv_2 _428_ (.Y(_404_),
    .A(net7));
 sg13g2_inv_1 _429_ (.Y(_044_),
    .A(net4));
 sg13g2_inv_1 _430_ (.Y(_045_),
    .A(net3));
 sg13g2_inv_1 _431_ (.Y(_046_),
    .A(net75));
 sg13g2_inv_1 _432_ (.Y(_047_),
    .A(net74));
 sg13g2_inv_1 _433_ (.Y(_048_),
    .A(\square_y_pos[3] ));
 sg13g2_inv_1 _434_ (.Y(_049_),
    .A(net71));
 sg13g2_inv_2 _435_ (.Y(_050_),
    .A(\square_y_pos[6] ));
 sg13g2_inv_1 _436_ (.Y(_051_),
    .A(\square_y_pos[7] ));
 sg13g2_inv_1 _437_ (.Y(_052_),
    .A(\square_y_pos[8] ));
 sg13g2_inv_2 _438_ (.Y(_053_),
    .A(vert_dir));
 sg13g2_inv_2 _439_ (.Y(_054_),
    .A(\square_x_pos[2] ));
 sg13g2_inv_1 _440_ (.Y(_055_),
    .A(\square_x_pos[3] ));
 sg13g2_inv_2 _441_ (.Y(_056_),
    .A(\square_x_pos[4] ));
 sg13g2_inv_1 _442_ (.Y(_057_),
    .A(\square_x_pos[5] ));
 sg13g2_inv_2 _443_ (.Y(_058_),
    .A(\square_x_pos[6] ));
 sg13g2_inv_2 _444_ (.Y(_059_),
    .A(\square_x_pos[7] ));
 sg13g2_inv_1 _445_ (.Y(_060_),
    .A(\square_x_pos[8] ));
 sg13g2_inv_1 _446_ (.Y(_061_),
    .A(net78));
 sg13g2_inv_1 _447_ (.Y(_062_),
    .A(net90));
 sg13g2_inv_1 _448_ (.Y(_063_),
    .A(\hvsync_gen.vpos[7] ));
 sg13g2_inv_2 _449_ (.Y(_064_),
    .A(net62));
 sg13g2_inv_2 _450_ (.Y(_065_),
    .A(net56));
 sg13g2_inv_1 _451_ (.Y(_066_),
    .A(\hvsync_gen.hpos[4] ));
 sg13g2_nand2_1 _452_ (.Y(_067_),
    .A(net100),
    .B(\hvsync_gen.vpos[6] ));
 sg13g2_nand4_1 _453_ (.B(net100),
    .C(net62),
    .A(\hvsync_gen.vpos[5] ),
    .Y(_068_),
    .D(net105));
 sg13g2_nor2_1 _454_ (.A(net79),
    .B(net78),
    .Y(_069_));
 sg13g2_nor2_1 _455_ (.A(\hvsync_gen.vpos[4] ),
    .B(net88),
    .Y(_070_));
 sg13g2_nand4_1 _456_ (.B(_061_),
    .C(net52),
    .A(net79),
    .Y(_071_),
    .D(_070_));
 sg13g2_nor2_1 _457_ (.A(_068_),
    .B(net53),
    .Y(_001_));
 sg13g2_nor3_1 _458_ (.A(net56),
    .B(\hvsync_gen.hpos[4] ),
    .C(net96),
    .Y(_072_));
 sg13g2_and3_1 _459_ (.X(_073_),
    .A(net56),
    .B(net104),
    .C(net96));
 sg13g2_nand2_1 _460_ (.Y(_074_),
    .A(net82),
    .B(net80));
 sg13g2_nor4_1 _461_ (.A(net81),
    .B(_072_),
    .C(_073_),
    .D(_074_),
    .Y(_000_));
 sg13g2_or2_1 _462_ (.X(_075_),
    .B(net81),
    .A(net82));
 sg13g2_nand2_1 _463_ (.Y(_076_),
    .A(net80),
    .B(_075_));
 sg13g2_nand3b_1 _464_ (.B(_068_),
    .C(_076_),
    .Y(_077_),
    .A_N(net88));
 sg13g2_nand4_1 _465_ (.B(net78),
    .C(net90),
    .A(net79),
    .Y(_078_),
    .D(\hvsync_gen.vpos[8] ));
 sg13g2_o21ai_1 _466_ (.B1(net91),
    .Y(_079_),
    .A1(_067_),
    .A2(_078_));
 sg13g2_nor4_1 _467_ (.A(net90),
    .B(\hvsync_gen.vpos[7] ),
    .C(\hvsync_gen.vpos[6] ),
    .D(\hvsync_gen.vpos[8] ),
    .Y(_080_));
 sg13g2_a21oi_1 _468_ (.A1(_069_),
    .A2(_080_),
    .Y(_081_),
    .B1(net91));
 sg13g2_nor2_1 _469_ (.A(\hvsync_gen.vpos[5] ),
    .B(_081_),
    .Y(_082_));
 sg13g2_nor4_1 _470_ (.A(net83),
    .B(\hvsync_gen.hpos[1] ),
    .C(net80),
    .D(_075_),
    .Y(_083_));
 sg13g2_a21oi_1 _471_ (.A1(_072_),
    .A2(_083_),
    .Y(_084_),
    .B1(\hvsync_gen.hpos[3] ));
 sg13g2_nand4_1 _472_ (.B(\hvsync_gen.hpos[1] ),
    .C(net80),
    .A(net83),
    .Y(_085_),
    .D(_073_));
 sg13g2_a21oi_1 _473_ (.A1(\hvsync_gen.hpos[3] ),
    .A2(_085_),
    .Y(_086_),
    .B1(_084_));
 sg13g2_a21oi_1 _474_ (.A1(_079_),
    .A2(_082_),
    .Y(_087_),
    .B1(_086_));
 sg13g2_nor2_2 _475_ (.A(_077_),
    .B(_087_),
    .Y(uo_out[6]));
 sg13g2_and3_2 _476_ (.X(_088_),
    .A(net75),
    .B(net74),
    .C(\square_y_pos[3] ));
 sg13g2_nor3_2 _477_ (.A(net72),
    .B(net71),
    .C(_088_),
    .Y(_089_));
 sg13g2_nor2_1 _478_ (.A(_050_),
    .B(_089_),
    .Y(_090_));
 sg13g2_xnor2_1 _479_ (.Y(_091_),
    .A(\square_y_pos[6] ),
    .B(_089_));
 sg13g2_inv_1 _480_ (.Y(_092_),
    .A(_091_));
 sg13g2_xor2_1 _481_ (.B(_088_),
    .A(net73),
    .X(_093_));
 sg13g2_nand2_1 _482_ (.Y(_094_),
    .A(net90),
    .B(_093_));
 sg13g2_nand2b_1 _483_ (.Y(_095_),
    .B(\square_y_pos[0] ),
    .A_N(\hvsync_gen.vpos[0] ));
 sg13g2_nand2_1 _484_ (.Y(_096_),
    .A(net79),
    .B(_095_));
 sg13g2_nor2_1 _485_ (.A(net79),
    .B(_095_),
    .Y(_097_));
 sg13g2_xor2_1 _486_ (.B(net74),
    .A(net75),
    .X(_098_));
 sg13g2_xnor2_1 _487_ (.Y(_099_),
    .A(net75),
    .B(net74));
 sg13g2_a221oi_1 _488_ (.B2(_061_),
    .C1(_097_),
    .B1(_098_),
    .A1(_046_),
    .Y(_100_),
    .A2(_096_));
 sg13g2_a21oi_1 _489_ (.A1(net75),
    .A2(net74),
    .Y(_101_),
    .B1(\square_y_pos[3] ));
 sg13g2_nor2_1 _490_ (.A(_088_),
    .B(_101_),
    .Y(_102_));
 sg13g2_inv_1 _491_ (.Y(_103_),
    .A(_102_));
 sg13g2_a221oi_1 _492_ (.B2(net91),
    .C1(_100_),
    .B1(_103_),
    .A1(net78),
    .Y(_104_),
    .A2(_099_));
 sg13g2_nand2b_1 _493_ (.Y(_105_),
    .B(_102_),
    .A_N(net91));
 sg13g2_o21ai_1 _494_ (.B1(_105_),
    .Y(_106_),
    .A1(net90),
    .A2(_093_));
 sg13g2_o21ai_1 _495_ (.B1(_094_),
    .Y(_107_),
    .A1(_104_),
    .A2(_106_));
 sg13g2_o21ai_1 _496_ (.B1(net71),
    .Y(_108_),
    .A1(net72),
    .A2(_088_));
 sg13g2_nor2b_2 _497_ (.A(_089_),
    .B_N(_108_),
    .Y(_109_));
 sg13g2_o21ai_1 _498_ (.B1(_107_),
    .Y(_110_),
    .A1(net89),
    .A2(_109_));
 sg13g2_a22oi_1 _499_ (.Y(_111_),
    .B1(_109_),
    .B2(net89),
    .A2(_092_),
    .A1(\hvsync_gen.vpos[6] ));
 sg13g2_a22oi_1 _500_ (.Y(_112_),
    .B1(_110_),
    .B2(_111_),
    .A2(_091_),
    .A1(_064_));
 sg13g2_xnor2_1 _501_ (.Y(_113_),
    .A(\square_y_pos[7] ),
    .B(_090_));
 sg13g2_a21o_1 _502_ (.A2(_113_),
    .A1(\hvsync_gen.vpos[7] ),
    .B1(_112_),
    .X(_114_));
 sg13g2_nand3_1 _503_ (.B(\square_y_pos[8] ),
    .C(_090_),
    .A(\square_y_pos[7] ),
    .Y(_115_));
 sg13g2_a21o_1 _504_ (.A2(_090_),
    .A1(\square_y_pos[7] ),
    .B1(\square_y_pos[8] ),
    .X(_116_));
 sg13g2_nand2_1 _505_ (.Y(_117_),
    .A(_115_),
    .B(_116_));
 sg13g2_nor2_1 _506_ (.A(\hvsync_gen.vpos[7] ),
    .B(_113_),
    .Y(_118_));
 sg13g2_nand2b_1 _507_ (.Y(_119_),
    .B(_115_),
    .A_N(\square_y_pos[9] ));
 sg13g2_xor2_1 _508_ (.B(_115_),
    .A(\square_y_pos[9] ),
    .X(_120_));
 sg13g2_or2_1 _509_ (.X(_121_),
    .B(_120_),
    .A(net88));
 sg13g2_xor2_1 _510_ (.B(_117_),
    .A(\hvsync_gen.vpos[8] ),
    .X(_122_));
 sg13g2_a21oi_1 _511_ (.A1(net88),
    .A2(_120_),
    .Y(_123_),
    .B1(_118_));
 sg13g2_nand4_1 _512_ (.B(_121_),
    .C(_122_),
    .A(_114_),
    .Y(_124_),
    .D(_123_));
 sg13g2_a221oi_1 _513_ (.B2(net75),
    .C1(_097_),
    .B1(_096_),
    .A1(net74),
    .Y(_125_),
    .A2(_061_));
 sg13g2_a221oi_1 _514_ (.B2(_048_),
    .C1(_125_),
    .B1(net91),
    .A1(_047_),
    .Y(_126_),
    .A2(net78));
 sg13g2_nor2_1 _515_ (.A(_049_),
    .B(net89),
    .Y(_127_));
 sg13g2_nand2b_1 _516_ (.Y(_128_),
    .B(net90),
    .A_N(net72));
 sg13g2_nor2b_1 _517_ (.A(net90),
    .B_N(net73),
    .Y(_129_));
 sg13g2_o21ai_1 _518_ (.B1(_128_),
    .Y(_130_),
    .A1(_048_),
    .A2(net91));
 sg13g2_nor4_1 _519_ (.A(_126_),
    .B(_127_),
    .C(_129_),
    .D(_130_),
    .Y(_131_));
 sg13g2_a22oi_1 _520_ (.Y(_132_),
    .B1(\hvsync_gen.vpos[6] ),
    .B2(_050_),
    .A2(net89),
    .A1(_049_));
 sg13g2_o21ai_1 _521_ (.B1(_132_),
    .Y(_133_),
    .A1(_127_),
    .A2(_128_));
 sg13g2_a22oi_1 _522_ (.Y(_134_),
    .B1(_064_),
    .B2(\square_y_pos[6] ),
    .A2(_063_),
    .A1(\square_y_pos[7] ));
 sg13g2_o21ai_1 _523_ (.B1(_134_),
    .Y(_135_),
    .A1(_131_),
    .A2(_133_));
 sg13g2_o21ai_1 _524_ (.B1(_135_),
    .Y(_136_),
    .A1(\square_y_pos[7] ),
    .A2(_063_));
 sg13g2_nor2b_1 _525_ (.A(\square_y_pos[8] ),
    .B_N(\hvsync_gen.vpos[8] ),
    .Y(_137_));
 sg13g2_nand2b_1 _526_ (.Y(_138_),
    .B(\square_y_pos[9] ),
    .A_N(net88));
 sg13g2_o21ai_1 _527_ (.B1(_138_),
    .Y(_139_),
    .A1(_052_),
    .A2(\hvsync_gen.vpos[8] ));
 sg13g2_nor2_1 _528_ (.A(_137_),
    .B(_139_),
    .Y(_140_));
 sg13g2_nor2b_1 _529_ (.A(\square_y_pos[9] ),
    .B_N(net88),
    .Y(_141_));
 sg13g2_a221oi_1 _530_ (.B2(_136_),
    .C1(_141_),
    .B1(_140_),
    .A1(_137_),
    .Y(_142_),
    .A2(_138_));
 sg13g2_nand3_1 _531_ (.B(_117_),
    .C(_121_),
    .A(\hvsync_gen.vpos[8] ),
    .Y(_143_));
 sg13g2_nand2b_1 _532_ (.Y(_144_),
    .B(\square_x_pos[9] ),
    .A_N(net80));
 sg13g2_nand2b_1 _533_ (.Y(_145_),
    .B(_144_),
    .A_N(_077_));
 sg13g2_nand2_1 _534_ (.Y(_146_),
    .A(net76),
    .B(\square_x_pos[2] ));
 sg13g2_and3_2 _535_ (.X(_147_),
    .A(net76),
    .B(\square_x_pos[2] ),
    .C(\square_x_pos[3] ));
 sg13g2_nor3_1 _536_ (.A(\square_x_pos[4] ),
    .B(\square_x_pos[5] ),
    .C(_147_),
    .Y(_148_));
 sg13g2_nand2b_1 _537_ (.Y(_149_),
    .B(\square_x_pos[6] ),
    .A_N(_148_));
 sg13g2_nor2_1 _538_ (.A(_059_),
    .B(_149_),
    .Y(_150_));
 sg13g2_nand2_1 _539_ (.Y(_151_),
    .A(\square_x_pos[8] ),
    .B(_150_));
 sg13g2_nand2b_1 _540_ (.Y(_152_),
    .B(net80),
    .A_N(\square_x_pos[9] ));
 sg13g2_xnor2_1 _541_ (.Y(_153_),
    .A(\square_x_pos[8] ),
    .B(_150_));
 sg13g2_nand2_1 _542_ (.Y(_154_),
    .A(net81),
    .B(_153_));
 sg13g2_and2_1 _543_ (.A(net47),
    .B(net61),
    .X(_155_));
 sg13g2_xnor2_1 _544_ (.Y(_156_),
    .A(net76),
    .B(\square_x_pos[2] ));
 sg13g2_nor2_1 _545_ (.A(net83),
    .B(_156_),
    .Y(_157_));
 sg13g2_nor2_1 _546_ (.A(net47),
    .B(net61),
    .Y(_158_));
 sg13g2_nand2_1 _547_ (.Y(_159_),
    .A(net76),
    .B(\hvsync_gen.hpos[1] ));
 sg13g2_nand2b_1 _548_ (.Y(_160_),
    .B(\square_x_pos[0] ),
    .A_N(\hvsync_gen.hpos[0] ));
 sg13g2_o21ai_1 _549_ (.B1(_160_),
    .Y(_161_),
    .A1(net76),
    .A2(\hvsync_gen.hpos[1] ));
 sg13g2_a21o_1 _550_ (.A2(_161_),
    .A1(_159_),
    .B1(_157_),
    .X(_162_));
 sg13g2_xnor2_1 _551_ (.Y(_163_),
    .A(\square_x_pos[3] ),
    .B(_146_));
 sg13g2_xnor2_1 _552_ (.Y(_164_),
    .A(_055_),
    .B(_146_));
 sg13g2_a22oi_1 _553_ (.Y(_165_),
    .B1(_164_),
    .B2(\hvsync_gen.hpos[3] ),
    .A2(_156_),
    .A1(net83));
 sg13g2_nor2_1 _554_ (.A(\hvsync_gen.hpos[3] ),
    .B(_164_),
    .Y(_166_));
 sg13g2_xnor2_1 _555_ (.Y(_167_),
    .A(_056_),
    .B(_147_));
 sg13g2_inv_1 _556_ (.Y(_168_),
    .A(_167_));
 sg13g2_a221oi_1 _557_ (.B2(_066_),
    .C1(_166_),
    .B1(_168_),
    .A1(_162_),
    .Y(_169_),
    .A2(_165_));
 sg13g2_o21ai_1 _558_ (.B1(\square_x_pos[5] ),
    .Y(_170_),
    .A1(\square_x_pos[4] ),
    .A2(_147_));
 sg13g2_nand2b_1 _559_ (.Y(_171_),
    .B(_170_),
    .A_N(_148_));
 sg13g2_inv_1 _560_ (.Y(_172_),
    .A(_171_));
 sg13g2_a221oi_1 _561_ (.B2(\hvsync_gen.hpos[5] ),
    .C1(_169_),
    .B1(_172_),
    .A1(\hvsync_gen.hpos[4] ),
    .Y(_173_),
    .A2(_167_));
 sg13g2_xnor2_1 _562_ (.Y(_174_),
    .A(_058_),
    .B(_148_));
 sg13g2_nand2_1 _563_ (.Y(_175_),
    .A(_065_),
    .B(_171_));
 sg13g2_o21ai_1 _564_ (.B1(_175_),
    .Y(_176_),
    .A1(\hvsync_gen.hpos[6] ),
    .A2(_174_));
 sg13g2_xnor2_1 _565_ (.Y(_177_),
    .A(_059_),
    .B(_149_));
 sg13g2_a22oi_1 _566_ (.Y(_178_),
    .B1(_177_),
    .B2(net82),
    .A2(_174_),
    .A1(\hvsync_gen.hpos[6] ));
 sg13g2_o21ai_1 _567_ (.B1(_178_),
    .Y(_179_),
    .A1(_173_),
    .A2(_176_));
 sg13g2_or2_1 _568_ (.X(_180_),
    .B(_177_),
    .A(net82));
 sg13g2_o21ai_1 _569_ (.B1(_180_),
    .Y(_181_),
    .A1(net81),
    .A2(_153_));
 sg13g2_nand2b_1 _570_ (.Y(_182_),
    .B(_179_),
    .A_N(_181_));
 sg13g2_nand2_1 _571_ (.Y(_183_),
    .A(_144_),
    .B(_151_));
 sg13g2_a22oi_1 _572_ (.Y(_184_),
    .B1(_183_),
    .B2(_152_),
    .A2(_182_),
    .A1(_154_));
 sg13g2_nand2b_1 _573_ (.Y(_185_),
    .B(net76),
    .A_N(\hvsync_gen.hpos[1] ));
 sg13g2_nor2b_1 _574_ (.A(net76),
    .B_N(\hvsync_gen.hpos[1] ),
    .Y(_186_));
 sg13g2_a221oi_1 _575_ (.B2(_185_),
    .C1(_186_),
    .B1(_160_),
    .A1(_054_),
    .Y(_187_),
    .A2(\hvsync_gen.hpos[2] ));
 sg13g2_nand2b_1 _576_ (.Y(_188_),
    .B(\square_x_pos[3] ),
    .A_N(\hvsync_gen.hpos[3] ));
 sg13g2_o21ai_1 _577_ (.B1(_188_),
    .Y(_189_),
    .A1(_054_),
    .A2(\hvsync_gen.hpos[2] ));
 sg13g2_a22oi_1 _578_ (.Y(_190_),
    .B1(\hvsync_gen.hpos[4] ),
    .B2(_056_),
    .A2(\hvsync_gen.hpos[3] ),
    .A1(_055_));
 sg13g2_o21ai_1 _579_ (.B1(_190_),
    .Y(_191_),
    .A1(_187_),
    .A2(_189_));
 sg13g2_a22oi_1 _580_ (.Y(_192_),
    .B1(_066_),
    .B2(\square_x_pos[4] ),
    .A2(_065_),
    .A1(\square_x_pos[5] ));
 sg13g2_nor2_1 _581_ (.A(\square_x_pos[5] ),
    .B(_065_),
    .Y(_193_));
 sg13g2_a221oi_1 _582_ (.B2(_192_),
    .C1(_193_),
    .B1(_191_),
    .A1(_058_),
    .Y(_194_),
    .A2(\hvsync_gen.hpos[6] ));
 sg13g2_nand2b_1 _583_ (.Y(_195_),
    .B(\square_x_pos[7] ),
    .A_N(net82));
 sg13g2_o21ai_1 _584_ (.B1(_195_),
    .Y(_196_),
    .A1(_058_),
    .A2(\hvsync_gen.hpos[6] ));
 sg13g2_a22oi_1 _585_ (.Y(_197_),
    .B1(net81),
    .B2(_060_),
    .A2(net82),
    .A1(_059_));
 sg13g2_o21ai_1 _586_ (.B1(_197_),
    .Y(_198_),
    .A1(_194_),
    .A2(_196_));
 sg13g2_o21ai_1 _587_ (.B1(_152_),
    .Y(_199_),
    .A1(_060_),
    .A2(\hvsync_gen.hpos[8] ));
 sg13g2_nand2b_1 _588_ (.Y(_200_),
    .B(_198_),
    .A_N(_199_));
 sg13g2_o21ai_1 _589_ (.B1(_200_),
    .Y(_201_),
    .A1(_151_),
    .A2(_152_));
 sg13g2_nand2_1 _590_ (.Y(_202_),
    .A(_143_),
    .B(_201_));
 sg13g2_nor4_1 _591_ (.A(_142_),
    .B(_145_),
    .C(_184_),
    .D(_202_),
    .Y(_203_));
 sg13g2_a21o_2 _592_ (.A2(_203_),
    .A1(_124_),
    .B1(uo_out[6]),
    .X(uo_out[5]));
 sg13g2_and3_2 _593_ (.X(_204_),
    .A(net83),
    .B(net58),
    .C(_155_));
 sg13g2_nand2_2 _594_ (.Y(_205_),
    .A(net104),
    .B(_204_));
 sg13g2_inv_1 _595_ (.Y(_206_),
    .A(_205_));
 sg13g2_nand3b_1 _596_ (.B(\hvsync_gen.hpos[9] ),
    .C(net81),
    .Y(_207_),
    .A_N(\hvsync_gen.hpos[7] ));
 sg13g2_nor4_2 _597_ (.A(net56),
    .B(\hvsync_gen.hpos[6] ),
    .C(_205_),
    .Y(_208_),
    .D(_207_));
 sg13g2_nor2b_2 _598_ (.A(_208_),
    .B_N(net94),
    .Y(_209_));
 sg13g2_nand2b_2 _599_ (.Y(_210_),
    .B(net94),
    .A_N(_208_));
 sg13g2_nand2_1 _600_ (.Y(_211_),
    .A(net52),
    .B(net67));
 sg13g2_nand3_1 _601_ (.B(net79),
    .C(net78),
    .A(net55),
    .Y(_212_));
 sg13g2_nand4_1 _602_ (.B(net79),
    .C(net78),
    .A(net55),
    .Y(_213_),
    .D(net91));
 sg13g2_xor2_1 _603_ (.B(_212_),
    .A(net52),
    .X(_214_));
 sg13g2_nand4_1 _604_ (.B(net91),
    .C(\hvsync_gen.vpos[9] ),
    .A(net78),
    .Y(_215_),
    .D(_080_));
 sg13g2_nor4_1 _605_ (.A(\hvsync_gen.vpos[0] ),
    .B(net79),
    .C(net89),
    .D(_215_),
    .Y(_216_));
 sg13g2_nand3b_1 _606_ (.B(net57),
    .C(net94),
    .Y(_217_),
    .A_N(_216_));
 sg13g2_o21ai_1 _607_ (.B1(_211_),
    .Y(_002_),
    .A1(_214_),
    .A2(net66));
 sg13g2_nand2_1 _608_ (.Y(_218_),
    .A(net90),
    .B(net67));
 sg13g2_nor2_1 _609_ (.A(_062_),
    .B(_213_),
    .Y(_219_));
 sg13g2_xnor2_1 _610_ (.Y(_220_),
    .A(_062_),
    .B(_213_));
 sg13g2_o21ai_1 _611_ (.B1(_218_),
    .Y(_003_),
    .A1(net66),
    .A2(_220_));
 sg13g2_nand2_1 _612_ (.Y(_221_),
    .A(net89),
    .B(net67));
 sg13g2_nand2_1 _613_ (.Y(_222_),
    .A(net89),
    .B(_219_));
 sg13g2_inv_1 _614_ (.Y(_223_),
    .A(_222_));
 sg13g2_xnor2_1 _615_ (.Y(_224_),
    .A(net89),
    .B(_219_));
 sg13g2_o21ai_1 _616_ (.B1(_221_),
    .Y(_004_),
    .A1(net66),
    .A2(_224_));
 sg13g2_nand2_1 _617_ (.Y(_225_),
    .A(net62),
    .B(net67));
 sg13g2_xnor2_1 _618_ (.Y(_226_),
    .A(_064_),
    .B(_222_));
 sg13g2_o21ai_1 _619_ (.B1(_225_),
    .Y(_005_),
    .A1(net66),
    .A2(_226_));
 sg13g2_a21oi_1 _620_ (.A1(net62),
    .A2(_223_),
    .Y(_227_),
    .B1(net100));
 sg13g2_nor2_1 _621_ (.A(_067_),
    .B(_222_),
    .Y(_228_));
 sg13g2_nor3_1 _622_ (.A(net66),
    .B(_227_),
    .C(_228_),
    .Y(_229_));
 sg13g2_a21o_1 _623_ (.A2(net67),
    .A1(net100),
    .B1(_229_),
    .X(_006_));
 sg13g2_nor3_1 _624_ (.A(_062_),
    .B(_068_),
    .C(_213_),
    .Y(_230_));
 sg13g2_o21ai_1 _625_ (.B1(_210_),
    .Y(_231_),
    .A1(net66),
    .A2(_230_));
 sg13g2_nor2b_1 _626_ (.A(net66),
    .B_N(_228_),
    .Y(_232_));
 sg13g2_o21ai_1 _627_ (.B1(_231_),
    .Y(_233_),
    .A1(net105),
    .A2(_232_));
 sg13g2_inv_1 _628_ (.Y(_007_),
    .A(net106));
 sg13g2_nand2_1 _629_ (.Y(_234_),
    .A(net88),
    .B(_231_));
 sg13g2_nand2b_1 _630_ (.Y(_235_),
    .B(_230_),
    .A_N(net66));
 sg13g2_o21ai_1 _631_ (.B1(_234_),
    .Y(_008_),
    .A1(net88),
    .A2(_235_));
 sg13g2_nor3_1 _632_ (.A(_044_),
    .B(_088_),
    .C(_101_),
    .Y(_236_));
 sg13g2_o21ai_1 _633_ (.B1(_044_),
    .Y(_237_),
    .A1(_088_),
    .A2(_101_));
 sg13g2_nor2b_1 _634_ (.A(net75),
    .B_N(net2),
    .Y(_238_));
 sg13g2_and2_1 _635_ (.A(net1),
    .B(\square_y_pos[0] ),
    .X(_239_));
 sg13g2_nand2b_1 _636_ (.Y(_240_),
    .B(net75),
    .A_N(net2));
 sg13g2_a221oi_1 _637_ (.B2(_240_),
    .C1(_238_),
    .B1(_239_),
    .A1(net3),
    .Y(_241_),
    .A2(_098_));
 sg13g2_a21oi_1 _638_ (.A1(_045_),
    .A2(_099_),
    .Y(_242_),
    .B1(_241_));
 sg13g2_o21ai_1 _639_ (.B1(_237_),
    .Y(_243_),
    .A1(_236_),
    .A2(_242_));
 sg13g2_o21ai_1 _640_ (.B1(_109_),
    .Y(_244_),
    .A1(_093_),
    .A2(_243_));
 sg13g2_and2_1 _641_ (.A(\square_y_pos[7] ),
    .B(_091_),
    .X(_245_));
 sg13g2_and2_1 _642_ (.A(\square_y_pos[8] ),
    .B(_245_),
    .X(_246_));
 sg13g2_a21oi_1 _643_ (.A1(_244_),
    .A2(_246_),
    .Y(_247_),
    .B1(_119_));
 sg13g2_a21o_1 _644_ (.A2(_243_),
    .A1(_093_),
    .B1(_109_),
    .X(_248_));
 sg13g2_nand2_1 _645_ (.Y(_249_),
    .A(net4),
    .B(\square_y_pos[3] ));
 sg13g2_xor2_1 _646_ (.B(\square_y_pos[3] ),
    .A(net4),
    .X(_250_));
 sg13g2_nor2_1 _647_ (.A(_045_),
    .B(_047_),
    .Y(_251_));
 sg13g2_xor2_1 _648_ (.B(net74),
    .A(net3),
    .X(_252_));
 sg13g2_nand2b_1 _649_ (.Y(_253_),
    .B(_240_),
    .A_N(_238_));
 sg13g2_and2_1 _650_ (.A(net2),
    .B(\square_y_pos[1] ),
    .X(_254_));
 sg13g2_a21o_1 _651_ (.A2(_253_),
    .A1(_239_),
    .B1(_254_),
    .X(_255_));
 sg13g2_a21oi_1 _652_ (.A1(_252_),
    .A2(_255_),
    .Y(_256_),
    .B1(_251_));
 sg13g2_nand2b_1 _653_ (.Y(_257_),
    .B(_250_),
    .A_N(_256_));
 sg13g2_xnor2_1 _654_ (.Y(_258_),
    .A(_250_),
    .B(_256_));
 sg13g2_xor2_1 _655_ (.B(_255_),
    .A(_252_),
    .X(_259_));
 sg13g2_nor2b_1 _656_ (.A(\square_y_pos[0] ),
    .B_N(net1),
    .Y(_260_));
 sg13g2_xor2_1 _657_ (.B(\square_y_pos[0] ),
    .A(net1),
    .X(_261_));
 sg13g2_nor2_1 _658_ (.A(\square_y_pos[9] ),
    .B(_261_),
    .Y(_262_));
 sg13g2_xor2_1 _659_ (.B(_253_),
    .A(_239_),
    .X(_263_));
 sg13g2_and4_1 _660_ (.A(_245_),
    .B(_259_),
    .C(_262_),
    .D(_263_),
    .X(_264_));
 sg13g2_and4_1 _661_ (.A(_244_),
    .B(_248_),
    .C(_258_),
    .D(_264_),
    .X(_265_));
 sg13g2_nor2_1 _662_ (.A(vert_dir),
    .B(_258_),
    .Y(_266_));
 sg13g2_nor3_2 _663_ (.A(vert_dir),
    .B(_247_),
    .C(_265_),
    .Y(_267_));
 sg13g2_nor4_1 _664_ (.A(net2),
    .B(net1),
    .C(net4),
    .D(net3),
    .Y(_268_));
 sg13g2_nand2b_1 _665_ (.Y(_269_),
    .B(_267_),
    .A_N(_268_));
 sg13g2_a21o_1 _666_ (.A2(_260_),
    .A1(_240_),
    .B1(_238_),
    .X(_270_));
 sg13g2_or2_1 _667_ (.X(_271_),
    .B(_270_),
    .A(_252_));
 sg13g2_nand2_1 _668_ (.Y(_272_),
    .A(_045_),
    .B(\square_y_pos[2] ));
 sg13g2_a21oi_1 _669_ (.A1(_271_),
    .A2(_272_),
    .Y(_273_),
    .B1(_250_));
 sg13g2_a21oi_1 _670_ (.A1(_044_),
    .A2(\square_y_pos[3] ),
    .Y(_274_),
    .B1(_273_));
 sg13g2_nor3_1 _671_ (.A(net72),
    .B(net71),
    .C(\square_y_pos[6] ),
    .Y(_275_));
 sg13g2_nand3_1 _672_ (.B(_274_),
    .C(_275_),
    .A(_051_),
    .Y(_276_));
 sg13g2_nor3_1 _673_ (.A(\square_y_pos[8] ),
    .B(\square_y_pos[9] ),
    .C(_276_),
    .Y(_277_));
 sg13g2_o21ai_1 _674_ (.B1(_269_),
    .Y(_009_),
    .A1(_053_),
    .A2(_277_));
 sg13g2_nor2_1 _675_ (.A(net47),
    .B(_210_),
    .Y(_010_));
 sg13g2_nor3_1 _676_ (.A(_155_),
    .B(_158_),
    .C(_210_),
    .Y(_011_));
 sg13g2_o21ai_1 _677_ (.B1(net67),
    .Y(_278_),
    .A1(net83),
    .A2(_155_));
 sg13g2_a21oi_1 _678_ (.A1(net83),
    .A2(_155_),
    .Y(_012_),
    .B1(_278_));
 sg13g2_a21oi_1 _679_ (.A1(net83),
    .A2(_155_),
    .Y(_279_),
    .B1(net58));
 sg13g2_nor3_1 _680_ (.A(_204_),
    .B(_210_),
    .C(net59),
    .Y(_013_));
 sg13g2_o21ai_1 _681_ (.B1(net93),
    .Y(_280_),
    .A1(net104),
    .A2(_204_));
 sg13g2_nor2_1 _682_ (.A(_206_),
    .B(_280_),
    .Y(_014_));
 sg13g2_xnor2_1 _683_ (.Y(_281_),
    .A(_065_),
    .B(_205_));
 sg13g2_nor2_1 _684_ (.A(_210_),
    .B(_281_),
    .Y(_015_));
 sg13g2_and2_1 _685_ (.A(_073_),
    .B(_204_),
    .X(_282_));
 sg13g2_a21oi_1 _686_ (.A1(net56),
    .A2(_206_),
    .Y(_283_),
    .B1(net96));
 sg13g2_nor3_1 _687_ (.A(_210_),
    .B(_282_),
    .C(net97),
    .Y(_016_));
 sg13g2_and2_1 _688_ (.A(net82),
    .B(_282_),
    .X(_284_));
 sg13g2_nor2_1 _689_ (.A(net82),
    .B(_282_),
    .Y(_285_));
 sg13g2_nor3_1 _690_ (.A(_210_),
    .B(_284_),
    .C(_285_),
    .Y(_017_));
 sg13g2_and2_1 _691_ (.A(net81),
    .B(_284_),
    .X(_286_));
 sg13g2_nor2_1 _692_ (.A(net81),
    .B(_284_),
    .Y(_287_));
 sg13g2_nor3_1 _693_ (.A(_210_),
    .B(_286_),
    .C(_287_),
    .Y(_018_));
 sg13g2_o21ai_1 _694_ (.B1(net67),
    .Y(_288_),
    .A1(net80),
    .A2(_286_));
 sg13g2_a21oi_1 _695_ (.A1(net80),
    .A2(_286_),
    .Y(_019_),
    .B1(_288_));
 sg13g2_nor2b_1 _696_ (.A(\square_x_pos[0] ),
    .B_N(net5),
    .Y(_289_));
 sg13g2_xor2_1 _697_ (.B(\square_x_pos[0] ),
    .A(net5),
    .X(_290_));
 sg13g2_nand2_1 _698_ (.Y(_291_),
    .A(net8),
    .B(\square_x_pos[3] ));
 sg13g2_xnor2_1 _699_ (.Y(_292_),
    .A(net8),
    .B(\square_x_pos[3] ));
 sg13g2_or2_1 _700_ (.X(_293_),
    .B(\square_x_pos[2] ),
    .A(net7));
 sg13g2_nor2_1 _701_ (.A(_404_),
    .B(_054_),
    .Y(_294_));
 sg13g2_nand2_1 _702_ (.Y(_295_),
    .A(net7),
    .B(\square_x_pos[2] ));
 sg13g2_and2_1 _703_ (.A(_293_),
    .B(_295_),
    .X(_296_));
 sg13g2_nand2b_1 _704_ (.Y(_297_),
    .B(net76),
    .A_N(net6));
 sg13g2_nor2b_1 _705_ (.A(net77),
    .B_N(net6),
    .Y(_298_));
 sg13g2_a21oi_1 _706_ (.A1(_289_),
    .A2(_297_),
    .Y(_299_),
    .B1(_298_));
 sg13g2_a221oi_1 _707_ (.B2(_289_),
    .C1(_298_),
    .B1(_297_),
    .A1(_293_),
    .Y(_300_),
    .A2(_295_));
 sg13g2_nor2_1 _708_ (.A(net7),
    .B(_054_),
    .Y(_301_));
 sg13g2_o21ai_1 _709_ (.B1(_292_),
    .Y(_302_),
    .A1(_300_),
    .A2(_301_));
 sg13g2_nand2_1 _710_ (.Y(_303_),
    .A(_403_),
    .B(\square_x_pos[3] ));
 sg13g2_nand3_1 _711_ (.B(_302_),
    .C(_303_),
    .A(_056_),
    .Y(_304_));
 sg13g2_nand4_1 _712_ (.B(_057_),
    .C(_302_),
    .A(_056_),
    .Y(_305_),
    .D(_303_));
 sg13g2_nor2_1 _713_ (.A(\square_x_pos[6] ),
    .B(_305_),
    .Y(_306_));
 sg13g2_nand2_2 _714_ (.Y(_307_),
    .A(net68),
    .B(_306_));
 sg13g2_inv_1 _715_ (.Y(_308_),
    .A(_307_));
 sg13g2_nor2_1 _716_ (.A(\square_x_pos[7] ),
    .B(_307_),
    .Y(_309_));
 sg13g2_nor3_1 _717_ (.A(\square_x_pos[7] ),
    .B(\square_x_pos[8] ),
    .C(_307_),
    .Y(_310_));
 sg13g2_nor4_1 _718_ (.A(\square_x_pos[7] ),
    .B(\square_x_pos[8] ),
    .C(\square_x_pos[9] ),
    .D(_307_),
    .Y(_311_));
 sg13g2_and2_1 _719_ (.A(net5),
    .B(\square_x_pos[0] ),
    .X(_312_));
 sg13g2_nand2_1 _720_ (.Y(_313_),
    .A(net5),
    .B(\square_x_pos[0] ));
 sg13g2_xnor2_1 _721_ (.Y(_314_),
    .A(net6),
    .B(net77));
 sg13g2_nand2_1 _722_ (.Y(_315_),
    .A(net6),
    .B(net77));
 sg13g2_o21ai_1 _723_ (.B1(_315_),
    .Y(_316_),
    .A1(_313_),
    .A2(_314_));
 sg13g2_a21oi_1 _724_ (.A1(_296_),
    .A2(_316_),
    .Y(_317_),
    .B1(_294_));
 sg13g2_o21ai_1 _725_ (.B1(_291_),
    .Y(_318_),
    .A1(_292_),
    .A2(_317_));
 sg13g2_inv_1 _726_ (.Y(_319_),
    .A(_318_));
 sg13g2_nand3_1 _727_ (.B(\square_x_pos[5] ),
    .C(_318_),
    .A(\square_x_pos[4] ),
    .Y(_320_));
 sg13g2_or2_1 _728_ (.X(_321_),
    .B(_320_),
    .A(_058_));
 sg13g2_xnor2_1 _729_ (.Y(_322_),
    .A(_058_),
    .B(_320_));
 sg13g2_a21o_1 _730_ (.A2(_318_),
    .A1(\square_x_pos[4] ),
    .B1(\square_x_pos[5] ),
    .X(_323_));
 sg13g2_and2_1 _731_ (.A(_320_),
    .B(_323_),
    .X(_324_));
 sg13g2_nand2_1 _732_ (.Y(_325_),
    .A(_404_),
    .B(_156_));
 sg13g2_nor2_1 _733_ (.A(_404_),
    .B(_156_),
    .Y(_326_));
 sg13g2_a21o_1 _734_ (.A2(_312_),
    .A1(_297_),
    .B1(_298_),
    .X(_327_));
 sg13g2_a221oi_1 _735_ (.B2(_327_),
    .C1(_326_),
    .B1(_325_),
    .A1(net8),
    .Y(_328_),
    .A2(_163_));
 sg13g2_a21oi_1 _736_ (.A1(_403_),
    .A2(_164_),
    .Y(_329_),
    .B1(_328_));
 sg13g2_and2_1 _737_ (.A(_168_),
    .B(_171_),
    .X(_330_));
 sg13g2_nand3b_1 _738_ (.B(_329_),
    .C(_330_),
    .Y(_331_),
    .A_N(_174_));
 sg13g2_xor2_1 _739_ (.B(_317_),
    .A(_292_),
    .X(_332_));
 sg13g2_xnor2_1 _740_ (.Y(_333_),
    .A(_296_),
    .B(_316_));
 sg13g2_xnor2_1 _741_ (.Y(_334_),
    .A(_313_),
    .B(_314_));
 sg13g2_nor4_1 _742_ (.A(\square_x_pos[8] ),
    .B(_290_),
    .C(_333_),
    .D(_334_),
    .Y(_335_));
 sg13g2_nand2_1 _743_ (.Y(_336_),
    .A(_332_),
    .B(_335_));
 sg13g2_a21o_1 _744_ (.A2(_331_),
    .A1(_177_),
    .B1(_336_),
    .X(_337_));
 sg13g2_xnor2_1 _745_ (.Y(_338_),
    .A(_168_),
    .B(_329_));
 sg13g2_o21ai_1 _746_ (.B1(_338_),
    .Y(_339_),
    .A1(_177_),
    .A2(_331_));
 sg13g2_or4_1 _747_ (.A(_322_),
    .B(_324_),
    .C(_337_),
    .D(_339_),
    .X(_340_));
 sg13g2_and3_1 _748_ (.X(_341_),
    .A(_059_),
    .B(_060_),
    .C(_149_));
 sg13g2_nand2b_1 _749_ (.Y(_342_),
    .B(\square_x_pos[9] ),
    .A_N(net68));
 sg13g2_a21oi_2 _750_ (.B1(_342_),
    .Y(_343_),
    .A2(_341_),
    .A1(_331_));
 sg13g2_a21oi_2 _751_ (.B1(_311_),
    .Y(_344_),
    .A2(_343_),
    .A1(_340_));
 sg13g2_mux2_1 _752_ (.A0(\square_x_pos[0] ),
    .A1(_290_),
    .S(net65),
    .X(_020_));
 sg13g2_nand2_1 _753_ (.Y(_345_),
    .A(net5),
    .B(net70));
 sg13g2_xor2_1 _754_ (.B(_345_),
    .A(_334_),
    .X(_346_));
 sg13g2_mux2_1 _755_ (.A0(net77),
    .A1(_346_),
    .S(net65),
    .X(_021_));
 sg13g2_nor2_1 _756_ (.A(\square_x_pos[2] ),
    .B(net65),
    .Y(_347_));
 sg13g2_nor2_1 _757_ (.A(net70),
    .B(_333_),
    .Y(_348_));
 sg13g2_xnor2_1 _758_ (.Y(_349_),
    .A(_296_),
    .B(_299_));
 sg13g2_a21oi_1 _759_ (.A1(net70),
    .A2(_349_),
    .Y(_350_),
    .B1(_348_));
 sg13g2_a21oi_1 _760_ (.A1(_344_),
    .A2(_350_),
    .Y(_022_),
    .B1(_347_));
 sg13g2_nand2b_1 _761_ (.Y(_351_),
    .B(_332_),
    .A_N(net69));
 sg13g2_nor3_1 _762_ (.A(_292_),
    .B(_300_),
    .C(_301_),
    .Y(_352_));
 sg13g2_nand2_1 _763_ (.Y(_353_),
    .A(net69),
    .B(_302_));
 sg13g2_o21ai_1 _764_ (.B1(_351_),
    .Y(_354_),
    .A1(_352_),
    .A2(_353_));
 sg13g2_mux2_1 _765_ (.A0(\square_x_pos[3] ),
    .A1(_354_),
    .S(net65),
    .X(_023_));
 sg13g2_nand3_1 _766_ (.B(_302_),
    .C(_303_),
    .A(net69),
    .Y(_355_));
 sg13g2_o21ai_1 _767_ (.B1(_355_),
    .Y(_356_),
    .A1(net69),
    .A2(_319_));
 sg13g2_nand2_1 _768_ (.Y(_357_),
    .A(net65),
    .B(_356_));
 sg13g2_xnor2_1 _769_ (.Y(_024_),
    .A(\square_x_pos[4] ),
    .B(_357_));
 sg13g2_a221oi_1 _770_ (.B2(_343_),
    .C1(_311_),
    .B1(_340_),
    .A1(net68),
    .Y(_358_),
    .A2(_305_));
 sg13g2_o21ai_1 _771_ (.B1(_358_),
    .Y(_359_),
    .A1(net68),
    .A2(_324_));
 sg13g2_a221oi_1 _772_ (.B2(_343_),
    .C1(_311_),
    .B1(_340_),
    .A1(net68),
    .Y(_360_),
    .A2(_304_));
 sg13g2_o21ai_1 _773_ (.B1(_359_),
    .Y(_025_),
    .A1(_057_),
    .A2(_360_));
 sg13g2_o21ai_1 _774_ (.B1(_307_),
    .Y(_361_),
    .A1(net68),
    .A2(_322_));
 sg13g2_mux2_1 _775_ (.A0(\square_x_pos[6] ),
    .A1(_361_),
    .S(_358_),
    .X(_026_));
 sg13g2_nor2_1 _776_ (.A(net68),
    .B(_321_),
    .Y(_362_));
 sg13g2_o21ai_1 _777_ (.B1(net65),
    .Y(_363_),
    .A1(_308_),
    .A2(_362_));
 sg13g2_xnor2_1 _778_ (.Y(_027_),
    .A(\square_x_pos[7] ),
    .B(_363_));
 sg13g2_nor3_1 _779_ (.A(net68),
    .B(_059_),
    .C(_321_),
    .Y(_364_));
 sg13g2_o21ai_1 _780_ (.B1(net65),
    .Y(_365_),
    .A1(_309_),
    .A2(_364_));
 sg13g2_xnor2_1 _781_ (.Y(_028_),
    .A(\square_x_pos[8] ),
    .B(_365_));
 sg13g2_a21oi_1 _782_ (.A1(\square_x_pos[8] ),
    .A2(_364_),
    .Y(_366_),
    .B1(_310_));
 sg13g2_nand2b_1 _783_ (.Y(_367_),
    .B(net65),
    .A_N(_366_));
 sg13g2_xnor2_1 _784_ (.Y(_029_),
    .A(\square_x_pos[9] ),
    .B(_367_));
 sg13g2_a21oi_2 _785_ (.B1(_267_),
    .Y(_368_),
    .A2(_277_),
    .A1(vert_dir));
 sg13g2_mux2_1 _786_ (.A0(\square_y_pos[0] ),
    .A1(_261_),
    .S(net64),
    .X(_030_));
 sg13g2_nand2_1 _787_ (.Y(_369_),
    .A(net1),
    .B(vert_dir));
 sg13g2_xnor2_1 _788_ (.Y(_370_),
    .A(_263_),
    .B(_369_));
 sg13g2_mux2_1 _789_ (.A0(\square_y_pos[1] ),
    .A1(_370_),
    .S(net64),
    .X(_031_));
 sg13g2_nand2_1 _790_ (.Y(_371_),
    .A(_053_),
    .B(_259_));
 sg13g2_xnor2_1 _791_ (.Y(_372_),
    .A(_252_),
    .B(_270_));
 sg13g2_o21ai_1 _792_ (.B1(_371_),
    .Y(_373_),
    .A1(_053_),
    .A2(_372_));
 sg13g2_mux2_1 _793_ (.A0(net74),
    .A1(_373_),
    .S(net64),
    .X(_032_));
 sg13g2_nand3_1 _794_ (.B(_271_),
    .C(_272_),
    .A(_250_),
    .Y(_374_));
 sg13g2_nand2b_1 _795_ (.Y(_375_),
    .B(_374_),
    .A_N(_273_));
 sg13g2_a21oi_1 _796_ (.A1(vert_dir),
    .A2(_375_),
    .Y(_376_),
    .B1(_266_));
 sg13g2_nand2_1 _797_ (.Y(_377_),
    .A(_368_),
    .B(_376_));
 sg13g2_o21ai_1 _798_ (.B1(_377_),
    .Y(_033_),
    .A1(_048_),
    .A2(net64));
 sg13g2_nand2_2 _799_ (.Y(_378_),
    .A(vert_dir),
    .B(_274_));
 sg13g2_inv_1 _800_ (.Y(_379_),
    .A(_378_));
 sg13g2_a21oi_1 _801_ (.A1(_249_),
    .A2(_257_),
    .Y(_380_),
    .B1(vert_dir));
 sg13g2_o21ai_1 _802_ (.B1(net64),
    .Y(_381_),
    .A1(_379_),
    .A2(_380_));
 sg13g2_xnor2_1 _803_ (.Y(_034_),
    .A(net73),
    .B(_381_));
 sg13g2_and2_1 _804_ (.A(net72),
    .B(_380_),
    .X(_382_));
 sg13g2_nor2_1 _805_ (.A(net73),
    .B(_378_),
    .Y(_383_));
 sg13g2_o21ai_1 _806_ (.B1(_368_),
    .Y(_384_),
    .A1(_382_),
    .A2(_383_));
 sg13g2_xnor2_1 _807_ (.Y(_035_),
    .A(\square_y_pos[5] ),
    .B(_384_));
 sg13g2_nor3_1 _808_ (.A(net72),
    .B(net71),
    .C(_378_),
    .Y(_385_));
 sg13g2_a21oi_1 _809_ (.A1(net71),
    .A2(_382_),
    .Y(_386_),
    .B1(_385_));
 sg13g2_nor2b_1 _810_ (.A(_386_),
    .B_N(net64),
    .Y(_387_));
 sg13g2_xnor2_1 _811_ (.Y(_036_),
    .A(_050_),
    .B(_387_));
 sg13g2_nor4_1 _812_ (.A(net72),
    .B(net71),
    .C(\square_y_pos[6] ),
    .D(_378_),
    .Y(_388_));
 sg13g2_nand4_1 _813_ (.B(net71),
    .C(\square_y_pos[6] ),
    .A(net72),
    .Y(_389_),
    .D(_380_));
 sg13g2_nand2b_1 _814_ (.Y(_390_),
    .B(_389_),
    .A_N(_388_));
 sg13g2_nand2_1 _815_ (.Y(_391_),
    .A(net64),
    .B(_390_));
 sg13g2_xnor2_1 _816_ (.Y(_037_),
    .A(\square_y_pos[7] ),
    .B(_391_));
 sg13g2_a22oi_1 _817_ (.Y(_392_),
    .B1(_276_),
    .B2(_389_),
    .A2(_053_),
    .A1(_051_));
 sg13g2_nand2_1 _818_ (.Y(_393_),
    .A(net64),
    .B(_392_));
 sg13g2_xnor2_1 _819_ (.Y(_038_),
    .A(\square_y_pos[8] ),
    .B(_393_));
 sg13g2_nor3_1 _820_ (.A(\square_y_pos[8] ),
    .B(_267_),
    .C(_276_),
    .Y(_394_));
 sg13g2_nor2b_1 _821_ (.A(_394_),
    .B_N(\square_y_pos[9] ),
    .Y(_039_));
 sg13g2_nor3_1 _822_ (.A(net6),
    .B(net5),
    .C(net8),
    .Y(_395_));
 sg13g2_a21oi_1 _823_ (.A1(_404_),
    .A2(_395_),
    .Y(_396_),
    .B1(_344_));
 sg13g2_xor2_1 _824_ (.B(_396_),
    .A(net69),
    .X(_040_));
 sg13g2_nand2_1 _825_ (.Y(_397_),
    .A(net55),
    .B(net67));
 sg13g2_o21ai_1 _826_ (.B1(_397_),
    .Y(_041_),
    .A1(net55),
    .A2(_217_));
 sg13g2_nand2_1 _827_ (.Y(_398_),
    .A(net50),
    .B(_209_));
 sg13g2_xnor2_1 _828_ (.Y(_399_),
    .A(\hvsync_gen.vpos[0] ),
    .B(net50));
 sg13g2_o21ai_1 _829_ (.B1(_398_),
    .Y(_042_),
    .A1(_217_),
    .A2(_399_));
 sg13g2_nand2_1 _830_ (.Y(_400_),
    .A(net48),
    .B(_209_));
 sg13g2_a21o_1 _831_ (.A2(\hvsync_gen.vpos[1] ),
    .A1(\hvsync_gen.vpos[0] ),
    .B1(net48),
    .X(_401_));
 sg13g2_nand2_1 _832_ (.Y(_402_),
    .A(_212_),
    .B(_401_));
 sg13g2_o21ai_1 _833_ (.B1(_400_),
    .Y(_043_),
    .A1(_217_),
    .A2(_402_));
 sg13g2_dfrbpq_2 _834_ (.RESET_B(net25),
    .D(_002_),
    .Q(\hvsync_gen.vpos[3] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _835_ (.RESET_B(net45),
    .D(_003_),
    .Q(\hvsync_gen.vpos[4] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _836_ (.RESET_B(net44),
    .D(_004_),
    .Q(\hvsync_gen.vpos[5] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _837_ (.RESET_B(net42),
    .D(net63),
    .Q(\hvsync_gen.vpos[6] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _838_ (.RESET_B(net40),
    .D(net101),
    .Q(\hvsync_gen.vpos[7] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _839_ (.RESET_B(net38),
    .D(_007_),
    .Q(\hvsync_gen.vpos[8] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _840_ (.RESET_B(net46),
    .D(net108),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_1 _841_ (.RESET_B(net36),
    .D(net54),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_2_3__leaf_clk));
 sg13g2_dfrbpq_2 _842_ (.RESET_B(net94),
    .D(_009_),
    .Q(vert_dir),
    .CLK(net86));
 sg13g2_dfrbpq_2 _843_ (.RESET_B(net35),
    .D(_010_),
    .Q(\hvsync_gen.hpos[0] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _844_ (.RESET_B(net34),
    .D(_011_),
    .Q(\hvsync_gen.hpos[1] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _845_ (.RESET_B(net33),
    .D(_012_),
    .Q(\hvsync_gen.hpos[2] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _846_ (.RESET_B(net32),
    .D(net60),
    .Q(\hvsync_gen.hpos[3] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _847_ (.RESET_B(net31),
    .D(_014_),
    .Q(\hvsync_gen.hpos[4] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _848_ (.RESET_B(net30),
    .D(_015_),
    .Q(\hvsync_gen.hpos[5] ),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _849_ (.RESET_B(net29),
    .D(_016_),
    .Q(\hvsync_gen.hpos[6] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _850_ (.RESET_B(net28),
    .D(_017_),
    .Q(\hvsync_gen.hpos[7] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _851_ (.RESET_B(net27),
    .D(_018_),
    .Q(\hvsync_gen.hpos[8] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_1 _852_ (.RESET_B(net26),
    .D(_019_),
    .Q(\hvsync_gen.hpos[9] ),
    .CLK(clknet_2_0__leaf_clk));
 sg13g2_dfrbpq_2 _853_ (.RESET_B(net93),
    .D(_020_),
    .Q(\square_x_pos[0] ),
    .CLK(net85));
 sg13g2_dfrbpq_1 _854_ (.RESET_B(net93),
    .D(_021_),
    .Q(\square_x_pos[1] ),
    .CLK(net85));
 sg13g2_dfrbpq_2 _855_ (.RESET_B(net92),
    .D(_022_),
    .Q(\square_x_pos[2] ),
    .CLK(net84));
 sg13g2_dfrbpq_2 _856_ (.RESET_B(net92),
    .D(_023_),
    .Q(\square_x_pos[3] ),
    .CLK(net84));
 sg13g2_dfrbpq_2 _857_ (.RESET_B(net92),
    .D(_024_),
    .Q(\square_x_pos[4] ),
    .CLK(net84));
 sg13g2_dfrbpq_2 _858_ (.RESET_B(net93),
    .D(_025_),
    .Q(\square_x_pos[5] ),
    .CLK(net85));
 sg13g2_dfrbpq_2 _859_ (.RESET_B(net92),
    .D(_026_),
    .Q(\square_x_pos[6] ),
    .CLK(net84));
 sg13g2_dfrbpq_2 _860_ (.RESET_B(net92),
    .D(_027_),
    .Q(\square_x_pos[7] ),
    .CLK(net84));
 sg13g2_dfrbpq_2 _861_ (.RESET_B(net92),
    .D(_028_),
    .Q(\square_x_pos[8] ),
    .CLK(net84));
 sg13g2_dfrbpq_2 _862_ (.RESET_B(net92),
    .D(_029_),
    .Q(\square_x_pos[9] ),
    .CLK(net84));
 sg13g2_dfrbpq_2 _863_ (.RESET_B(net95),
    .D(_030_),
    .Q(\square_y_pos[0] ),
    .CLK(net86));
 sg13g2_dfrbpq_2 _864_ (.RESET_B(net95),
    .D(_031_),
    .Q(\square_y_pos[1] ),
    .CLK(net86));
 sg13g2_dfrbpq_1 _865_ (.RESET_B(net95),
    .D(_032_),
    .Q(\square_y_pos[2] ),
    .CLK(net87));
 sg13g2_dfrbpq_2 _866_ (.RESET_B(net95),
    .D(_033_),
    .Q(\square_y_pos[3] ),
    .CLK(net86));
 sg13g2_dfrbpq_1 _867_ (.RESET_B(net95),
    .D(_034_),
    .Q(\square_y_pos[4] ),
    .CLK(net87));
 sg13g2_dfrbpq_2 _868_ (.RESET_B(net95),
    .D(_035_),
    .Q(\square_y_pos[5] ),
    .CLK(net87));
 sg13g2_dfrbpq_2 _869_ (.RESET_B(net94),
    .D(_036_),
    .Q(\square_y_pos[6] ),
    .CLK(net86));
 sg13g2_dfrbpq_2 _870_ (.RESET_B(net94),
    .D(_037_),
    .Q(\square_y_pos[7] ),
    .CLK(net86));
 sg13g2_dfrbpq_2 _871_ (.RESET_B(net94),
    .D(_038_),
    .Q(\square_y_pos[8] ),
    .CLK(net86));
 sg13g2_dfrbpq_2 _872_ (.RESET_B(net94),
    .D(_039_),
    .Q(\square_y_pos[9] ),
    .CLK(net86));
 sg13g2_dfrbpq_1 _873_ (.RESET_B(net92),
    .D(_040_),
    .Q(horz_dir),
    .CLK(net84));
 sg13g2_dfrbpq_1 _874_ (.RESET_B(net43),
    .D(net99),
    .Q(hsync),
    .CLK(clknet_2_1__leaf_clk));
 sg13g2_dfrbpq_2 _875_ (.RESET_B(net41),
    .D(_041_),
    .Q(\hvsync_gen.vpos[0] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _876_ (.RESET_B(net37),
    .D(net51),
    .Q(\hvsync_gen.vpos[1] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_dfrbpq_2 _877_ (.RESET_B(net39),
    .D(net49),
    .Q(\hvsync_gen.vpos[2] ),
    .CLK(clknet_2_2__leaf_clk));
 sg13g2_tiehi _852__26 (.L_HI(net26));
 sg13g2_tiehi _851__27 (.L_HI(net27));
 sg13g2_tiehi _850__28 (.L_HI(net28));
 sg13g2_tiehi _849__29 (.L_HI(net29));
 sg13g2_tiehi _848__30 (.L_HI(net30));
 sg13g2_tiehi _847__31 (.L_HI(net31));
 sg13g2_tiehi _846__32 (.L_HI(net32));
 sg13g2_tiehi _845__33 (.L_HI(net33));
 sg13g2_tiehi _844__34 (.L_HI(net34));
 sg13g2_tiehi _843__35 (.L_HI(net35));
 sg13g2_tiehi _841__36 (.L_HI(net36));
 sg13g2_tiehi _876__37 (.L_HI(net37));
 sg13g2_tiehi _839__38 (.L_HI(net38));
 sg13g2_tiehi _877__39 (.L_HI(net39));
 sg13g2_tiehi _838__40 (.L_HI(net40));
 sg13g2_tiehi _875__41 (.L_HI(net41));
 sg13g2_tiehi _837__42 (.L_HI(net42));
 sg13g2_tiehi _874__43 (.L_HI(net43));
 sg13g2_tiehi _836__44 (.L_HI(net44));
 sg13g2_tiehi _835__45 (.L_HI(net45));
 sg13g2_tiehi _840__46 (.L_HI(net46));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_vga_example_10 (.L_LO(net10));
 sg13g2_tielo tt_um_vga_example_11 (.L_LO(net11));
 sg13g2_tielo tt_um_vga_example_12 (.L_LO(net12));
 sg13g2_tielo tt_um_vga_example_13 (.L_LO(net13));
 sg13g2_tielo tt_um_vga_example_14 (.L_LO(net14));
 sg13g2_tielo tt_um_vga_example_15 (.L_LO(net15));
 sg13g2_tielo tt_um_vga_example_16 (.L_LO(net16));
 sg13g2_tielo tt_um_vga_example_17 (.L_LO(net17));
 sg13g2_tielo tt_um_vga_example_18 (.L_LO(net18));
 sg13g2_tielo tt_um_vga_example_19 (.L_LO(net19));
 sg13g2_tielo tt_um_vga_example_20 (.L_LO(net20));
 sg13g2_tielo tt_um_vga_example_21 (.L_LO(net21));
 sg13g2_tielo tt_um_vga_example_22 (.L_LO(net22));
 sg13g2_tielo tt_um_vga_example_23 (.L_LO(net23));
 sg13g2_tielo tt_um_vga_example_24 (.L_LO(net24));
 sg13g2_tiehi _834__25 (.L_HI(net25));
 sg13g2_buf_1 _916_ (.A(uo_out[5]),
    .X(uo_out[0]));
 sg13g2_buf_1 _917_ (.A(uo_out[6]),
    .X(uo_out[1]));
 sg13g2_buf_1 _918_ (.A(uo_out[6]),
    .X(uo_out[2]));
 sg13g2_buf_1 _919_ (.A(net85),
    .X(uo_out[3]));
 sg13g2_buf_1 _920_ (.A(uo_out[6]),
    .X(uo_out[4]));
 sg13g2_buf_1 _921_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout64 (.A(_368_),
    .X(net64));
 sg13g2_buf_8 fanout65 (.A(_344_),
    .X(net65));
 sg13g2_buf_8 fanout66 (.A(_217_),
    .X(net66));
 sg13g2_buf_8 fanout67 (.A(_209_),
    .X(net67));
 sg13g2_buf_8 fanout68 (.A(net70),
    .X(net68));
 sg13g2_buf_1 fanout69 (.A(net70),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(horz_dir),
    .X(net70));
 sg13g2_buf_8 fanout71 (.A(\square_y_pos[5] ),
    .X(net71));
 sg13g2_buf_8 fanout72 (.A(net73),
    .X(net72));
 sg13g2_buf_8 fanout73 (.A(\square_y_pos[4] ),
    .X(net73));
 sg13g2_buf_8 fanout74 (.A(\square_y_pos[2] ),
    .X(net74));
 sg13g2_buf_8 fanout75 (.A(\square_y_pos[1] ),
    .X(net75));
 sg13g2_buf_8 fanout76 (.A(\square_x_pos[1] ),
    .X(net76));
 sg13g2_buf_1 fanout77 (.A(\square_x_pos[1] ),
    .X(net77));
 sg13g2_buf_8 fanout78 (.A(net48),
    .X(net78));
 sg13g2_buf_8 fanout79 (.A(net50),
    .X(net79));
 sg13g2_buf_8 fanout80 (.A(net103),
    .X(net80));
 sg13g2_buf_8 fanout81 (.A(net98),
    .X(net81));
 sg13g2_buf_8 fanout82 (.A(net111),
    .X(net82));
 sg13g2_buf_8 fanout83 (.A(net102),
    .X(net83));
 sg13g2_buf_8 fanout84 (.A(net85),
    .X(net84));
 sg13g2_buf_8 fanout85 (.A(net87),
    .X(net85));
 sg13g2_buf_8 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_8 fanout87 (.A(\hvsync_gen.vsync ),
    .X(net87));
 sg13g2_buf_8 fanout88 (.A(net107),
    .X(net88));
 sg13g2_buf_8 fanout89 (.A(net110),
    .X(net89));
 sg13g2_buf_8 fanout90 (.A(net109),
    .X(net90));
 sg13g2_buf_8 fanout91 (.A(net52),
    .X(net91));
 sg13g2_buf_8 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_8 fanout93 (.A(rst_n),
    .X(net93));
 sg13g2_buf_8 fanout94 (.A(rst_n),
    .X(net94));
 sg13g2_buf_8 fanout95 (.A(rst_n),
    .X(net95));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_tielo tt_um_vga_example_9 (.L_LO(net9));
 sg13g2_buf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_2_0__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_2_1__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\hvsync_gen.hpos[0] ),
    .X(net47));
 sg13g2_dlygate4sd3_1 hold2 (.A(\hvsync_gen.vpos[2] ),
    .X(net48));
 sg13g2_dlygate4sd3_1 hold3 (.A(_043_),
    .X(net49));
 sg13g2_dlygate4sd3_1 hold4 (.A(\hvsync_gen.vpos[1] ),
    .X(net50));
 sg13g2_dlygate4sd3_1 hold5 (.A(_042_),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold6 (.A(\hvsync_gen.vpos[3] ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold7 (.A(_071_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold8 (.A(_001_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold9 (.A(\hvsync_gen.vpos[0] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold10 (.A(\hvsync_gen.hpos[5] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold11 (.A(_208_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold12 (.A(\hvsync_gen.hpos[3] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold13 (.A(_279_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold14 (.A(_013_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold15 (.A(\hvsync_gen.hpos[1] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold16 (.A(\hvsync_gen.vpos[6] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold17 (.A(_005_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold18 (.A(\hvsync_gen.hpos[6] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold19 (.A(_283_),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold20 (.A(\hvsync_gen.hpos[8] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold21 (.A(_000_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold22 (.A(\hvsync_gen.vpos[7] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold23 (.A(_006_),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold24 (.A(\hvsync_gen.hpos[2] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold25 (.A(\hvsync_gen.hpos[9] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold26 (.A(\hvsync_gen.hpos[4] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold27 (.A(\hvsync_gen.vpos[8] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold28 (.A(_233_),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold29 (.A(\hvsync_gen.vpos[9] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold30 (.A(_008_),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold31 (.A(\hvsync_gen.vpos[4] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold32 (.A(\hvsync_gen.vpos[5] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold33 (.A(\hvsync_gen.hpos[7] ),
    .X(net111));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_8 FILLER_10_315 ();
 sg13g2_decap_8 FILLER_10_322 ();
 sg13g2_decap_8 FILLER_10_329 ();
 sg13g2_decap_8 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_343 ();
 sg13g2_decap_8 FILLER_10_350 ();
 sg13g2_decap_8 FILLER_10_357 ();
 sg13g2_decap_8 FILLER_10_364 ();
 sg13g2_decap_8 FILLER_10_371 ();
 sg13g2_decap_8 FILLER_10_378 ();
 sg13g2_decap_8 FILLER_10_385 ();
 sg13g2_decap_8 FILLER_10_392 ();
 sg13g2_decap_8 FILLER_10_399 ();
 sg13g2_fill_2 FILLER_10_406 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_fill_2 FILLER_11_406 ();
 sg13g2_fill_1 FILLER_11_408 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_fill_2 FILLER_14_406 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_8 FILLER_15_308 ();
 sg13g2_decap_8 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_322 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_decap_8 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_343 ();
 sg13g2_decap_8 FILLER_15_350 ();
 sg13g2_decap_8 FILLER_15_357 ();
 sg13g2_decap_8 FILLER_15_364 ();
 sg13g2_decap_8 FILLER_15_371 ();
 sg13g2_decap_8 FILLER_15_378 ();
 sg13g2_decap_8 FILLER_15_385 ();
 sg13g2_decap_8 FILLER_15_392 ();
 sg13g2_decap_8 FILLER_15_399 ();
 sg13g2_fill_2 FILLER_15_406 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_fill_2 FILLER_16_406 ();
 sg13g2_fill_1 FILLER_16_408 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_fill_2 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_fill_2 FILLER_20_263 ();
 sg13g2_fill_1 FILLER_20_265 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_4 FILLER_20_403 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_4 FILLER_21_133 ();
 sg13g2_fill_1 FILLER_21_137 ();
 sg13g2_decap_4 FILLER_21_169 ();
 sg13g2_fill_2 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_202 ();
 sg13g2_fill_1 FILLER_21_204 ();
 sg13g2_decap_8 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_216 ();
 sg13g2_decap_8 FILLER_21_223 ();
 sg13g2_decap_4 FILLER_21_230 ();
 sg13g2_fill_2 FILLER_21_234 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_4 FILLER_21_312 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_2 FILLER_21_322 ();
 sg13g2_decap_4 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_8 FILLER_21_383 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_4 FILLER_22_105 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_114 ();
 sg13g2_decap_4 FILLER_22_121 ();
 sg13g2_fill_1 FILLER_22_125 ();
 sg13g2_fill_2 FILLER_22_139 ();
 sg13g2_fill_1 FILLER_22_141 ();
 sg13g2_decap_8 FILLER_22_152 ();
 sg13g2_decap_4 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_163 ();
 sg13g2_fill_1 FILLER_22_288 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_4 FILLER_22_342 ();
 sg13g2_fill_1 FILLER_22_346 ();
 sg13g2_fill_2 FILLER_22_355 ();
 sg13g2_fill_1 FILLER_22_357 ();
 sg13g2_decap_8 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_393 ();
 sg13g2_decap_8 FILLER_22_400 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_4 FILLER_23_98 ();
 sg13g2_fill_2 FILLER_23_153 ();
 sg13g2_fill_1 FILLER_23_155 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_2 FILLER_23_215 ();
 sg13g2_decap_4 FILLER_23_226 ();
 sg13g2_fill_1 FILLER_23_230 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_4 FILLER_23_249 ();
 sg13g2_fill_1 FILLER_23_258 ();
 sg13g2_decap_8 FILLER_23_296 ();
 sg13g2_decap_4 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_307 ();
 sg13g2_fill_2 FILLER_23_321 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_fill_1 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_390 ();
 sg13g2_decap_8 FILLER_23_397 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_4 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_4 FILLER_24_119 ();
 sg13g2_fill_2 FILLER_24_123 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_4 FILLER_24_261 ();
 sg13g2_fill_2 FILLER_24_265 ();
 sg13g2_fill_2 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_decap_4 FILLER_24_283 ();
 sg13g2_decap_4 FILLER_24_302 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_fill_2 FILLER_24_334 ();
 sg13g2_fill_1 FILLER_24_336 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_392 ();
 sg13g2_decap_8 FILLER_24_399 ();
 sg13g2_fill_2 FILLER_24_406 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_fill_2 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_152 ();
 sg13g2_fill_1 FILLER_25_159 ();
 sg13g2_fill_1 FILLER_25_217 ();
 sg13g2_fill_2 FILLER_25_227 ();
 sg13g2_fill_2 FILLER_25_271 ();
 sg13g2_fill_1 FILLER_25_284 ();
 sg13g2_fill_2 FILLER_25_296 ();
 sg13g2_fill_1 FILLER_25_298 ();
 sg13g2_fill_2 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_325 ();
 sg13g2_fill_2 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_345 ();
 sg13g2_fill_2 FILLER_25_359 ();
 sg13g2_fill_1 FILLER_25_361 ();
 sg13g2_fill_2 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_fill_2 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_4 FILLER_26_77 ();
 sg13g2_fill_1 FILLER_26_109 ();
 sg13g2_fill_1 FILLER_26_164 ();
 sg13g2_fill_2 FILLER_26_199 ();
 sg13g2_fill_2 FILLER_26_278 ();
 sg13g2_fill_1 FILLER_26_284 ();
 sg13g2_fill_1 FILLER_26_290 ();
 sg13g2_fill_1 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_fill_2 FILLER_26_406 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_4 FILLER_27_56 ();
 sg13g2_decap_4 FILLER_27_68 ();
 sg13g2_decap_8 FILLER_27_85 ();
 sg13g2_decap_8 FILLER_27_92 ();
 sg13g2_decap_8 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_108 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_fill_2 FILLER_27_126 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_fill_2 FILLER_27_134 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_fill_1 FILLER_27_177 ();
 sg13g2_decap_4 FILLER_27_202 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_4 FILLER_27_217 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_1 FILLER_27_281 ();
 sg13g2_fill_1 FILLER_27_288 ();
 sg13g2_fill_1 FILLER_27_329 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_fill_1 FILLER_27_350 ();
 sg13g2_fill_2 FILLER_27_360 ();
 sg13g2_fill_1 FILLER_27_362 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_2 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_82 ();
 sg13g2_fill_2 FILLER_28_89 ();
 sg13g2_fill_1 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_96 ();
 sg13g2_fill_2 FILLER_28_140 ();
 sg13g2_fill_2 FILLER_28_159 ();
 sg13g2_fill_2 FILLER_28_166 ();
 sg13g2_fill_2 FILLER_28_177 ();
 sg13g2_fill_1 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_1 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_190 ();
 sg13g2_fill_2 FILLER_28_207 ();
 sg13g2_decap_8 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_227 ();
 sg13g2_decap_4 FILLER_28_232 ();
 sg13g2_fill_2 FILLER_28_236 ();
 sg13g2_fill_2 FILLER_28_244 ();
 sg13g2_fill_1 FILLER_28_256 ();
 sg13g2_decap_8 FILLER_28_261 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_decap_4 FILLER_28_279 ();
 sg13g2_fill_2 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_306 ();
 sg13g2_fill_1 FILLER_28_308 ();
 sg13g2_fill_2 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_314 ();
 sg13g2_fill_2 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_328 ();
 sg13g2_fill_2 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_338 ();
 sg13g2_fill_1 FILLER_28_355 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_fill_2 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_4 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_decap_8 FILLER_29_107 ();
 sg13g2_decap_8 FILLER_29_114 ();
 sg13g2_decap_4 FILLER_29_121 ();
 sg13g2_fill_2 FILLER_29_125 ();
 sg13g2_decap_8 FILLER_29_132 ();
 sg13g2_decap_8 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_146 ();
 sg13g2_fill_1 FILLER_29_148 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_fill_1 FILLER_29_157 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_4 FILLER_29_176 ();
 sg13g2_fill_1 FILLER_29_180 ();
 sg13g2_fill_2 FILLER_29_226 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_fill_2 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_275 ();
 sg13g2_fill_1 FILLER_29_285 ();
 sg13g2_fill_2 FILLER_29_307 ();
 sg13g2_fill_2 FILLER_29_314 ();
 sg13g2_fill_2 FILLER_29_321 ();
 sg13g2_fill_1 FILLER_29_323 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_4 FILLER_29_383 ();
 sg13g2_fill_2 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_58 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_fill_1 FILLER_30_79 ();
 sg13g2_decap_8 FILLER_30_90 ();
 sg13g2_decap_8 FILLER_30_97 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_decap_4 FILLER_30_114 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_decap_4 FILLER_30_136 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_decap_4 FILLER_30_205 ();
 sg13g2_fill_2 FILLER_30_217 ();
 sg13g2_fill_1 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_228 ();
 sg13g2_decap_4 FILLER_30_235 ();
 sg13g2_fill_1 FILLER_30_244 ();
 sg13g2_decap_8 FILLER_30_253 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_fill_2 FILLER_30_277 ();
 sg13g2_fill_2 FILLER_30_286 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_297 ();
 sg13g2_decap_4 FILLER_30_303 ();
 sg13g2_fill_2 FILLER_30_307 ();
 sg13g2_decap_8 FILLER_30_321 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_fill_1 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_fill_2 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_75 ();
 sg13g2_decap_8 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_103 ();
 sg13g2_fill_1 FILLER_31_112 ();
 sg13g2_decap_4 FILLER_31_118 ();
 sg13g2_fill_2 FILLER_31_122 ();
 sg13g2_decap_4 FILLER_31_134 ();
 sg13g2_fill_1 FILLER_31_138 ();
 sg13g2_fill_1 FILLER_31_197 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_4 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_214 ();
 sg13g2_fill_2 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_235 ();
 sg13g2_decap_4 FILLER_31_260 ();
 sg13g2_fill_1 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_fill_2 FILLER_31_307 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_decap_4 FILLER_31_354 ();
 sg13g2_fill_2 FILLER_31_358 ();
 sg13g2_decap_8 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_375 ();
 sg13g2_fill_2 FILLER_31_384 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_56 ();
 sg13g2_fill_2 FILLER_32_78 ();
 sg13g2_decap_8 FILLER_32_101 ();
 sg13g2_decap_8 FILLER_32_108 ();
 sg13g2_decap_4 FILLER_32_115 ();
 sg13g2_decap_8 FILLER_32_138 ();
 sg13g2_decap_8 FILLER_32_145 ();
 sg13g2_fill_2 FILLER_32_152 ();
 sg13g2_fill_1 FILLER_32_154 ();
 sg13g2_decap_8 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_decap_4 FILLER_32_177 ();
 sg13g2_fill_2 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_211 ();
 sg13g2_fill_2 FILLER_32_218 ();
 sg13g2_decap_8 FILLER_32_229 ();
 sg13g2_fill_2 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_238 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_decap_4 FILLER_32_250 ();
 sg13g2_fill_2 FILLER_32_254 ();
 sg13g2_decap_8 FILLER_32_260 ();
 sg13g2_decap_4 FILLER_32_267 ();
 sg13g2_fill_1 FILLER_32_271 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_4 FILLER_32_291 ();
 sg13g2_fill_2 FILLER_32_295 ();
 sg13g2_decap_8 FILLER_32_301 ();
 sg13g2_decap_8 FILLER_32_308 ();
 sg13g2_decap_8 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_322 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_fill_2 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_342 ();
 sg13g2_decap_8 FILLER_32_349 ();
 sg13g2_decap_8 FILLER_32_356 ();
 sg13g2_decap_4 FILLER_32_363 ();
 sg13g2_fill_1 FILLER_32_367 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_fill_2 FILLER_33_28 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_2 FILLER_33_67 ();
 sg13g2_fill_1 FILLER_33_69 ();
 sg13g2_decap_8 FILLER_33_75 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_fill_2 FILLER_33_99 ();
 sg13g2_decap_8 FILLER_33_129 ();
 sg13g2_decap_4 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_144 ();
 sg13g2_fill_1 FILLER_33_148 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_180 ();
 sg13g2_decap_4 FILLER_33_187 ();
 sg13g2_fill_1 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_202 ();
 sg13g2_decap_8 FILLER_33_209 ();
 sg13g2_decap_8 FILLER_33_216 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_260 ();
 sg13g2_decap_4 FILLER_33_266 ();
 sg13g2_fill_1 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_281 ();
 sg13g2_fill_2 FILLER_33_306 ();
 sg13g2_fill_1 FILLER_33_308 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_fill_1 FILLER_33_353 ();
 sg13g2_decap_8 FILLER_33_382 ();
 sg13g2_decap_4 FILLER_33_389 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_65 ();
 sg13g2_fill_1 FILLER_34_78 ();
 sg13g2_decap_8 FILLER_34_88 ();
 sg13g2_fill_1 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_101 ();
 sg13g2_fill_1 FILLER_34_106 ();
 sg13g2_decap_8 FILLER_34_111 ();
 sg13g2_decap_8 FILLER_34_118 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_4 FILLER_34_135 ();
 sg13g2_fill_2 FILLER_34_139 ();
 sg13g2_decap_8 FILLER_34_160 ();
 sg13g2_decap_4 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_decap_8 FILLER_34_192 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_211 ();
 sg13g2_decap_8 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_232 ();
 sg13g2_decap_8 FILLER_34_239 ();
 sg13g2_decap_8 FILLER_34_246 ();
 sg13g2_decap_4 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_281 ();
 sg13g2_decap_4 FILLER_34_288 ();
 sg13g2_fill_1 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_329 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_408 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_2 FILLER_35_75 ();
 sg13g2_fill_1 FILLER_35_77 ();
 sg13g2_fill_2 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_125 ();
 sg13g2_decap_4 FILLER_35_144 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_1 FILLER_35_189 ();
 sg13g2_decap_4 FILLER_35_218 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_decap_4 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_4 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_304 ();
 sg13g2_fill_1 FILLER_35_306 ();
 sg13g2_decap_4 FILLER_35_311 ();
 sg13g2_fill_1 FILLER_35_315 ();
 sg13g2_fill_1 FILLER_35_325 ();
 sg13g2_decap_4 FILLER_35_331 ();
 sg13g2_fill_2 FILLER_35_346 ();
 sg13g2_fill_1 FILLER_35_348 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_4 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_406 ();
 sg13g2_fill_1 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_decap_4 FILLER_36_71 ();
 sg13g2_decap_8 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_92 ();
 sg13g2_fill_2 FILLER_36_106 ();
 sg13g2_fill_1 FILLER_36_108 ();
 sg13g2_fill_2 FILLER_36_122 ();
 sg13g2_fill_2 FILLER_36_132 ();
 sg13g2_fill_1 FILLER_36_134 ();
 sg13g2_fill_2 FILLER_36_140 ();
 sg13g2_decap_4 FILLER_36_148 ();
 sg13g2_fill_1 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_167 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_174 ();
 sg13g2_decap_8 FILLER_36_183 ();
 sg13g2_decap_8 FILLER_36_190 ();
 sg13g2_decap_4 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_201 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_fill_1 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_244 ();
 sg13g2_decap_8 FILLER_36_251 ();
 sg13g2_decap_4 FILLER_36_258 ();
 sg13g2_fill_2 FILLER_36_266 ();
 sg13g2_fill_2 FILLER_36_273 ();
 sg13g2_fill_1 FILLER_36_280 ();
 sg13g2_fill_2 FILLER_36_336 ();
 sg13g2_fill_1 FILLER_36_338 ();
 sg13g2_decap_4 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_4 FILLER_37_49 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_decap_8 FILLER_37_83 ();
 sg13g2_fill_1 FILLER_37_90 ();
 sg13g2_fill_2 FILLER_37_123 ();
 sg13g2_fill_2 FILLER_37_165 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_fill_1 FILLER_37_214 ();
 sg13g2_fill_1 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_decap_8 FILLER_37_269 ();
 sg13g2_decap_8 FILLER_37_276 ();
 sg13g2_decap_8 FILLER_37_283 ();
 sg13g2_decap_8 FILLER_37_290 ();
 sg13g2_decap_8 FILLER_37_297 ();
 sg13g2_decap_8 FILLER_37_304 ();
 sg13g2_fill_1 FILLER_37_311 ();
 sg13g2_fill_2 FILLER_37_325 ();
 sg13g2_fill_2 FILLER_37_342 ();
 sg13g2_fill_2 FILLER_37_354 ();
 sg13g2_decap_4 FILLER_37_365 ();
 sg13g2_decap_8 FILLER_37_379 ();
 sg13g2_decap_8 FILLER_37_386 ();
 sg13g2_decap_8 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_400 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_76 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_206 ();
 sg13g2_decap_8 FILLER_38_213 ();
 sg13g2_decap_8 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_227 ();
 sg13g2_decap_8 FILLER_38_241 ();
 sg13g2_decap_4 FILLER_38_248 ();
 sg13g2_fill_1 FILLER_38_280 ();
 sg13g2_fill_2 FILLER_38_309 ();
 sg13g2_fill_1 FILLER_38_311 ();
 sg13g2_decap_4 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_334 ();
 sg13g2_fill_2 FILLER_38_341 ();
 sg13g2_fill_1 FILLER_38_343 ();
 sg13g2_fill_1 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net9;
 assign uio_oe[1] = net10;
 assign uio_oe[2] = net11;
 assign uio_oe[3] = net12;
 assign uio_oe[4] = net13;
 assign uio_oe[5] = net14;
 assign uio_oe[6] = net15;
 assign uio_oe[7] = net16;
 assign uio_out[0] = net17;
 assign uio_out[1] = net18;
 assign uio_out[2] = net19;
 assign uio_out[3] = net20;
 assign uio_out[4] = net21;
 assign uio_out[5] = net22;
 assign uio_out[6] = net23;
 assign uio_out[7] = net24;
endmodule
