module tt_um_tt_tinyQV (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire net1435;
 wire clk_regs;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire \addr[0] ;
 wire \addr[10] ;
 wire \addr[11] ;
 wire \addr[12] ;
 wire \addr[13] ;
 wire \addr[14] ;
 wire \addr[15] ;
 wire \addr[16] ;
 wire \addr[17] ;
 wire \addr[18] ;
 wire \addr[19] ;
 wire \addr[1] ;
 wire \addr[20] ;
 wire \addr[21] ;
 wire \addr[22] ;
 wire \addr[23] ;
 wire \addr[24] ;
 wire \addr[25] ;
 wire \addr[26] ;
 wire \addr[27] ;
 wire \addr[2] ;
 wire \addr[3] ;
 wire \addr[4] ;
 wire \addr[5] ;
 wire \addr[6] ;
 wire \addr[7] ;
 wire \addr[8] ;
 wire \addr[9] ;
 wire \data_to_write[0] ;
 wire \data_to_write[10] ;
 wire \data_to_write[11] ;
 wire \data_to_write[12] ;
 wire \data_to_write[13] ;
 wire \data_to_write[14] ;
 wire \data_to_write[15] ;
 wire \data_to_write[16] ;
 wire \data_to_write[17] ;
 wire \data_to_write[18] ;
 wire \data_to_write[19] ;
 wire \data_to_write[1] ;
 wire \data_to_write[20] ;
 wire \data_to_write[21] ;
 wire \data_to_write[22] ;
 wire \data_to_write[23] ;
 wire \data_to_write[24] ;
 wire \data_to_write[25] ;
 wire \data_to_write[26] ;
 wire \data_to_write[27] ;
 wire \data_to_write[28] ;
 wire \data_to_write[29] ;
 wire \data_to_write[2] ;
 wire \data_to_write[30] ;
 wire \data_to_write[31] ;
 wire \data_to_write[3] ;
 wire \data_to_write[4] ;
 wire \data_to_write[5] ;
 wire \data_to_write[6] ;
 wire \data_to_write[7] ;
 wire \data_to_write[8] ;
 wire \data_to_write[9] ;
 wire debug_data_continue;
 wire debug_instr_valid;
 wire \debug_rd[0] ;
 wire \debug_rd[1] ;
 wire \debug_rd[2] ;
 wire \debug_rd[3] ;
 wire \debug_rd_r[0] ;
 wire \debug_rd_r[1] ;
 wire \debug_rd_r[2] ;
 wire \debug_rd_r[3] ;
 wire debug_register_data;
 wire debug_uart_txd;
 wire \gpio_out_sel[6] ;
 wire \gpio_out_sel[7] ;
 wire \i_debug_uart_tx.cycle_counter[0] ;
 wire \i_debug_uart_tx.cycle_counter[1] ;
 wire \i_debug_uart_tx.cycle_counter[2] ;
 wire \i_debug_uart_tx.cycle_counter[3] ;
 wire \i_debug_uart_tx.cycle_counter[4] ;
 wire \i_debug_uart_tx.data_to_send[0] ;
 wire \i_debug_uart_tx.data_to_send[1] ;
 wire \i_debug_uart_tx.data_to_send[2] ;
 wire \i_debug_uart_tx.data_to_send[3] ;
 wire \i_debug_uart_tx.data_to_send[4] ;
 wire \i_debug_uart_tx.data_to_send[5] ;
 wire \i_debug_uart_tx.data_to_send[6] ;
 wire \i_debug_uart_tx.data_to_send[7] ;
 wire \i_debug_uart_tx.fsm_state[0] ;
 wire \i_debug_uart_tx.fsm_state[1] ;
 wire \i_debug_uart_tx.fsm_state[2] ;
 wire \i_debug_uart_tx.fsm_state[3] ;
 wire \i_debug_uart_tx.resetn ;
 wire \i_peripherals.data_out[0] ;
 wire \i_peripherals.data_out[10] ;
 wire \i_peripherals.data_out[11] ;
 wire \i_peripherals.data_out[12] ;
 wire \i_peripherals.data_out[13] ;
 wire \i_peripherals.data_out[14] ;
 wire \i_peripherals.data_out[15] ;
 wire \i_peripherals.data_out[16] ;
 wire \i_peripherals.data_out[17] ;
 wire \i_peripherals.data_out[18] ;
 wire \i_peripherals.data_out[19] ;
 wire \i_peripherals.data_out[1] ;
 wire \i_peripherals.data_out[20] ;
 wire \i_peripherals.data_out[21] ;
 wire \i_peripherals.data_out[22] ;
 wire \i_peripherals.data_out[23] ;
 wire \i_peripherals.data_out[24] ;
 wire \i_peripherals.data_out[25] ;
 wire \i_peripherals.data_out[26] ;
 wire \i_peripherals.data_out[27] ;
 wire \i_peripherals.data_out[28] ;
 wire \i_peripherals.data_out[29] ;
 wire \i_peripherals.data_out[2] ;
 wire \i_peripherals.data_out[30] ;
 wire \i_peripherals.data_out[31] ;
 wire \i_peripherals.data_out[3] ;
 wire \i_peripherals.data_out[4] ;
 wire \i_peripherals.data_out[5] ;
 wire \i_peripherals.data_out[6] ;
 wire \i_peripherals.data_out[7] ;
 wire \i_peripherals.data_out[8] ;
 wire \i_peripherals.data_out[9] ;
 wire \i_peripherals.data_out_hold ;
 wire \i_peripherals.data_ready_r ;
 wire \i_peripherals.func_sel[0] ;
 wire \i_peripherals.func_sel[10] ;
 wire \i_peripherals.func_sel[11] ;
 wire \i_peripherals.func_sel[12] ;
 wire \i_peripherals.func_sel[13] ;
 wire \i_peripherals.func_sel[14] ;
 wire \i_peripherals.func_sel[15] ;
 wire \i_peripherals.func_sel[16] ;
 wire \i_peripherals.func_sel[17] ;
 wire \i_peripherals.func_sel[18] ;
 wire \i_peripherals.func_sel[19] ;
 wire \i_peripherals.func_sel[1] ;
 wire \i_peripherals.func_sel[20] ;
 wire \i_peripherals.func_sel[21] ;
 wire \i_peripherals.func_sel[22] ;
 wire \i_peripherals.func_sel[23] ;
 wire \i_peripherals.func_sel[24] ;
 wire \i_peripherals.func_sel[25] ;
 wire \i_peripherals.func_sel[26] ;
 wire \i_peripherals.func_sel[27] ;
 wire \i_peripherals.func_sel[28] ;
 wire \i_peripherals.func_sel[29] ;
 wire \i_peripherals.func_sel[2] ;
 wire \i_peripherals.func_sel[30] ;
 wire \i_peripherals.func_sel[31] ;
 wire \i_peripherals.func_sel[32] ;
 wire \i_peripherals.func_sel[33] ;
 wire \i_peripherals.func_sel[34] ;
 wire \i_peripherals.func_sel[35] ;
 wire \i_peripherals.func_sel[36] ;
 wire \i_peripherals.func_sel[37] ;
 wire \i_peripherals.func_sel[38] ;
 wire \i_peripherals.func_sel[39] ;
 wire \i_peripherals.func_sel[3] ;
 wire \i_peripherals.func_sel[40] ;
 wire \i_peripherals.func_sel[41] ;
 wire \i_peripherals.func_sel[42] ;
 wire \i_peripherals.func_sel[43] ;
 wire \i_peripherals.func_sel[44] ;
 wire \i_peripherals.func_sel[45] ;
 wire \i_peripherals.func_sel[46] ;
 wire \i_peripherals.func_sel[47] ;
 wire \i_peripherals.func_sel[4] ;
 wire \i_peripherals.func_sel[5] ;
 wire \i_peripherals.func_sel[6] ;
 wire \i_peripherals.func_sel[7] ;
 wire \i_peripherals.func_sel[8] ;
 wire \i_peripherals.func_sel[9] ;
 wire \i_peripherals.gpio_out[0] ;
 wire \i_peripherals.gpio_out[1] ;
 wire \i_peripherals.gpio_out[2] ;
 wire \i_peripherals.gpio_out[3] ;
 wire \i_peripherals.gpio_out[4] ;
 wire \i_peripherals.gpio_out[5] ;
 wire \i_peripherals.gpio_out[6] ;
 wire \i_peripherals.gpio_out[7] ;
 wire \i_peripherals.i_uart.baud_divider[0] ;
 wire \i_peripherals.i_uart.baud_divider[10] ;
 wire \i_peripherals.i_uart.baud_divider[11] ;
 wire \i_peripherals.i_uart.baud_divider[12] ;
 wire \i_peripherals.i_uart.baud_divider[1] ;
 wire \i_peripherals.i_uart.baud_divider[2] ;
 wire \i_peripherals.i_uart.baud_divider[3] ;
 wire \i_peripherals.i_uart.baud_divider[4] ;
 wire \i_peripherals.i_uart.baud_divider[5] ;
 wire \i_peripherals.i_uart.baud_divider[6] ;
 wire \i_peripherals.i_uart.baud_divider[7] ;
 wire \i_peripherals.i_uart.baud_divider[8] ;
 wire \i_peripherals.i_uart.baud_divider[9] ;
 wire \i_peripherals.i_uart.i_uart_rx.bit_sample ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[0] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[10] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[11] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[12] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[2] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[3] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[4] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[6] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[7] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[8] ;
 wire \i_peripherals.i_uart.i_uart_rx.cycle_counter[9] ;
 wire \i_peripherals.i_uart.i_uart_rx.fsm_state[0] ;
 wire \i_peripherals.i_uart.i_uart_rx.fsm_state[1] ;
 wire \i_peripherals.i_uart.i_uart_rx.fsm_state[2] ;
 wire \i_peripherals.i_uart.i_uart_rx.fsm_state[3] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[0] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[1] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[2] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[3] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[4] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[5] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[6] ;
 wire \i_peripherals.i_uart.i_uart_rx.recieved_data[7] ;
 wire \i_peripherals.i_uart.i_uart_rx.uart_rts ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[0] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[10] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[11] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[12] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[1] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[2] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[3] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[4] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[5] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[6] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[7] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[8] ;
 wire \i_peripherals.i_uart.i_uart_tx.cycle_counter[9] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[0] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[1] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[2] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[3] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[4] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[5] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[6] ;
 wire \i_peripherals.i_uart.i_uart_tx.data_to_send[7] ;
 wire \i_peripherals.i_uart.i_uart_tx.fsm_state[0] ;
 wire \i_peripherals.i_uart.i_uart_tx.fsm_state[1] ;
 wire \i_peripherals.i_uart.i_uart_tx.fsm_state[2] ;
 wire \i_peripherals.i_uart.i_uart_tx.fsm_state[3] ;
 wire \i_peripherals.i_uart.i_uart_tx.txd_reg ;
 wire \i_peripherals.i_uart.rxd_select ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[0] ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[1] ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[2] ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[3] ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[4] ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[5] ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[6] ;
 wire \i_peripherals.i_uart.uart_rx_buf_data[7] ;
 wire \i_peripherals.i_uart.uart_rx_buffered ;
 wire \i_peripherals.i_uart.ui_in[0] ;
 wire \i_peripherals.i_uart.ui_in[1] ;
 wire \i_peripherals.i_uart.ui_in[2] ;
 wire \i_peripherals.i_uart.ui_in[3] ;
 wire \i_peripherals.i_uart.ui_in[4] ;
 wire \i_peripherals.i_uart.ui_in[5] ;
 wire \i_peripherals.i_uart.ui_in[6] ;
 wire \i_peripherals.i_uart.ui_in[7] ;
 wire \i_peripherals.i_user_peri39._GEN[0] ;
 wire \i_peripherals.i_user_peri39._GEN[100] ;
 wire \i_peripherals.i_user_peri39._GEN[101] ;
 wire \i_peripherals.i_user_peri39._GEN[102] ;
 wire \i_peripherals.i_user_peri39._GEN[103] ;
 wire \i_peripherals.i_user_peri39._GEN[104] ;
 wire \i_peripherals.i_user_peri39._GEN[105] ;
 wire \i_peripherals.i_user_peri39._GEN[106] ;
 wire \i_peripherals.i_user_peri39._GEN[107] ;
 wire \i_peripherals.i_user_peri39._GEN[108] ;
 wire \i_peripherals.i_user_peri39._GEN[109] ;
 wire \i_peripherals.i_user_peri39._GEN[110] ;
 wire \i_peripherals.i_user_peri39._GEN[111] ;
 wire \i_peripherals.i_user_peri39._GEN[112] ;
 wire \i_peripherals.i_user_peri39._GEN[113] ;
 wire \i_peripherals.i_user_peri39._GEN[114] ;
 wire \i_peripherals.i_user_peri39._GEN[115] ;
 wire \i_peripherals.i_user_peri39._GEN[116] ;
 wire \i_peripherals.i_user_peri39._GEN[117] ;
 wire \i_peripherals.i_user_peri39._GEN[118] ;
 wire \i_peripherals.i_user_peri39._GEN[119] ;
 wire \i_peripherals.i_user_peri39._GEN[120] ;
 wire \i_peripherals.i_user_peri39._GEN[121] ;
 wire \i_peripherals.i_user_peri39._GEN[122] ;
 wire \i_peripherals.i_user_peri39._GEN[123] ;
 wire \i_peripherals.i_user_peri39._GEN[124] ;
 wire \i_peripherals.i_user_peri39._GEN[125] ;
 wire \i_peripherals.i_user_peri39._GEN[126] ;
 wire \i_peripherals.i_user_peri39._GEN[127] ;
 wire \i_peripherals.i_user_peri39._GEN[1] ;
 wire \i_peripherals.i_user_peri39._GEN[2] ;
 wire \i_peripherals.i_user_peri39._GEN[32] ;
 wire \i_peripherals.i_user_peri39._GEN[33] ;
 wire \i_peripherals.i_user_peri39._GEN[34] ;
 wire \i_peripherals.i_user_peri39._GEN[35] ;
 wire \i_peripherals.i_user_peri39._GEN[36] ;
 wire \i_peripherals.i_user_peri39._GEN[37] ;
 wire \i_peripherals.i_user_peri39._GEN[38] ;
 wire \i_peripherals.i_user_peri39._GEN[39] ;
 wire \i_peripherals.i_user_peri39._GEN[3] ;
 wire \i_peripherals.i_user_peri39._GEN[40] ;
 wire \i_peripherals.i_user_peri39._GEN[41] ;
 wire \i_peripherals.i_user_peri39._GEN[42] ;
 wire \i_peripherals.i_user_peri39._GEN[43] ;
 wire \i_peripherals.i_user_peri39._GEN[44] ;
 wire \i_peripherals.i_user_peri39._GEN[45] ;
 wire \i_peripherals.i_user_peri39._GEN[46] ;
 wire \i_peripherals.i_user_peri39._GEN[47] ;
 wire \i_peripherals.i_user_peri39._GEN[48] ;
 wire \i_peripherals.i_user_peri39._GEN[49] ;
 wire \i_peripherals.i_user_peri39._GEN[50] ;
 wire \i_peripherals.i_user_peri39._GEN[51] ;
 wire \i_peripherals.i_user_peri39._GEN[52] ;
 wire \i_peripherals.i_user_peri39._GEN[53] ;
 wire \i_peripherals.i_user_peri39._GEN[54] ;
 wire \i_peripherals.i_user_peri39._GEN[55] ;
 wire \i_peripherals.i_user_peri39._GEN[56] ;
 wire \i_peripherals.i_user_peri39._GEN[57] ;
 wire \i_peripherals.i_user_peri39._GEN[58] ;
 wire \i_peripherals.i_user_peri39._GEN[59] ;
 wire \i_peripherals.i_user_peri39._GEN[60] ;
 wire \i_peripherals.i_user_peri39._GEN[61] ;
 wire \i_peripherals.i_user_peri39._GEN[62] ;
 wire \i_peripherals.i_user_peri39._GEN[63] ;
 wire \i_peripherals.i_user_peri39._GEN[64] ;
 wire \i_peripherals.i_user_peri39._GEN[65] ;
 wire \i_peripherals.i_user_peri39._GEN[66] ;
 wire \i_peripherals.i_user_peri39._GEN[67] ;
 wire \i_peripherals.i_user_peri39._GEN[68] ;
 wire \i_peripherals.i_user_peri39._GEN[69] ;
 wire \i_peripherals.i_user_peri39._GEN[70] ;
 wire \i_peripherals.i_user_peri39._GEN[71] ;
 wire \i_peripherals.i_user_peri39._GEN[72] ;
 wire \i_peripherals.i_user_peri39._GEN[73] ;
 wire \i_peripherals.i_user_peri39._GEN[74] ;
 wire \i_peripherals.i_user_peri39._GEN[75] ;
 wire \i_peripherals.i_user_peri39._GEN[76] ;
 wire \i_peripherals.i_user_peri39._GEN[77] ;
 wire \i_peripherals.i_user_peri39._GEN[78] ;
 wire \i_peripherals.i_user_peri39._GEN[79] ;
 wire \i_peripherals.i_user_peri39._GEN[80] ;
 wire \i_peripherals.i_user_peri39._GEN[81] ;
 wire \i_peripherals.i_user_peri39._GEN[82] ;
 wire \i_peripherals.i_user_peri39._GEN[83] ;
 wire \i_peripherals.i_user_peri39._GEN[84] ;
 wire \i_peripherals.i_user_peri39._GEN[85] ;
 wire \i_peripherals.i_user_peri39._GEN[86] ;
 wire \i_peripherals.i_user_peri39._GEN[87] ;
 wire \i_peripherals.i_user_peri39._GEN[88] ;
 wire \i_peripherals.i_user_peri39._GEN[89] ;
 wire \i_peripherals.i_user_peri39._GEN[90] ;
 wire \i_peripherals.i_user_peri39._GEN[91] ;
 wire \i_peripherals.i_user_peri39._GEN[92] ;
 wire \i_peripherals.i_user_peri39._GEN[93] ;
 wire \i_peripherals.i_user_peri39._GEN[94] ;
 wire \i_peripherals.i_user_peri39._GEN[95] ;
 wire \i_peripherals.i_user_peri39.busy_counter[0] ;
 wire \i_peripherals.i_user_peri39.busy_counter[1] ;
 wire \i_peripherals.i_user_peri39.busy_counter[2] ;
 wire \i_peripherals.i_user_peri39.instr[0] ;
 wire \i_peripherals.i_user_peri39.instr[10] ;
 wire \i_peripherals.i_user_peri39.instr[11] ;
 wire \i_peripherals.i_user_peri39.instr[12] ;
 wire \i_peripherals.i_user_peri39.instr[13] ;
 wire \i_peripherals.i_user_peri39.instr[14] ;
 wire \i_peripherals.i_user_peri39.instr[15] ;
 wire \i_peripherals.i_user_peri39.instr[16] ;
 wire \i_peripherals.i_user_peri39.instr[17] ;
 wire \i_peripherals.i_user_peri39.instr[18] ;
 wire \i_peripherals.i_user_peri39.instr[19] ;
 wire \i_peripherals.i_user_peri39.instr[1] ;
 wire \i_peripherals.i_user_peri39.instr[20] ;
 wire \i_peripherals.i_user_peri39.instr[21] ;
 wire \i_peripherals.i_user_peri39.instr[22] ;
 wire \i_peripherals.i_user_peri39.instr[23] ;
 wire \i_peripherals.i_user_peri39.instr[24] ;
 wire \i_peripherals.i_user_peri39.instr[25] ;
 wire \i_peripherals.i_user_peri39.instr[26] ;
 wire \i_peripherals.i_user_peri39.instr[27] ;
 wire \i_peripherals.i_user_peri39.instr[28] ;
 wire \i_peripherals.i_user_peri39.instr[29] ;
 wire \i_peripherals.i_user_peri39.instr[2] ;
 wire \i_peripherals.i_user_peri39.instr[30] ;
 wire \i_peripherals.i_user_peri39.instr[31] ;
 wire \i_peripherals.i_user_peri39.instr[3] ;
 wire \i_peripherals.i_user_peri39.instr[4] ;
 wire \i_peripherals.i_user_peri39.instr[5] ;
 wire \i_peripherals.i_user_peri39.instr[6] ;
 wire \i_peripherals.i_user_peri39.instr[7] ;
 wire \i_peripherals.i_user_peri39.instr[8] ;
 wire \i_peripherals.i_user_peri39.instr[9] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[0] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[10] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[11] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[12] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[13] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[14] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[15] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[16] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[17] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[18] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[19] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[1] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[20] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[21] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[22] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[23] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[24] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[25] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[26] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[27] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[28] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[29] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[2] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[30] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[31] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[3] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[4] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[5] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[6] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[7] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[8] ;
 wire \i_peripherals.i_user_peri39.math_result_reg[9] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[0] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[10] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[11] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[12] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[13] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[14] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[15] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[16] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[17] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[18] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[19] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[1] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[20] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[21] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[22] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[23] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[24] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[25] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[26] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[27] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[28] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[29] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[2] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[30] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[31] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[32] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[3] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[4] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[5] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[6] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[7] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[8] ;
 wire \i_peripherals.i_user_peri39.stage1_math_rec[9] ;
 wire \i_tinyqv.cpu.additional_mem_ops[0] ;
 wire \i_tinyqv.cpu.additional_mem_ops[1] ;
 wire \i_tinyqv.cpu.additional_mem_ops[2] ;
 wire \i_tinyqv.cpu.addr_offset[2] ;
 wire \i_tinyqv.cpu.addr_offset[3] ;
 wire \i_tinyqv.cpu.alu_op[0] ;
 wire \i_tinyqv.cpu.alu_op[1] ;
 wire \i_tinyqv.cpu.alu_op[2] ;
 wire \i_tinyqv.cpu.alu_op[3] ;
 wire \i_tinyqv.cpu.counter[2] ;
 wire \i_tinyqv.cpu.counter[3] ;
 wire \i_tinyqv.cpu.counter[4] ;
 wire \i_tinyqv.cpu.data_read_n[0] ;
 wire \i_tinyqv.cpu.data_read_n[1] ;
 wire \i_tinyqv.cpu.data_ready_latch ;
 wire \i_tinyqv.cpu.data_ready_sync ;
 wire \i_tinyqv.cpu.data_write_n[0] ;
 wire \i_tinyqv.cpu.data_write_n[1] ;
 wire \i_tinyqv.cpu.i_core.cmp ;
 wire \i_tinyqv.cpu.i_core.cmp_out ;
 wire \i_tinyqv.cpu.i_core.cy ;
 wire \i_tinyqv.cpu.i_core.cy_out ;
 wire \i_tinyqv.cpu.i_core.cycle[0] ;
 wire \i_tinyqv.cpu.i_core.cycle[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[0] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[1] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[2] ;
 wire \i_tinyqv.cpu.i_core.cycle_count[3] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[4] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[5] ;
 wire \i_tinyqv.cpu.i_core.cycle_count_wide[6] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.cy ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_cycles.rstn ;
 wire \i_tinyqv.cpu.i_core.i_instrret.add ;
 wire \i_tinyqv.cpu.i_core.i_instrret.cy ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[0] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[1] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[2] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.data[3] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rd[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs1[3] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[0] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[1] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[2] ;
 wire \i_tinyqv.cpu.i_core.i_registers.rs2[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[10] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[11] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[12] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[13] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[14] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[15] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[16] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[17] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[18] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[19] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[20] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[21] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[22] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[23] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[24] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[25] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[26] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[27] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[28] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[29] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[30] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[31] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[4] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[5] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[6] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[7] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[8] ;
 wire \i_tinyqv.cpu.i_core.i_shift.a[9] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ;
 wire \i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[2] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[3] ;
 wire \i_tinyqv.cpu.i_core.i_shift.b[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[0] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[10] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[11] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[1] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[2] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[3] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[4] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[5] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[6] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[7] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[8] ;
 wire \i_tinyqv.cpu.i_core.imm_lo[9] ;
 wire \i_tinyqv.cpu.i_core.is_double_fault_r ;
 wire \i_tinyqv.cpu.i_core.is_interrupt ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[0] ;
 wire \i_tinyqv.cpu.i_core.last_interrupt_req[1] ;
 wire \i_tinyqv.cpu.i_core.load_done ;
 wire \i_tinyqv.cpu.i_core.load_top_bit ;
 wire \i_tinyqv.cpu.i_core.mcause[0] ;
 wire \i_tinyqv.cpu.i_core.mcause[1] ;
 wire \i_tinyqv.cpu.i_core.mcause[2] ;
 wire \i_tinyqv.cpu.i_core.mcause[3] ;
 wire \i_tinyqv.cpu.i_core.mcause[4] ;
 wire \i_tinyqv.cpu.i_core.mcause[5] ;
 wire \i_tinyqv.cpu.i_core.mem_op[0] ;
 wire \i_tinyqv.cpu.i_core.mem_op[1] ;
 wire \i_tinyqv.cpu.i_core.mem_op[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[0] ;
 wire \i_tinyqv.cpu.i_core.mepc[10] ;
 wire \i_tinyqv.cpu.i_core.mepc[11] ;
 wire \i_tinyqv.cpu.i_core.mepc[12] ;
 wire \i_tinyqv.cpu.i_core.mepc[13] ;
 wire \i_tinyqv.cpu.i_core.mepc[14] ;
 wire \i_tinyqv.cpu.i_core.mepc[15] ;
 wire \i_tinyqv.cpu.i_core.mepc[16] ;
 wire \i_tinyqv.cpu.i_core.mepc[17] ;
 wire \i_tinyqv.cpu.i_core.mepc[18] ;
 wire \i_tinyqv.cpu.i_core.mepc[19] ;
 wire \i_tinyqv.cpu.i_core.mepc[1] ;
 wire \i_tinyqv.cpu.i_core.mepc[20] ;
 wire \i_tinyqv.cpu.i_core.mepc[21] ;
 wire \i_tinyqv.cpu.i_core.mepc[22] ;
 wire \i_tinyqv.cpu.i_core.mepc[23] ;
 wire \i_tinyqv.cpu.i_core.mepc[2] ;
 wire \i_tinyqv.cpu.i_core.mepc[3] ;
 wire \i_tinyqv.cpu.i_core.mepc[4] ;
 wire \i_tinyqv.cpu.i_core.mepc[5] ;
 wire \i_tinyqv.cpu.i_core.mepc[6] ;
 wire \i_tinyqv.cpu.i_core.mepc[7] ;
 wire \i_tinyqv.cpu.i_core.mepc[8] ;
 wire \i_tinyqv.cpu.i_core.mepc[9] ;
 wire \i_tinyqv.cpu.i_core.mie[0] ;
 wire \i_tinyqv.cpu.i_core.mie[10] ;
 wire \i_tinyqv.cpu.i_core.mie[11] ;
 wire \i_tinyqv.cpu.i_core.mie[12] ;
 wire \i_tinyqv.cpu.i_core.mie[13] ;
 wire \i_tinyqv.cpu.i_core.mie[14] ;
 wire \i_tinyqv.cpu.i_core.mie[15] ;
 wire \i_tinyqv.cpu.i_core.mie[16] ;
 wire \i_tinyqv.cpu.i_core.mie[1] ;
 wire \i_tinyqv.cpu.i_core.mie[2] ;
 wire \i_tinyqv.cpu.i_core.mie[3] ;
 wire \i_tinyqv.cpu.i_core.mie[4] ;
 wire \i_tinyqv.cpu.i_core.mie[5] ;
 wire \i_tinyqv.cpu.i_core.mie[6] ;
 wire \i_tinyqv.cpu.i_core.mie[7] ;
 wire \i_tinyqv.cpu.i_core.mie[8] ;
 wire \i_tinyqv.cpu.i_core.mie[9] ;
 wire \i_tinyqv.cpu.i_core.mip[0] ;
 wire \i_tinyqv.cpu.i_core.mip[16] ;
 wire \i_tinyqv.cpu.i_core.mip[1] ;
 wire \i_tinyqv.cpu.i_core.mstatus_mie ;
 wire \i_tinyqv.cpu.i_core.mstatus_mpie ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[0] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[10] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[11] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[12] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[13] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[14] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[15] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[1] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[2] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[3] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[4] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[5] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[6] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[7] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[8] ;
 wire \i_tinyqv.cpu.i_core.multiplier.accum[9] ;
 wire \i_tinyqv.cpu.i_core.time_hi[0] ;
 wire \i_tinyqv.cpu.i_core.time_hi[1] ;
 wire \i_tinyqv.cpu.i_core.time_hi[2] ;
 wire \i_tinyqv.cpu.i_timer.cy ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.cy ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.data[0] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.data[1] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.data[2] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.data[3] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[10] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[11] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[12] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[13] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[14] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[15] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[16] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[17] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[18] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[19] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[20] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[21] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[22] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[23] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[24] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[25] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[26] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[27] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[28] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[29] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[30] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[31] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[4] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[5] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[6] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[7] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[8] ;
 wire \i_tinyqv.cpu.i_timer.i_mtime.reg_buf[9] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[0] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[10] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[11] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[12] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[13] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[14] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[15] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[16] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[17] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[18] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[19] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[1] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[20] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[21] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[22] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[23] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[24] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[25] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[26] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[27] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[28] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[29] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[2] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[30] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[31] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[3] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[4] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[5] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[6] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[7] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[8] ;
 wire \i_tinyqv.cpu.i_timer.mtimecmp[9] ;
 wire \i_tinyqv.cpu.i_timer.time_pulse_r ;
 wire \i_tinyqv.cpu.imm[12] ;
 wire \i_tinyqv.cpu.imm[13] ;
 wire \i_tinyqv.cpu.imm[14] ;
 wire \i_tinyqv.cpu.imm[15] ;
 wire \i_tinyqv.cpu.imm[16] ;
 wire \i_tinyqv.cpu.imm[17] ;
 wire \i_tinyqv.cpu.imm[18] ;
 wire \i_tinyqv.cpu.imm[19] ;
 wire \i_tinyqv.cpu.imm[20] ;
 wire \i_tinyqv.cpu.imm[21] ;
 wire \i_tinyqv.cpu.imm[22] ;
 wire \i_tinyqv.cpu.imm[23] ;
 wire \i_tinyqv.cpu.imm[24] ;
 wire \i_tinyqv.cpu.imm[25] ;
 wire \i_tinyqv.cpu.imm[26] ;
 wire \i_tinyqv.cpu.imm[27] ;
 wire \i_tinyqv.cpu.imm[28] ;
 wire \i_tinyqv.cpu.imm[29] ;
 wire \i_tinyqv.cpu.imm[30] ;
 wire \i_tinyqv.cpu.imm[31] ;
 wire \i_tinyqv.cpu.instr_data[0][0] ;
 wire \i_tinyqv.cpu.instr_data[0][10] ;
 wire \i_tinyqv.cpu.instr_data[0][11] ;
 wire \i_tinyqv.cpu.instr_data[0][12] ;
 wire \i_tinyqv.cpu.instr_data[0][13] ;
 wire \i_tinyqv.cpu.instr_data[0][14] ;
 wire \i_tinyqv.cpu.instr_data[0][15] ;
 wire \i_tinyqv.cpu.instr_data[0][1] ;
 wire \i_tinyqv.cpu.instr_data[0][2] ;
 wire \i_tinyqv.cpu.instr_data[0][3] ;
 wire \i_tinyqv.cpu.instr_data[0][4] ;
 wire \i_tinyqv.cpu.instr_data[0][5] ;
 wire \i_tinyqv.cpu.instr_data[0][6] ;
 wire \i_tinyqv.cpu.instr_data[0][7] ;
 wire \i_tinyqv.cpu.instr_data[0][8] ;
 wire \i_tinyqv.cpu.instr_data[0][9] ;
 wire \i_tinyqv.cpu.instr_data[1][0] ;
 wire \i_tinyqv.cpu.instr_data[1][10] ;
 wire \i_tinyqv.cpu.instr_data[1][11] ;
 wire \i_tinyqv.cpu.instr_data[1][12] ;
 wire \i_tinyqv.cpu.instr_data[1][13] ;
 wire \i_tinyqv.cpu.instr_data[1][14] ;
 wire \i_tinyqv.cpu.instr_data[1][15] ;
 wire \i_tinyqv.cpu.instr_data[1][1] ;
 wire \i_tinyqv.cpu.instr_data[1][2] ;
 wire \i_tinyqv.cpu.instr_data[1][3] ;
 wire \i_tinyqv.cpu.instr_data[1][4] ;
 wire \i_tinyqv.cpu.instr_data[1][5] ;
 wire \i_tinyqv.cpu.instr_data[1][6] ;
 wire \i_tinyqv.cpu.instr_data[1][7] ;
 wire \i_tinyqv.cpu.instr_data[1][8] ;
 wire \i_tinyqv.cpu.instr_data[1][9] ;
 wire \i_tinyqv.cpu.instr_data[2][0] ;
 wire \i_tinyqv.cpu.instr_data[2][10] ;
 wire \i_tinyqv.cpu.instr_data[2][11] ;
 wire \i_tinyqv.cpu.instr_data[2][12] ;
 wire \i_tinyqv.cpu.instr_data[2][13] ;
 wire \i_tinyqv.cpu.instr_data[2][14] ;
 wire \i_tinyqv.cpu.instr_data[2][15] ;
 wire \i_tinyqv.cpu.instr_data[2][1] ;
 wire \i_tinyqv.cpu.instr_data[2][2] ;
 wire \i_tinyqv.cpu.instr_data[2][3] ;
 wire \i_tinyqv.cpu.instr_data[2][4] ;
 wire \i_tinyqv.cpu.instr_data[2][5] ;
 wire \i_tinyqv.cpu.instr_data[2][6] ;
 wire \i_tinyqv.cpu.instr_data[2][7] ;
 wire \i_tinyqv.cpu.instr_data[2][8] ;
 wire \i_tinyqv.cpu.instr_data[2][9] ;
 wire \i_tinyqv.cpu.instr_data[3][0] ;
 wire \i_tinyqv.cpu.instr_data[3][10] ;
 wire \i_tinyqv.cpu.instr_data[3][11] ;
 wire \i_tinyqv.cpu.instr_data[3][12] ;
 wire \i_tinyqv.cpu.instr_data[3][13] ;
 wire \i_tinyqv.cpu.instr_data[3][14] ;
 wire \i_tinyqv.cpu.instr_data[3][15] ;
 wire \i_tinyqv.cpu.instr_data[3][1] ;
 wire \i_tinyqv.cpu.instr_data[3][2] ;
 wire \i_tinyqv.cpu.instr_data[3][3] ;
 wire \i_tinyqv.cpu.instr_data[3][4] ;
 wire \i_tinyqv.cpu.instr_data[3][5] ;
 wire \i_tinyqv.cpu.instr_data[3][6] ;
 wire \i_tinyqv.cpu.instr_data[3][7] ;
 wire \i_tinyqv.cpu.instr_data[3][8] ;
 wire \i_tinyqv.cpu.instr_data[3][9] ;
 wire \i_tinyqv.cpu.instr_data_in[0] ;
 wire \i_tinyqv.cpu.instr_data_in[10] ;
 wire \i_tinyqv.cpu.instr_data_in[11] ;
 wire \i_tinyqv.cpu.instr_data_in[12] ;
 wire \i_tinyqv.cpu.instr_data_in[13] ;
 wire \i_tinyqv.cpu.instr_data_in[14] ;
 wire \i_tinyqv.cpu.instr_data_in[15] ;
 wire \i_tinyqv.cpu.instr_data_in[1] ;
 wire \i_tinyqv.cpu.instr_data_in[2] ;
 wire \i_tinyqv.cpu.instr_data_in[3] ;
 wire \i_tinyqv.cpu.instr_data_in[4] ;
 wire \i_tinyqv.cpu.instr_data_in[5] ;
 wire \i_tinyqv.cpu.instr_data_in[6] ;
 wire \i_tinyqv.cpu.instr_data_in[7] ;
 wire \i_tinyqv.cpu.instr_data_in[8] ;
 wire \i_tinyqv.cpu.instr_data_in[9] ;
 wire \i_tinyqv.cpu.instr_data_start[10] ;
 wire \i_tinyqv.cpu.instr_data_start[11] ;
 wire \i_tinyqv.cpu.instr_data_start[12] ;
 wire \i_tinyqv.cpu.instr_data_start[13] ;
 wire \i_tinyqv.cpu.instr_data_start[14] ;
 wire \i_tinyqv.cpu.instr_data_start[15] ;
 wire \i_tinyqv.cpu.instr_data_start[16] ;
 wire \i_tinyqv.cpu.instr_data_start[17] ;
 wire \i_tinyqv.cpu.instr_data_start[18] ;
 wire \i_tinyqv.cpu.instr_data_start[19] ;
 wire \i_tinyqv.cpu.instr_data_start[20] ;
 wire \i_tinyqv.cpu.instr_data_start[21] ;
 wire \i_tinyqv.cpu.instr_data_start[22] ;
 wire \i_tinyqv.cpu.instr_data_start[23] ;
 wire \i_tinyqv.cpu.instr_data_start[3] ;
 wire \i_tinyqv.cpu.instr_data_start[4] ;
 wire \i_tinyqv.cpu.instr_data_start[5] ;
 wire \i_tinyqv.cpu.instr_data_start[6] ;
 wire \i_tinyqv.cpu.instr_data_start[7] ;
 wire \i_tinyqv.cpu.instr_data_start[8] ;
 wire \i_tinyqv.cpu.instr_data_start[9] ;
 wire \i_tinyqv.cpu.instr_fetch_running ;
 wire \i_tinyqv.cpu.instr_fetch_started ;
 wire \i_tinyqv.cpu.instr_fetch_stopped ;
 wire \i_tinyqv.cpu.instr_len[1] ;
 wire \i_tinyqv.cpu.instr_len[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[1] ;
 wire \i_tinyqv.cpu.instr_write_offset[2] ;
 wire \i_tinyqv.cpu.instr_write_offset[3] ;
 wire \i_tinyqv.cpu.is_alu_imm ;
 wire \i_tinyqv.cpu.is_alu_reg ;
 wire \i_tinyqv.cpu.is_auipc ;
 wire \i_tinyqv.cpu.is_branch ;
 wire \i_tinyqv.cpu.is_jal ;
 wire \i_tinyqv.cpu.is_jalr ;
 wire \i_tinyqv.cpu.is_load ;
 wire \i_tinyqv.cpu.is_lui ;
 wire \i_tinyqv.cpu.is_store ;
 wire \i_tinyqv.cpu.is_system ;
 wire \i_tinyqv.cpu.load_started ;
 wire \i_tinyqv.cpu.mem_op_increment_reg ;
 wire \i_tinyqv.cpu.no_write_in_progress ;
 wire \i_tinyqv.cpu.pc[1] ;
 wire \i_tinyqv.cpu.pc[2] ;
 wire \i_tinyqv.cpu.was_early_branch ;
 wire \i_tinyqv.mem.continue_txn ;
 wire \i_tinyqv.mem.data_from_read[16] ;
 wire \i_tinyqv.mem.data_from_read[17] ;
 wire \i_tinyqv.mem.data_from_read[18] ;
 wire \i_tinyqv.mem.data_from_read[19] ;
 wire \i_tinyqv.mem.data_from_read[20] ;
 wire \i_tinyqv.mem.data_from_read[21] ;
 wire \i_tinyqv.mem.data_from_read[22] ;
 wire \i_tinyqv.mem.data_from_read[23] ;
 wire \i_tinyqv.mem.data_stall ;
 wire \i_tinyqv.mem.data_txn_len[0] ;
 wire \i_tinyqv.mem.data_txn_len[1] ;
 wire \i_tinyqv.mem.instr_active ;
 wire \i_tinyqv.mem.q_ctrl.addr[0] ;
 wire \i_tinyqv.mem.q_ctrl.addr[10] ;
 wire \i_tinyqv.mem.q_ctrl.addr[11] ;
 wire \i_tinyqv.mem.q_ctrl.addr[12] ;
 wire \i_tinyqv.mem.q_ctrl.addr[13] ;
 wire \i_tinyqv.mem.q_ctrl.addr[14] ;
 wire \i_tinyqv.mem.q_ctrl.addr[15] ;
 wire \i_tinyqv.mem.q_ctrl.addr[16] ;
 wire \i_tinyqv.mem.q_ctrl.addr[17] ;
 wire \i_tinyqv.mem.q_ctrl.addr[18] ;
 wire \i_tinyqv.mem.q_ctrl.addr[19] ;
 wire \i_tinyqv.mem.q_ctrl.addr[1] ;
 wire \i_tinyqv.mem.q_ctrl.addr[20] ;
 wire \i_tinyqv.mem.q_ctrl.addr[21] ;
 wire \i_tinyqv.mem.q_ctrl.addr[22] ;
 wire \i_tinyqv.mem.q_ctrl.addr[23] ;
 wire \i_tinyqv.mem.q_ctrl.addr[2] ;
 wire \i_tinyqv.mem.q_ctrl.addr[3] ;
 wire \i_tinyqv.mem.q_ctrl.addr[4] ;
 wire \i_tinyqv.mem.q_ctrl.addr[5] ;
 wire \i_tinyqv.mem.q_ctrl.addr[6] ;
 wire \i_tinyqv.mem.q_ctrl.addr[7] ;
 wire \i_tinyqv.mem.q_ctrl.addr[8] ;
 wire \i_tinyqv.mem.q_ctrl.addr[9] ;
 wire \i_tinyqv.mem.q_ctrl.data_ready ;
 wire \i_tinyqv.mem.q_ctrl.data_req ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ;
 wire \i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[0] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[1] ;
 wire \i_tinyqv.mem.q_ctrl.fsm_state[2] ;
 wire \i_tinyqv.mem.q_ctrl.is_writing ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_a_sel ;
 wire \i_tinyqv.mem.q_ctrl.last_ram_b_sel ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ;
 wire \i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[0] ;
 wire \i_tinyqv.mem.q_ctrl.read_cycles_count[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_neg ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_out ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_pos ;
 wire \i_tinyqv.mem.q_ctrl.spi_clk_use_neg ;
 wire \i_tinyqv.mem.q_ctrl.spi_data_oe[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_flash_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ;
 wire \i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_a_select ;
 wire \i_tinyqv.mem.q_ctrl.spi_ram_b_select ;
 wire \i_tinyqv.mem.q_ctrl.stop_txn_reg ;
 wire \i_tinyqv.mem.qspi_data_buf[10] ;
 wire \i_tinyqv.mem.qspi_data_buf[11] ;
 wire \i_tinyqv.mem.qspi_data_buf[12] ;
 wire \i_tinyqv.mem.qspi_data_buf[13] ;
 wire \i_tinyqv.mem.qspi_data_buf[14] ;
 wire \i_tinyqv.mem.qspi_data_buf[15] ;
 wire \i_tinyqv.mem.qspi_data_buf[24] ;
 wire \i_tinyqv.mem.qspi_data_buf[25] ;
 wire \i_tinyqv.mem.qspi_data_buf[26] ;
 wire \i_tinyqv.mem.qspi_data_buf[27] ;
 wire \i_tinyqv.mem.qspi_data_buf[28] ;
 wire \i_tinyqv.mem.qspi_data_buf[29] ;
 wire \i_tinyqv.mem.qspi_data_buf[30] ;
 wire \i_tinyqv.mem.qspi_data_buf[31] ;
 wire \i_tinyqv.mem.qspi_data_buf[8] ;
 wire \i_tinyqv.mem.qspi_data_buf[9] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[0] ;
 wire \i_tinyqv.mem.qspi_data_byte_idx[1] ;
 wire \i_tinyqv.mem.qspi_write_done ;
 wire \time_count[0] ;
 wire \time_count[1] ;
 wire \time_count[2] ;
 wire \time_count[3] ;
 wire \time_count[4] ;
 wire \time_count[5] ;
 wire \time_count[6] ;
 wire \time_limit[2] ;
 wire \time_limit[3] ;
 wire \time_limit[4] ;
 wire \time_limit[5] ;
 wire \time_limit[6] ;
 wire \ui_in_sync0[0] ;
 wire \ui_in_sync0[1] ;
 wire \ui_in_sync0[2] ;
 wire \ui_in_sync0[3] ;
 wire \ui_in_sync0[4] ;
 wire \ui_in_sync0[5] ;
 wire \ui_in_sync0[6] ;
 wire \ui_in_sync0[7] ;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire clknet_leaf_0_clk_regs;
 wire clknet_leaf_1_clk_regs;
 wire clknet_leaf_2_clk_regs;
 wire clknet_leaf_3_clk_regs;
 wire clknet_leaf_4_clk_regs;
 wire clknet_leaf_5_clk_regs;
 wire clknet_leaf_6_clk_regs;
 wire clknet_leaf_7_clk_regs;
 wire clknet_leaf_8_clk_regs;
 wire clknet_leaf_9_clk_regs;
 wire clknet_leaf_10_clk_regs;
 wire clknet_leaf_11_clk_regs;
 wire clknet_leaf_12_clk_regs;
 wire clknet_leaf_13_clk_regs;
 wire clknet_leaf_14_clk_regs;
 wire clknet_leaf_15_clk_regs;
 wire clknet_leaf_16_clk_regs;
 wire clknet_leaf_17_clk_regs;
 wire clknet_leaf_18_clk_regs;
 wire clknet_leaf_19_clk_regs;
 wire clknet_leaf_20_clk_regs;
 wire clknet_leaf_21_clk_regs;
 wire clknet_leaf_22_clk_regs;
 wire clknet_leaf_23_clk_regs;
 wire clknet_leaf_24_clk_regs;
 wire clknet_leaf_25_clk_regs;
 wire clknet_leaf_26_clk_regs;
 wire clknet_leaf_27_clk_regs;
 wire clknet_leaf_28_clk_regs;
 wire clknet_leaf_29_clk_regs;
 wire clknet_leaf_30_clk_regs;
 wire clknet_leaf_31_clk_regs;
 wire clknet_leaf_32_clk_regs;
 wire clknet_leaf_33_clk_regs;
 wire clknet_leaf_34_clk_regs;
 wire clknet_leaf_35_clk_regs;
 wire clknet_leaf_36_clk_regs;
 wire clknet_leaf_37_clk_regs;
 wire clknet_leaf_38_clk_regs;
 wire clknet_leaf_39_clk_regs;
 wire clknet_leaf_40_clk_regs;
 wire clknet_leaf_41_clk_regs;
 wire clknet_leaf_42_clk_regs;
 wire clknet_leaf_43_clk_regs;
 wire clknet_leaf_44_clk_regs;
 wire clknet_leaf_45_clk_regs;
 wire clknet_leaf_46_clk_regs;
 wire clknet_leaf_47_clk_regs;
 wire clknet_leaf_48_clk_regs;
 wire clknet_leaf_49_clk_regs;
 wire clknet_leaf_50_clk_regs;
 wire clknet_leaf_51_clk_regs;
 wire clknet_leaf_52_clk_regs;
 wire clknet_leaf_53_clk_regs;
 wire clknet_leaf_54_clk_regs;
 wire clknet_leaf_55_clk_regs;
 wire clknet_leaf_56_clk_regs;
 wire clknet_leaf_57_clk_regs;
 wire clknet_leaf_58_clk_regs;
 wire clknet_leaf_59_clk_regs;
 wire clknet_leaf_60_clk_regs;
 wire clknet_leaf_61_clk_regs;
 wire clknet_leaf_62_clk_regs;
 wire clknet_leaf_63_clk_regs;
 wire clknet_leaf_64_clk_regs;
 wire clknet_leaf_65_clk_regs;
 wire clknet_leaf_66_clk_regs;
 wire clknet_leaf_67_clk_regs;
 wire clknet_leaf_68_clk_regs;
 wire clknet_leaf_69_clk_regs;
 wire clknet_leaf_70_clk_regs;
 wire clknet_leaf_71_clk_regs;
 wire clknet_leaf_72_clk_regs;
 wire clknet_leaf_73_clk_regs;
 wire clknet_leaf_74_clk_regs;
 wire clknet_leaf_75_clk_regs;
 wire clknet_leaf_76_clk_regs;
 wire clknet_leaf_77_clk_regs;
 wire clknet_leaf_78_clk_regs;
 wire clknet_leaf_79_clk_regs;
 wire clknet_leaf_80_clk_regs;
 wire clknet_leaf_81_clk_regs;
 wire clknet_leaf_82_clk_regs;
 wire clknet_leaf_83_clk_regs;
 wire clknet_leaf_84_clk_regs;
 wire clknet_leaf_85_clk_regs;
 wire clknet_leaf_86_clk_regs;
 wire clknet_leaf_87_clk_regs;
 wire clknet_leaf_88_clk_regs;
 wire clknet_leaf_89_clk_regs;
 wire clknet_leaf_90_clk_regs;
 wire clknet_leaf_91_clk_regs;
 wire clknet_leaf_92_clk_regs;
 wire clknet_leaf_93_clk_regs;
 wire clknet_leaf_94_clk_regs;
 wire clknet_leaf_95_clk_regs;
 wire clknet_leaf_96_clk_regs;
 wire clknet_leaf_97_clk_regs;
 wire clknet_leaf_98_clk_regs;
 wire clknet_leaf_99_clk_regs;
 wire clknet_leaf_100_clk_regs;
 wire clknet_leaf_101_clk_regs;
 wire clknet_leaf_102_clk_regs;
 wire clknet_leaf_103_clk_regs;
 wire clknet_leaf_104_clk_regs;
 wire clknet_leaf_105_clk_regs;
 wire clknet_leaf_106_clk_regs;
 wire clknet_leaf_107_clk_regs;
 wire clknet_leaf_108_clk_regs;
 wire clknet_leaf_109_clk_regs;
 wire clknet_leaf_110_clk_regs;
 wire clknet_leaf_111_clk_regs;
 wire clknet_leaf_112_clk_regs;
 wire clknet_leaf_113_clk_regs;
 wire clknet_leaf_114_clk_regs;
 wire clknet_leaf_115_clk_regs;
 wire clknet_leaf_116_clk_regs;
 wire clknet_leaf_117_clk_regs;
 wire clknet_leaf_118_clk_regs;
 wire clknet_leaf_119_clk_regs;
 wire clknet_leaf_120_clk_regs;
 wire clknet_leaf_121_clk_regs;
 wire clknet_leaf_122_clk_regs;
 wire clknet_leaf_123_clk_regs;
 wire clknet_leaf_124_clk_regs;
 wire clknet_leaf_125_clk_regs;
 wire clknet_leaf_126_clk_regs;
 wire clknet_leaf_127_clk_regs;
 wire clknet_leaf_128_clk_regs;
 wire clknet_leaf_129_clk_regs;
 wire clknet_leaf_130_clk_regs;
 wire clknet_leaf_131_clk_regs;
 wire clknet_leaf_132_clk_regs;
 wire clknet_leaf_133_clk_regs;
 wire clknet_leaf_134_clk_regs;
 wire clknet_leaf_135_clk_regs;
 wire clknet_leaf_136_clk_regs;
 wire clknet_leaf_137_clk_regs;
 wire clknet_leaf_138_clk_regs;
 wire clknet_leaf_139_clk_regs;
 wire clknet_leaf_140_clk_regs;
 wire clknet_leaf_141_clk_regs;
 wire clknet_leaf_142_clk_regs;
 wire clknet_leaf_143_clk_regs;
 wire clknet_leaf_144_clk_regs;
 wire clknet_leaf_145_clk_regs;
 wire clknet_leaf_146_clk_regs;
 wire clknet_leaf_147_clk_regs;
 wire clknet_leaf_148_clk_regs;
 wire clknet_leaf_149_clk_regs;
 wire clknet_leaf_150_clk_regs;
 wire clknet_leaf_151_clk_regs;
 wire clknet_leaf_152_clk_regs;
 wire clknet_leaf_153_clk_regs;
 wire clknet_leaf_154_clk_regs;
 wire clknet_leaf_155_clk_regs;
 wire clknet_leaf_156_clk_regs;
 wire clknet_leaf_157_clk_regs;
 wire clknet_leaf_158_clk_regs;
 wire clknet_leaf_159_clk_regs;
 wire clknet_leaf_160_clk_regs;
 wire clknet_leaf_161_clk_regs;
 wire clknet_leaf_162_clk_regs;
 wire clknet_leaf_163_clk_regs;
 wire clknet_leaf_164_clk_regs;
 wire clknet_leaf_165_clk_regs;
 wire clknet_leaf_166_clk_regs;
 wire clknet_leaf_167_clk_regs;
 wire clknet_leaf_168_clk_regs;
 wire clknet_leaf_169_clk_regs;
 wire clknet_leaf_170_clk_regs;
 wire clknet_leaf_171_clk_regs;
 wire clknet_leaf_172_clk_regs;
 wire clknet_leaf_173_clk_regs;
 wire clknet_leaf_174_clk_regs;
 wire clknet_leaf_175_clk_regs;
 wire clknet_leaf_176_clk_regs;
 wire clknet_leaf_177_clk_regs;
 wire clknet_0_clk_regs;
 wire clknet_3_0_0_clk_regs;
 wire clknet_3_1_0_clk_regs;
 wire clknet_3_2_0_clk_regs;
 wire clknet_3_3_0_clk_regs;
 wire clknet_3_4_0_clk_regs;
 wire clknet_3_5_0_clk_regs;
 wire clknet_3_6_0_clk_regs;
 wire clknet_3_7_0_clk_regs;
 wire clknet_5_0__leaf_clk_regs;
 wire clknet_5_1__leaf_clk_regs;
 wire clknet_5_2__leaf_clk_regs;
 wire clknet_5_3__leaf_clk_regs;
 wire clknet_5_4__leaf_clk_regs;
 wire clknet_5_5__leaf_clk_regs;
 wire clknet_5_6__leaf_clk_regs;
 wire clknet_5_7__leaf_clk_regs;
 wire clknet_5_8__leaf_clk_regs;
 wire clknet_5_9__leaf_clk_regs;
 wire clknet_5_10__leaf_clk_regs;
 wire clknet_5_11__leaf_clk_regs;
 wire clknet_5_12__leaf_clk_regs;
 wire clknet_5_13__leaf_clk_regs;
 wire clknet_5_14__leaf_clk_regs;
 wire clknet_5_15__leaf_clk_regs;
 wire clknet_5_16__leaf_clk_regs;
 wire clknet_5_17__leaf_clk_regs;
 wire clknet_5_18__leaf_clk_regs;
 wire clknet_5_19__leaf_clk_regs;
 wire clknet_5_20__leaf_clk_regs;
 wire clknet_5_21__leaf_clk_regs;
 wire clknet_5_22__leaf_clk_regs;
 wire clknet_5_23__leaf_clk_regs;
 wire clknet_5_24__leaf_clk_regs;
 wire clknet_5_25__leaf_clk_regs;
 wire clknet_5_26__leaf_clk_regs;
 wire clknet_5_27__leaf_clk_regs;
 wire clknet_5_28__leaf_clk_regs;
 wire clknet_5_29__leaf_clk_regs;
 wire clknet_5_30__leaf_clk_regs;
 wire clknet_5_31__leaf_clk_regs;
 wire delaynet_0_clk;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire net3649;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3653;
 wire net3654;
 wire net3655;
 wire net3656;
 wire net3657;
 wire net3658;
 wire net3659;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3668;
 wire net3669;
 wire net3670;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3677;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3688;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3702;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3725;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3782;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3808;
 wire net3809;
 wire net3810;
 wire net3811;
 wire net3812;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3821;
 wire net3822;
 wire net3823;
 wire net3824;
 wire net3825;
 wire net3826;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3848;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3858;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3869;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3878;
 wire net3879;
 wire net3880;
 wire net3881;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3889;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3901;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3911;
 wire net3912;
 wire net3913;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3920;
 wire net3921;
 wire net3922;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3927;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3931;
 wire net3932;
 wire net3933;
 wire net3934;
 wire net3935;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3939;
 wire net3940;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3953;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3965;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3973;
 wire net3974;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3979;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3983;
 wire net3984;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3988;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net3992;
 wire net3993;
 wire net3994;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net3999;
 wire net4000;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4004;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4008;
 wire net4009;
 wire net4010;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4016;
 wire net4017;
 wire net4018;
 wire net4019;
 wire net4020;
 wire net4021;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4028;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4037;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4041;
 wire net4042;
 wire net4043;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4052;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4061;
 wire net4062;
 wire net4063;
 wire net4064;
 wire net4065;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4069;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4075;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4084;
 wire net4085;
 wire net4086;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4106;
 wire net4107;
 wire net4108;
 wire net4109;
 wire net4110;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4114;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4122;
 wire net4123;
 wire net4124;
 wire net4125;
 wire net4126;
 wire net4127;
 wire net4128;
 wire net4129;
 wire net4130;
 wire net4131;
 wire net4132;
 wire net4133;
 wire net4134;
 wire net4135;
 wire net4136;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4143;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4147;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4157;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4161;
 wire net4162;
 wire net4163;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;

 sg13g2_inv_4 _08658_ (.A(net2358),
    .Y(_00923_));
 sg13g2_inv_2 _08659_ (.Y(_00924_),
    .A(net2362));
 sg13g2_inv_1 _08660_ (.Y(_00925_),
    .A(net3767));
 sg13g2_inv_1 _08661_ (.Y(_00926_),
    .A(\i_tinyqv.cpu.is_jalr ));
 sg13g2_inv_1 _08662_ (.Y(_00927_),
    .A(net3652));
 sg13g2_inv_2 _08663_ (.Y(_00928_),
    .A(net3444));
 sg13g2_inv_1 _08664_ (.Y(_00929_),
    .A(net3043));
 sg13g2_inv_1 _08665_ (.Y(_00930_),
    .A(net3154));
 sg13g2_inv_1 _08666_ (.Y(_00931_),
    .A(net3309));
 sg13g2_inv_1 _08667_ (.Y(_00932_),
    .A(net3197));
 sg13g2_inv_1 _08668_ (.Y(_00933_),
    .A(net3168));
 sg13g2_inv_1 _08669_ (.Y(_00934_),
    .A(net3219));
 sg13g2_inv_1 _08670_ (.Y(_00935_),
    .A(net3095));
 sg13g2_inv_1 _08671_ (.Y(_00936_),
    .A(net3237));
 sg13g2_inv_1 _08672_ (.Y(_00937_),
    .A(net3172));
 sg13g2_inv_1 _08673_ (.Y(_00938_),
    .A(net3176));
 sg13g2_inv_1 _08674_ (.Y(_00939_),
    .A(net2991));
 sg13g2_inv_1 _08675_ (.Y(_00940_),
    .A(net3376));
 sg13g2_inv_2 _08676_ (.Y(_00941_),
    .A(net3827));
 sg13g2_inv_1 _08677_ (.Y(_00942_),
    .A(net3666));
 sg13g2_inv_1 _08678_ (.Y(_00943_),
    .A(\addr[5] ));
 sg13g2_inv_1 _08679_ (.Y(_00944_),
    .A(net3163));
 sg13g2_inv_1 _08680_ (.Y(_00945_),
    .A(net2775));
 sg13g2_inv_1 _08681_ (.Y(_00946_),
    .A(net4154));
 sg13g2_inv_1 _08682_ (.Y(_00947_),
    .A(\i_tinyqv.cpu.data_write_n[1] ));
 sg13g2_inv_4 _08683_ (.A(net3281),
    .Y(_00948_));
 sg13g2_inv_4 _08684_ (.A(net3327),
    .Y(_00949_));
 sg13g2_inv_4 _08685_ (.A(net3317),
    .Y(_00950_));
 sg13g2_inv_4 _08686_ (.A(net3229),
    .Y(_00951_));
 sg13g2_inv_4 _08687_ (.A(net3386),
    .Y(_00952_));
 sg13g2_inv_4 _08688_ (.A(net3329),
    .Y(_00953_));
 sg13g2_inv_4 _08689_ (.A(net3196),
    .Y(_00954_));
 sg13g2_inv_4 _08690_ (.A(net3225),
    .Y(_00955_));
 sg13g2_inv_4 _08691_ (.A(net3591),
    .Y(_00956_));
 sg13g2_inv_4 _08692_ (.A(net3643),
    .Y(_00957_));
 sg13g2_inv_4 _08693_ (.A(net3642),
    .Y(_00958_));
 sg13g2_inv_4 _08694_ (.A(net3772),
    .Y(_00959_));
 sg13g2_inv_4 _08695_ (.A(net3607),
    .Y(_00960_));
 sg13g2_inv_4 _08696_ (.A(net3480),
    .Y(_00961_));
 sg13g2_inv_4 _08697_ (.A(net3674),
    .Y(_00962_));
 sg13g2_inv_4 _08698_ (.A(net3435),
    .Y(_00963_));
 sg13g2_inv_4 _08699_ (.A(\data_to_write[14] ),
    .Y(_00964_));
 sg13g2_inv_4 _08700_ (.A(net3590),
    .Y(_00965_));
 sg13g2_inv_2 _08701_ (.Y(_00966_),
    .A(\data_to_write[9] ));
 sg13g2_inv_2 _08702_ (.Y(_00967_),
    .A(\data_to_write[7] ));
 sg13g2_inv_8 _08703_ (.Y(_00968_),
    .A(net4082));
 sg13g2_inv_4 _08704_ (.A(net2389),
    .Y(_00969_));
 sg13g2_inv_4 _08705_ (.A(net2392),
    .Y(_00970_));
 sg13g2_inv_8 _08706_ (.Y(_00971_),
    .A(net2393));
 sg13g2_inv_8 _08707_ (.Y(_00972_),
    .A(net2396));
 sg13g2_inv_8 _08708_ (.Y(_00973_),
    .A(net2397));
 sg13g2_inv_4 _08709_ (.A(net2399),
    .Y(_00974_));
 sg13g2_inv_2 _08710_ (.Y(_00975_),
    .A(net3963));
 sg13g2_inv_2 _08711_ (.Y(_00976_),
    .A(net3972));
 sg13g2_inv_1 _08712_ (.Y(_00977_),
    .A(net4070));
 sg13g2_inv_4 _08713_ (.A(net3820),
    .Y(_00978_));
 sg13g2_inv_2 _08714_ (.Y(_00979_),
    .A(\i_tinyqv.cpu.instr_data_start[12] ));
 sg13g2_inv_2 _08715_ (.Y(_00980_),
    .A(\i_tinyqv.cpu.instr_data_start[9] ));
 sg13g2_inv_2 _08716_ (.Y(_00981_),
    .A(net4063));
 sg13g2_inv_1 _08717_ (.Y(_00982_),
    .A(net4077));
 sg13g2_inv_2 _08718_ (.Y(_00983_),
    .A(net2437));
 sg13g2_inv_1 _08719_ (.Y(_00984_),
    .A(net3707));
 sg13g2_inv_2 _08720_ (.Y(_00985_),
    .A(net4028));
 sg13g2_inv_2 _08721_ (.Y(_00986_),
    .A(net3784));
 sg13g2_inv_1 _08722_ (.Y(_00987_),
    .A(net3892));
 sg13g2_inv_2 _08723_ (.Y(_00988_),
    .A(net3727));
 sg13g2_inv_1 _08724_ (.Y(_00989_),
    .A(\i_peripherals.i_uart.baud_divider[9] ));
 sg13g2_inv_2 _08725_ (.Y(_00990_),
    .A(net3690));
 sg13g2_inv_1 _08726_ (.Y(_00991_),
    .A(net2783));
 sg13g2_inv_1 _08727_ (.Y(_00992_),
    .A(net2920));
 sg13g2_inv_1 _08728_ (.Y(_00993_),
    .A(net2796));
 sg13g2_inv_1 _08729_ (.Y(_00994_),
    .A(net2845));
 sg13g2_inv_1 _08730_ (.Y(_00995_),
    .A(net3074));
 sg13g2_inv_1 _08731_ (.Y(_00996_),
    .A(net2763));
 sg13g2_inv_1 _08732_ (.Y(_00997_),
    .A(net2890));
 sg13g2_inv_1 _08733_ (.Y(_00998_),
    .A(net2821));
 sg13g2_inv_1 _08734_ (.Y(_00999_),
    .A(net3065));
 sg13g2_inv_1 _08735_ (.Y(_01000_),
    .A(net2753));
 sg13g2_inv_1 _08736_ (.Y(_01001_),
    .A(net2755));
 sg13g2_inv_1 _08737_ (.Y(_01002_),
    .A(net2803));
 sg13g2_inv_1 _08738_ (.Y(_01003_),
    .A(net2761));
 sg13g2_inv_1 _08739_ (.Y(_01004_),
    .A(net2915));
 sg13g2_inv_1 _08740_ (.Y(_01005_),
    .A(net2759));
 sg13g2_inv_1 _08741_ (.Y(_01006_),
    .A(net2767));
 sg13g2_inv_1 _08742_ (.Y(_01007_),
    .A(net3024));
 sg13g2_inv_1 _08743_ (.Y(_01008_),
    .A(net2846));
 sg13g2_inv_1 _08744_ (.Y(_01009_),
    .A(net2815));
 sg13g2_inv_1 _08745_ (.Y(_01010_),
    .A(net2748));
 sg13g2_inv_1 _08746_ (.Y(_01011_),
    .A(net2765));
 sg13g2_inv_1 _08747_ (.Y(_01012_),
    .A(net2888));
 sg13g2_inv_1 _08748_ (.Y(_01013_),
    .A(net2790));
 sg13g2_inv_1 _08749_ (.Y(_01014_),
    .A(net2869));
 sg13g2_inv_1 _08750_ (.Y(_01015_),
    .A(net2777));
 sg13g2_inv_1 _08751_ (.Y(_01016_),
    .A(net2824));
 sg13g2_inv_1 _08752_ (.Y(_01017_),
    .A(net2948));
 sg13g2_inv_1 _08753_ (.Y(_01018_),
    .A(net2757));
 sg13g2_inv_1 _08754_ (.Y(_01019_),
    .A(net3102));
 sg13g2_inv_1 _08755_ (.Y(_01020_),
    .A(\i_tinyqv.cpu.i_core.mie[4] ));
 sg13g2_inv_1 _08756_ (.Y(_01021_),
    .A(\i_tinyqv.cpu.i_core.mie[7] ));
 sg13g2_inv_1 _08757_ (.Y(_01022_),
    .A(net3182));
 sg13g2_inv_1 _08758_ (.Y(_01023_),
    .A(net3988));
 sg13g2_inv_1 _08759_ (.Y(_01024_),
    .A(\i_debug_uart_tx.cycle_counter[3] ));
 sg13g2_inv_1 _08760_ (.Y(_01025_),
    .A(net2773));
 sg13g2_inv_1 _08761_ (.Y(_01026_),
    .A(net2892));
 sg13g2_inv_1 _08762_ (.Y(_01027_),
    .A(net2769));
 sg13g2_inv_1 _08763_ (.Y(_01028_),
    .A(net3091));
 sg13g2_inv_1 _08764_ (.Y(_01029_),
    .A(net2941));
 sg13g2_inv_1 _08765_ (.Y(_01030_),
    .A(net2946));
 sg13g2_inv_1 _08766_ (.Y(_01031_),
    .A(net3187));
 sg13g2_inv_1 _08767_ (.Y(_01032_),
    .A(net3264));
 sg13g2_inv_1 _08768_ (.Y(_01033_),
    .A(net3136));
 sg13g2_inv_1 _08769_ (.Y(_01034_),
    .A(net3266));
 sg13g2_inv_1 _08770_ (.Y(_01035_),
    .A(net3093));
 sg13g2_inv_1 _08771_ (.Y(_01036_),
    .A(net2966));
 sg13g2_inv_1 _08772_ (.Y(_01037_),
    .A(net3054));
 sg13g2_inv_1 _08773_ (.Y(_01038_),
    .A(net2884));
 sg13g2_inv_2 _08774_ (.Y(_01039_),
    .A(net3758));
 sg13g2_inv_1 _08775_ (.Y(_01040_),
    .A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[12] ));
 sg13g2_inv_1 _08776_ (.Y(_01041_),
    .A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[11] ));
 sg13g2_inv_1 _08777_ (.Y(_01042_),
    .A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[4] ));
 sg13g2_inv_1 _08778_ (.Y(_01043_),
    .A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[3] ));
 sg13g2_inv_1 _08779_ (.Y(_01044_),
    .A(net3337));
 sg13g2_inv_2 _08780_ (.Y(_01045_),
    .A(net3216));
 sg13g2_inv_1 _08781_ (.Y(_01046_),
    .A(net3063));
 sg13g2_inv_2 _08782_ (.Y(_01047_),
    .A(net3921));
 sg13g2_inv_2 _08783_ (.Y(_01048_),
    .A(net4015));
 sg13g2_inv_2 _08784_ (.Y(_01049_),
    .A(\i_peripherals.i_uart.baud_divider[5] ));
 sg13g2_inv_1 _08785_ (.Y(_01050_),
    .A(net3986));
 sg13g2_inv_1 _08786_ (.Y(_01051_),
    .A(\i_peripherals.i_uart.baud_divider[3] ));
 sg13g2_inv_2 _08787_ (.Y(_01052_),
    .A(net3877));
 sg13g2_inv_2 _08788_ (.Y(_01053_),
    .A(\i_peripherals.i_uart.baud_divider[1] ));
 sg13g2_inv_1 _08789_ (.Y(_01054_),
    .A(net3702));
 sg13g2_inv_1 _08790_ (.Y(_01055_),
    .A(net3022));
 sg13g2_inv_1 _08791_ (.Y(_01056_),
    .A(net3747));
 sg13g2_inv_1 _08792_ (.Y(_01057_),
    .A(\i_peripherals.i_user_peri39.instr[15] ));
 sg13g2_inv_1 _08793_ (.Y(_01058_),
    .A(net2805));
 sg13g2_inv_1 _08794_ (.Y(_01059_),
    .A(net2779));
 sg13g2_inv_1 _08795_ (.Y(_01060_),
    .A(net2751));
 sg13g2_inv_1 _08796_ (.Y(_01061_),
    .A(net3463));
 sg13g2_inv_1 _08797_ (.Y(_01062_),
    .A(net2771));
 sg13g2_inv_1 _08798_ (.Y(_01063_),
    .A(net3003));
 sg13g2_inv_1 _08799_ (.Y(_01064_),
    .A(net2835));
 sg13g2_inv_1 _08800_ (.Y(_01065_),
    .A(net2492));
 sg13g2_inv_1 _08801_ (.Y(_01066_),
    .A(net2997));
 sg13g2_inv_1 _08802_ (.Y(_01067_),
    .A(net2378));
 sg13g2_inv_2 _08803_ (.Y(_01068_),
    .A(net3995));
 sg13g2_inv_1 _08804_ (.Y(_01069_),
    .A(net3621));
 sg13g2_inv_1 _08805_ (.Y(_01070_),
    .A(net3887));
 sg13g2_inv_1 _08806_ (.Y(_01071_),
    .A(net3788));
 sg13g2_inv_2 _08807_ (.Y(_01072_),
    .A(net3965));
 sg13g2_inv_1 _08808_ (.Y(_01073_),
    .A(\i_tinyqv.cpu.imm[12] ));
 sg13g2_inv_1 _08809_ (.Y(_01074_),
    .A(net3961));
 sg13g2_inv_1 _08810_ (.Y(_01075_),
    .A(net2906));
 sg13g2_inv_2 _08811_ (.Y(_01076_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ));
 sg13g2_inv_2 _08812_ (.Y(_01077_),
    .A(\i_tinyqv.cpu.instr_write_offset[1] ));
 sg13g2_inv_2 _08813_ (.Y(_01078_),
    .A(net2435));
 sg13g2_inv_1 _08814_ (.Y(_01079_),
    .A(\i_peripherals.i_user_peri39._GEN[79] ));
 sg13g2_inv_1 _08815_ (.Y(_01080_),
    .A(\i_peripherals.i_user_peri39._GEN[83] ));
 sg13g2_inv_1 _08816_ (.Y(_01081_),
    .A(\i_peripherals.i_user_peri39._GEN[91] ));
 sg13g2_inv_1 _08817_ (.Y(_01082_),
    .A(\i_peripherals.i_user_peri39._GEN[89] ));
 sg13g2_inv_1 _08818_ (.Y(_01083_),
    .A(\i_peripherals.i_user_peri39._GEN[90] ));
 sg13g2_inv_1 _08819_ (.Y(_01084_),
    .A(\i_peripherals.i_user_peri39._GEN[92] ));
 sg13g2_inv_1 _08820_ (.Y(_01085_),
    .A(\i_peripherals.i_user_peri39._GEN[93] ));
 sg13g2_inv_1 _08821_ (.Y(_01086_),
    .A(\i_peripherals.i_user_peri39._GEN[94] ));
 sg13g2_inv_1 _08822_ (.Y(_01087_),
    .A(net2870));
 sg13g2_inv_1 _08823_ (.Y(_01088_),
    .A(net2929));
 sg13g2_inv_1 _08824_ (.Y(_01089_),
    .A(net3166));
 sg13g2_inv_1 _08825_ (.Y(_01090_),
    .A(\i_tinyqv.cpu.instr_data[2][0] ));
 sg13g2_inv_1 _08826_ (.Y(_01091_),
    .A(net2907));
 sg13g2_inv_1 _08827_ (.Y(_01092_),
    .A(net2943));
 sg13g2_inv_1 _08828_ (.Y(_01093_),
    .A(net2989));
 sg13g2_inv_1 _08829_ (.Y(_01094_),
    .A(\i_tinyqv.cpu.instr_data[2][1] ));
 sg13g2_inv_1 _08830_ (.Y(_01095_),
    .A(net4088));
 sg13g2_inv_1 _08831_ (.Y(_01096_),
    .A(net3232));
 sg13g2_inv_1 _08832_ (.Y(_01097_),
    .A(net3516));
 sg13g2_inv_1 _08833_ (.Y(_01098_),
    .A(net2265));
 sg13g2_inv_1 _08834_ (.Y(_01099_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[2] ));
 sg13g2_inv_1 _08835_ (.Y(_01100_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[3] ));
 sg13g2_inv_1 _08836_ (.Y(_01101_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[4] ));
 sg13g2_inv_1 _08837_ (.Y(_01102_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[6] ));
 sg13g2_inv_1 _08838_ (.Y(_01103_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[9] ));
 sg13g2_inv_1 _08839_ (.Y(_01104_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[10] ));
 sg13g2_inv_1 _08840_ (.Y(_01105_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[11] ));
 sg13g2_inv_1 _08841_ (.Y(_01106_),
    .A(net4037));
 sg13g2_inv_2 _08842_ (.Y(_01107_),
    .A(net3983));
 sg13g2_inv_1 _08843_ (.Y(_01108_),
    .A(net4020));
 sg13g2_inv_2 _08844_ (.Y(_01109_),
    .A(net4091));
 sg13g2_inv_1 _08845_ (.Y(_01110_),
    .A(\i_tinyqv.cpu.instr_fetch_stopped ));
 sg13g2_inv_1 _08846_ (.Y(_01111_),
    .A(\i_tinyqv.cpu.i_timer.mtimecmp[5] ));
 sg13g2_inv_1 _08847_ (.Y(_01112_),
    .A(\i_tinyqv.cpu.i_timer.i_mtime.data[1] ));
 sg13g2_inv_1 _08848_ (.Y(_01113_),
    .A(\i_tinyqv.cpu.i_timer.i_mtime.data[0] ));
 sg13g2_inv_1 _08849_ (.Y(_01114_),
    .A(\i_tinyqv.cpu.i_timer.cy ));
 sg13g2_inv_1 _08850_ (.Y(_01115_),
    .A(net4033));
 sg13g2_inv_1 _08851_ (.Y(_01116_),
    .A(net4045));
 sg13g2_inv_2 _08852_ (.Y(_01117_),
    .A(\i_tinyqv.cpu.instr_data_in[0] ));
 sg13g2_inv_4 _08853_ (.A(net3045),
    .Y(_01118_));
 sg13g2_inv_2 _08854_ (.Y(_01119_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[28] ));
 sg13g2_inv_1 _08855_ (.Y(_01120_),
    .A(net2476));
 sg13g2_inv_1 _08856_ (.Y(_01121_),
    .A(net2468));
 sg13g2_inv_1 _08857_ (.Y(_01122_),
    .A(net3311));
 sg13g2_inv_1 _08858_ (.Y(_01123_),
    .A(\i_tinyqv.cpu.instr_data_in[1] ));
 sg13g2_inv_8 _08859_ (.Y(_01124_),
    .A(\i_tinyqv.cpu.instr_data_in[9] ));
 sg13g2_inv_4 _08860_ (.A(net4099),
    .Y(_01125_));
 sg13g2_inv_1 _08861_ (.Y(_01126_),
    .A(\i_tinyqv.mem.qspi_data_buf[9] ));
 sg13g2_inv_1 _08862_ (.Y(_01127_),
    .A(net3087));
 sg13g2_inv_1 _08863_ (.Y(_01128_),
    .A(net4134));
 sg13g2_inv_8 _08864_ (.Y(_01129_),
    .A(net3996));
 sg13g2_inv_1 _08865_ (.Y(_01130_),
    .A(\i_tinyqv.mem.qspi_data_buf[10] ));
 sg13g2_inv_1 _08866_ (.Y(_01131_),
    .A(\i_tinyqv.mem.data_from_read[18] ));
 sg13g2_inv_1 _08867_ (.Y(_01132_),
    .A(net3254));
 sg13g2_inv_8 _08868_ (.Y(_01133_),
    .A(\i_tinyqv.cpu.instr_data_in[11] ));
 sg13g2_inv_4 _08869_ (.A(net3932),
    .Y(_01134_));
 sg13g2_inv_1 _08870_ (.Y(_01135_),
    .A(net2787));
 sg13g2_inv_1 _08871_ (.Y(_01136_),
    .A(\i_tinyqv.mem.qspi_data_buf[15] ));
 sg13g2_inv_1 _08872_ (.Y(_01137_),
    .A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ));
 sg13g2_inv_1 _08873_ (.Y(_01138_),
    .A(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ));
 sg13g2_inv_1 _08874_ (.Y(_01139_),
    .A(net3841));
 sg13g2_inv_1 _08875_ (.Y(_01140_),
    .A(net2451));
 sg13g2_inv_1 _08876_ (.Y(_01141_),
    .A(net3871));
 sg13g2_inv_4 _08877_ (.A(net2443),
    .Y(_01142_));
 sg13g2_inv_1 _08878_ (.Y(_01143_),
    .A(net3803));
 sg13g2_inv_2 _08879_ (.Y(_01144_),
    .A(net3759));
 sg13g2_inv_1 _08880_ (.Y(_01145_),
    .A(net3470));
 sg13g2_inv_1 _08881_ (.Y(_01146_),
    .A(net3395));
 sg13g2_inv_1 _08882_ (.Y(_01147_),
    .A(net3328));
 sg13g2_inv_1 _08883_ (.Y(_01148_),
    .A(net3416));
 sg13g2_inv_2 _08884_ (.Y(_01149_),
    .A(\i_peripherals.i_uart.i_uart_tx.txd_reg ));
 sg13g2_inv_1 _08885_ (.Y(_01150_),
    .A(net6));
 sg13g2_inv_1 _08886_ (.Y(_01151_),
    .A(net7));
 sg13g2_inv_1 _08887_ (.Y(_01152_),
    .A(net3099));
 sg13g2_inv_1 _08888_ (.Y(_01153_),
    .A(net3174));
 sg13g2_inv_1 _08889_ (.Y(_01154_),
    .A(net2809));
 sg13g2_inv_1 _08890_ (.Y(_01155_),
    .A(net2916));
 sg13g2_inv_1 _08891_ (.Y(_01156_),
    .A(net2685));
 sg13g2_inv_1 _15914__2 (.Y(net1435),
    .A(clknet_1_0__leaf_clk));
 sg13g2_nand2b_2 _08893_ (.Y(_01157_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ));
 sg13g2_nor3_2 _08894_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .C(_01157_),
    .Y(_01158_));
 sg13g2_nand2b_2 _08895_ (.Y(_01159_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ));
 sg13g2_nand2_2 _08896_ (.Y(_01160_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ));
 sg13g2_nor2_2 _08897_ (.A(_01159_),
    .B(_01160_),
    .Y(_01161_));
 sg13g2_nor2b_1 _08898_ (.A(net2384),
    .B_N(net2379),
    .Y(_01162_));
 sg13g2_nand2b_1 _08899_ (.Y(_01163_),
    .B(net2379),
    .A_N(net2382));
 sg13g2_nor2_2 _08900_ (.A(net2337),
    .B(net2324),
    .Y(_01164_));
 sg13g2_nor3_1 _08901_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .C(_01159_),
    .Y(_01165_));
 sg13g2_nand2b_2 _08902_ (.Y(_01166_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ));
 sg13g2_nor2_2 _08903_ (.A(_01159_),
    .B(_01166_),
    .Y(_01167_));
 sg13g2_nor2_2 _08904_ (.A(_01157_),
    .B(_01159_),
    .Y(_01168_));
 sg13g2_nand2_2 _08905_ (.Y(_01169_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_nor2_2 _08906_ (.A(_01166_),
    .B(_01169_),
    .Y(_01170_));
 sg13g2_nor3_2 _08907_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .C(_01166_),
    .Y(_01171_));
 sg13g2_nand2b_2 _08908_ (.Y(_01172_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ));
 sg13g2_nor2_2 _08909_ (.A(_01157_),
    .B(_01172_),
    .Y(_01173_));
 sg13g2_nor2_2 _08910_ (.A(_01166_),
    .B(_01172_),
    .Y(_01174_));
 sg13g2_nor2_2 _08911_ (.A(_01157_),
    .B(_01169_),
    .Y(_01175_));
 sg13g2_nor3_2 _08912_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .C(_01169_),
    .Y(_01176_));
 sg13g2_nor2_2 _08913_ (.A(_01160_),
    .B(_01169_),
    .Y(_01177_));
 sg13g2_nor3_2 _08914_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .C(_01172_),
    .Y(_01178_));
 sg13g2_nor2_2 _08915_ (.A(_01160_),
    .B(_01172_),
    .Y(_01179_));
 sg13g2_a22oi_1 _08916_ (.Y(_01180_),
    .B1(_01178_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .A2(_01171_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ));
 sg13g2_a22oi_1 _08917_ (.Y(_01181_),
    .B1(_01176_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .A2(_01174_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ));
 sg13g2_a22oi_1 _08918_ (.Y(_01182_),
    .B1(_01179_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .A2(_01168_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ));
 sg13g2_a22oi_1 _08919_ (.Y(_01183_),
    .B1(_01177_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .A2(_01170_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ));
 sg13g2_nand4_1 _08920_ (.B(_01181_),
    .C(_01182_),
    .A(_01180_),
    .Y(_01184_),
    .D(_01183_));
 sg13g2_a22oi_1 _08921_ (.Y(_01185_),
    .B1(_01164_),
    .B2(_01165_),
    .A2(_01158_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_a22oi_1 _08922_ (.Y(_01186_),
    .B1(_01175_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .A2(_01167_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ));
 sg13g2_a22oi_1 _08923_ (.Y(_01187_),
    .B1(_01173_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .A2(_01161_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_nand3_1 _08924_ (.B(_01186_),
    .C(_01187_),
    .A(_01185_),
    .Y(_01188_));
 sg13g2_or2_1 _08925_ (.X(_01189_),
    .B(_01188_),
    .A(_01184_));
 sg13g2_inv_2 _08926_ (.Y(_01190_),
    .A(_01189_));
 sg13g2_nand2_1 _08927_ (.Y(_01191_),
    .A(net2355),
    .B(\i_tinyqv.cpu.is_auipc ));
 sg13g2_o21ai_1 _08928_ (.B1(net2355),
    .Y(_01192_),
    .A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_auipc ));
 sg13g2_nand2_2 _08929_ (.Y(_01193_),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .B(net2371));
 sg13g2_nor2_2 _08930_ (.A(net2354),
    .B(_01193_),
    .Y(_01194_));
 sg13g2_nand3_1 _08931_ (.B(net2369),
    .C(net2371),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .Y(_01195_));
 sg13g2_nor2b_1 _08932_ (.A(net2379),
    .B_N(net2382),
    .Y(_01196_));
 sg13g2_nand2b_1 _08933_ (.Y(_01197_),
    .B(net2384),
    .A_N(net2379));
 sg13g2_nor2_1 _08934_ (.A(net2382),
    .B(net2379),
    .Y(_01198_));
 sg13g2_or2_1 _08935_ (.X(_01199_),
    .B(net2380),
    .A(net2384));
 sg13g2_a22oi_1 _08936_ (.Y(_01200_),
    .B1(net2313),
    .B2(net2418),
    .A2(net2318),
    .A1(net2416));
 sg13g2_and2_1 _08937_ (.A(net2382),
    .B(net2379),
    .X(_01201_));
 sg13g2_nand2_1 _08938_ (.Y(_01202_),
    .A(net2382),
    .B(net2380));
 sg13g2_a22oi_1 _08939_ (.Y(_01203_),
    .B1(net2309),
    .B2(\i_tinyqv.cpu.instr_data_start[15] ),
    .A2(net2326),
    .A1(\i_tinyqv.cpu.instr_data_start[11] ));
 sg13g2_a21oi_1 _08940_ (.A1(_01200_),
    .A2(_01203_),
    .Y(_01204_),
    .B1(net2375));
 sg13g2_nor2_2 _08941_ (.A(net2381),
    .B(net2336),
    .Y(_01205_));
 sg13g2_nor2_2 _08942_ (.A(net2337),
    .B(net2317),
    .Y(_01206_));
 sg13g2_nand2_2 _08943_ (.Y(_01207_),
    .A(net2375),
    .B(net2318));
 sg13g2_nor2_2 _08944_ (.A(net2336),
    .B(_01199_),
    .Y(_01208_));
 sg13g2_a22oi_1 _08945_ (.Y(_01209_),
    .B1(net2243),
    .B2(net2410),
    .A2(net2244),
    .A1(\i_tinyqv.cpu.instr_data_start[23] ));
 sg13g2_nand2b_1 _08946_ (.Y(_01210_),
    .B(_01209_),
    .A_N(_01204_));
 sg13g2_o21ai_1 _08947_ (.B1(net2323),
    .Y(_01211_),
    .A1(_01192_),
    .A2(_01210_));
 sg13g2_a21o_2 _08948_ (.A2(_01192_),
    .A1(_01190_),
    .B1(_01211_),
    .X(_01212_));
 sg13g2_nand2_1 _08949_ (.Y(_01213_),
    .A(net2371),
    .B(net2323));
 sg13g2_o21ai_1 _08950_ (.B1(net2323),
    .Y(_01214_),
    .A1(\i_tinyqv.cpu.alu_op[3] ),
    .A2(net2371));
 sg13g2_nor2_1 _08951_ (.A(_00923_),
    .B(_00927_),
    .Y(_01215_));
 sg13g2_nand2_2 _08952_ (.Y(_01216_),
    .A(net2356),
    .B(\i_tinyqv.cpu.is_branch ));
 sg13g2_o21ai_1 _08953_ (.B1(net2355),
    .Y(_01217_),
    .A1(\i_tinyqv.cpu.is_branch ),
    .A2(\i_tinyqv.cpu.is_alu_reg ));
 sg13g2_and2_1 _08954_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(net2314),
    .X(_01218_));
 sg13g2_a21oi_1 _08955_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .A2(net2320),
    .Y(_01219_),
    .B1(net2376));
 sg13g2_a221oi_1 _08956_ (.B2(\i_tinyqv.cpu.imm[15] ),
    .C1(_01218_),
    .B1(net2308),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .Y(_01220_),
    .A2(net2325));
 sg13g2_a22oi_1 _08957_ (.Y(_01221_),
    .B1(net2314),
    .B2(\i_tinyqv.cpu.imm[19] ),
    .A2(net2325),
    .A1(\i_tinyqv.cpu.imm[27] ));
 sg13g2_a221oi_1 _08958_ (.B2(\i_tinyqv.cpu.imm[31] ),
    .C1(net2338),
    .B1(net2308),
    .A1(\i_tinyqv.cpu.imm[23] ),
    .Y(_01222_),
    .A2(net2320));
 sg13g2_a22oi_1 _08959_ (.Y(_01223_),
    .B1(_01221_),
    .B2(_01222_),
    .A2(_01220_),
    .A1(_01219_));
 sg13g2_nand2_1 _08960_ (.Y(_01224_),
    .A(_01217_),
    .B(_01223_));
 sg13g2_nand2b_2 _08961_ (.Y(_01225_),
    .B(net2361),
    .A_N(net2360));
 sg13g2_nand2_2 _08962_ (.Y(_01226_),
    .A(net2359),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ));
 sg13g2_nor2_2 _08963_ (.A(_01225_),
    .B(_01226_),
    .Y(_01227_));
 sg13g2_nand2b_2 _08964_ (.Y(_01228_),
    .B(net2359),
    .A_N(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ));
 sg13g2_nand2b_2 _08965_ (.Y(_01229_),
    .B(net2360),
    .A_N(net2361));
 sg13g2_nor2_2 _08966_ (.A(_01228_),
    .B(_01229_),
    .Y(_01230_));
 sg13g2_a22oi_1 _08967_ (.Y(_01231_),
    .B1(_01230_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .A2(_01227_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ));
 sg13g2_nand2_2 _08968_ (.Y(_01232_),
    .A(net2360),
    .B(net2361));
 sg13g2_nand2b_2 _08969_ (.Y(_01233_),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .A_N(net2359));
 sg13g2_nor2_2 _08970_ (.A(_01232_),
    .B(_01233_),
    .Y(_01234_));
 sg13g2_nor3_2 _08971_ (.A(net2359),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .C(_01225_),
    .Y(_01235_));
 sg13g2_nor2_2 _08972_ (.A(_01226_),
    .B(_01229_),
    .Y(_01236_));
 sg13g2_nor2_2 _08973_ (.A(_01226_),
    .B(_01232_),
    .Y(_01237_));
 sg13g2_a22oi_1 _08974_ (.Y(_01238_),
    .B1(_01237_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .A2(_01236_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ));
 sg13g2_nor3_2 _08975_ (.A(net2359),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .C(_01229_),
    .Y(_01239_));
 sg13g2_nor3_2 _08976_ (.A(net2360),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .C(_01226_),
    .Y(_01240_));
 sg13g2_nor2_2 _08977_ (.A(_01229_),
    .B(_01233_),
    .Y(_01241_));
 sg13g2_nor2_2 _08978_ (.A(_01225_),
    .B(_01228_),
    .Y(_01242_));
 sg13g2_nor2_2 _08979_ (.A(_01225_),
    .B(_01233_),
    .Y(_01243_));
 sg13g2_nor2_2 _08980_ (.A(_01228_),
    .B(_01232_),
    .Y(_01244_));
 sg13g2_nor3_2 _08981_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .C(_01233_),
    .Y(_01245_));
 sg13g2_a22oi_1 _08982_ (.Y(_01246_),
    .B1(_01245_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .A2(_01240_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ));
 sg13g2_a22oi_1 _08983_ (.Y(_01247_),
    .B1(_01243_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .A2(_01234_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ));
 sg13g2_nor3_1 _08984_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .C(_01228_),
    .Y(_01248_));
 sg13g2_a22oi_1 _08985_ (.Y(_01249_),
    .B1(_01248_),
    .B2(_01164_),
    .A2(_01244_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ));
 sg13g2_a22oi_1 _08986_ (.Y(_01250_),
    .B1(_01241_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .A2(_01239_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ));
 sg13g2_nand4_1 _08987_ (.B(_01247_),
    .C(_01249_),
    .A(_01231_),
    .Y(_01251_),
    .D(_01250_));
 sg13g2_a22oi_1 _08988_ (.Y(_01252_),
    .B1(_01242_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .A2(_01235_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ));
 sg13g2_nand3_1 _08989_ (.B(_01246_),
    .C(_01252_),
    .A(_01238_),
    .Y(_01253_));
 sg13g2_nor2_2 _08990_ (.A(_01251_),
    .B(_01253_),
    .Y(_01254_));
 sg13g2_o21ai_1 _08991_ (.B1(_01224_),
    .Y(_01255_),
    .A1(_01217_),
    .A2(_01254_));
 sg13g2_inv_1 _08992_ (.Y(_01256_),
    .A(_01255_));
 sg13g2_xor2_1 _08993_ (.B(_01255_),
    .A(_01214_),
    .X(_01257_));
 sg13g2_a22oi_1 _08994_ (.Y(_01258_),
    .B1(_01175_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A2(_01161_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ));
 sg13g2_a22oi_1 _08995_ (.Y(_01259_),
    .B1(_01177_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .A2(_01158_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ));
 sg13g2_a22oi_1 _08996_ (.Y(_01260_),
    .B1(_01178_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A2(_01176_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ));
 sg13g2_nand3_1 _08997_ (.B(_01259_),
    .C(_01260_),
    .A(_01258_),
    .Y(_01261_));
 sg13g2_a22oi_1 _08998_ (.Y(_01262_),
    .B1(_01173_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .A2(_01171_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_a22oi_1 _08999_ (.Y(_01263_),
    .B1(_01179_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .A2(_01170_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_nor3_1 _09000_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .C(_01160_),
    .Y(_01264_));
 sg13g2_nor2_2 _09001_ (.A(net2376),
    .B(net2324),
    .Y(_01265_));
 sg13g2_a22oi_1 _09002_ (.Y(_01266_),
    .B1(_01264_),
    .B2(_01265_),
    .A2(_01168_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_a22oi_1 _09003_ (.Y(_01267_),
    .B1(_01174_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A2(_01167_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ));
 sg13g2_nand4_1 _09004_ (.B(_01263_),
    .C(_01266_),
    .A(_01262_),
    .Y(_01268_),
    .D(_01267_));
 sg13g2_nor2_2 _09005_ (.A(_01261_),
    .B(_01268_),
    .Y(_01269_));
 sg13g2_a22oi_1 _09006_ (.Y(_01270_),
    .B1(net2313),
    .B2(\i_tinyqv.cpu.pc[2] ),
    .A2(net2318),
    .A1(\i_tinyqv.cpu.instr_data_start[6] ));
 sg13g2_a22oi_1 _09007_ (.Y(_01271_),
    .B1(net2309),
    .B2(net2413),
    .A2(net2326),
    .A1(net2415));
 sg13g2_a21oi_1 _09008_ (.A1(_01270_),
    .A2(_01271_),
    .Y(_01272_),
    .B1(net2375));
 sg13g2_a22oi_1 _09009_ (.Y(_01273_),
    .B1(net2243),
    .B2(\i_tinyqv.cpu.instr_data_start[18] ),
    .A2(net2244),
    .A1(\i_tinyqv.cpu.instr_data_start[22] ));
 sg13g2_nand2b_1 _09010_ (.Y(_01274_),
    .B(_01273_),
    .A_N(_01272_));
 sg13g2_o21ai_1 _09011_ (.B1(net2323),
    .Y(_01275_),
    .A1(_01192_),
    .A2(_01274_));
 sg13g2_a21oi_2 _09012_ (.B1(_01275_),
    .Y(_01276_),
    .A2(_01269_),
    .A1(_01192_));
 sg13g2_a22oi_1 _09013_ (.Y(_01277_),
    .B1(net2308),
    .B2(\i_tinyqv.cpu.imm[30] ),
    .A2(net2313),
    .A1(\i_tinyqv.cpu.imm[18] ));
 sg13g2_a221oi_1 _09014_ (.B2(\i_tinyqv.cpu.imm[22] ),
    .C1(net2338),
    .B1(net2320),
    .A1(\i_tinyqv.cpu.imm[26] ),
    .Y(_01278_),
    .A2(net2325));
 sg13g2_a21oi_1 _09015_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .A2(net2313),
    .Y(_01279_),
    .B1(net2376));
 sg13g2_and2_1 _09016_ (.A(\i_tinyqv.cpu.imm[14] ),
    .B(net2308),
    .X(_01280_));
 sg13g2_a221oi_1 _09017_ (.B2(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .C1(_01280_),
    .B1(net2320),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .Y(_01281_),
    .A2(net2325));
 sg13g2_a22oi_1 _09018_ (.Y(_01282_),
    .B1(_01279_),
    .B2(_01281_),
    .A2(_01278_),
    .A1(_01277_));
 sg13g2_nor3_1 _09019_ (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .B(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .C(_01232_),
    .Y(_01283_));
 sg13g2_a22oi_1 _09020_ (.Y(_01284_),
    .B1(_01244_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .A2(_01227_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ));
 sg13g2_a22oi_1 _09021_ (.Y(_01285_),
    .B1(_01243_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .A2(_01230_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ));
 sg13g2_a22oi_1 _09022_ (.Y(_01286_),
    .B1(_01245_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .A2(_01241_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ));
 sg13g2_a22oi_1 _09023_ (.Y(_01287_),
    .B1(_01240_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .A2(_01237_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ));
 sg13g2_nand3_1 _09024_ (.B(_01286_),
    .C(_01287_),
    .A(_01285_),
    .Y(_01288_));
 sg13g2_a221oi_1 _09025_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .C1(_01288_),
    .B1(_01242_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .Y(_01289_),
    .A2(_01239_));
 sg13g2_a22oi_1 _09026_ (.Y(_01290_),
    .B1(_01265_),
    .B2(_01283_),
    .A2(_01234_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ));
 sg13g2_a22oi_1 _09027_ (.Y(_01291_),
    .B1(_01236_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .A2(_01235_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ));
 sg13g2_nand4_1 _09028_ (.B(_01289_),
    .C(_01290_),
    .A(_01284_),
    .Y(_01292_),
    .D(_01291_));
 sg13g2_mux2_1 _09029_ (.A0(_01292_),
    .A1(_01282_),
    .S(_01217_),
    .X(_01293_));
 sg13g2_xor2_1 _09030_ (.B(_01293_),
    .A(_01214_),
    .X(_01294_));
 sg13g2_inv_1 _09031_ (.Y(_01295_),
    .A(_01294_));
 sg13g2_nand2_1 _09032_ (.Y(_01296_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .B(_01158_));
 sg13g2_a22oi_1 _09033_ (.Y(_01297_),
    .B1(_01178_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A2(_01167_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ));
 sg13g2_a22oi_1 _09034_ (.Y(_01298_),
    .B1(_01179_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A2(_01171_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_a22oi_1 _09035_ (.Y(_01299_),
    .B1(_01168_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .A2(_01161_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ));
 sg13g2_a22oi_1 _09036_ (.Y(_01300_),
    .B1(_01176_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .A2(_01170_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ));
 sg13g2_nand3_1 _09037_ (.B(_01299_),
    .C(_01300_),
    .A(_01298_),
    .Y(_01301_));
 sg13g2_a22oi_1 _09038_ (.Y(_01302_),
    .B1(_01177_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .A2(_01173_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ));
 sg13g2_a22oi_1 _09039_ (.Y(_01303_),
    .B1(_01175_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A2(_01174_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ));
 sg13g2_nand4_1 _09040_ (.B(_01297_),
    .C(_01302_),
    .A(_01296_),
    .Y(_01304_),
    .D(_01303_));
 sg13g2_or2_1 _09041_ (.X(_01305_),
    .B(_01304_),
    .A(_01301_));
 sg13g2_a22oi_1 _09042_ (.Y(_01306_),
    .B1(net2313),
    .B2(\i_tinyqv.cpu.pc[1] ),
    .A2(net2319),
    .A1(\i_tinyqv.cpu.instr_data_start[5] ));
 sg13g2_a22oi_1 _09043_ (.Y(_01307_),
    .B1(net2309),
    .B2(\i_tinyqv.cpu.instr_data_start[13] ),
    .A2(net2326),
    .A1(\i_tinyqv.cpu.instr_data_start[9] ));
 sg13g2_nand2_1 _09044_ (.Y(_01308_),
    .A(_01306_),
    .B(_01307_));
 sg13g2_a22oi_1 _09045_ (.Y(_01309_),
    .B1(_01308_),
    .B2(net2336),
    .A2(net2243),
    .A1(net2411));
 sg13g2_o21ai_1 _09046_ (.B1(_01309_),
    .Y(_01310_),
    .A1(_00976_),
    .A2(_01207_));
 sg13g2_mux2_1 _09047_ (.A0(_01310_),
    .A1(_01305_),
    .S(_01192_),
    .X(_01311_));
 sg13g2_nand2_2 _09048_ (.Y(_01312_),
    .A(net2323),
    .B(_01311_));
 sg13g2_a22oi_1 _09049_ (.Y(_01313_),
    .B1(net2314),
    .B2(\i_tinyqv.cpu.imm[17] ),
    .A2(net2325),
    .A1(\i_tinyqv.cpu.imm[25] ));
 sg13g2_a221oi_1 _09050_ (.B2(\i_tinyqv.cpu.imm[29] ),
    .C1(net2338),
    .B1(net2308),
    .A1(\i_tinyqv.cpu.imm[21] ),
    .Y(_01314_),
    .A2(net2320));
 sg13g2_and2_1 _09051_ (.A(net2439),
    .B(net2315),
    .X(_01315_));
 sg13g2_a21oi_1 _09052_ (.A1(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .A2(net2325),
    .Y(_01316_),
    .B1(net2376));
 sg13g2_a221oi_1 _09053_ (.B2(\i_tinyqv.cpu.imm[13] ),
    .C1(_01315_),
    .B1(net2308),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .Y(_01317_),
    .A2(net2320));
 sg13g2_a22oi_1 _09054_ (.Y(_01318_),
    .B1(_01316_),
    .B2(_01317_),
    .A2(_01314_),
    .A1(_01313_));
 sg13g2_nand2_1 _09055_ (.Y(_01319_),
    .A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .B(_01230_));
 sg13g2_a22oi_1 _09056_ (.Y(_01320_),
    .B1(_01234_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .A2(_01227_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ));
 sg13g2_a22oi_1 _09057_ (.Y(_01321_),
    .B1(_01241_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .A2(_01237_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ));
 sg13g2_a22oi_1 _09058_ (.Y(_01322_),
    .B1(_01243_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .A2(_01240_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ));
 sg13g2_a22oi_1 _09059_ (.Y(_01323_),
    .B1(_01236_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .A2(_01235_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ));
 sg13g2_nand3_1 _09060_ (.B(_01322_),
    .C(_01323_),
    .A(_01320_),
    .Y(_01324_));
 sg13g2_a22oi_1 _09061_ (.Y(_01325_),
    .B1(_01244_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .A2(_01242_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ));
 sg13g2_a22oi_1 _09062_ (.Y(_01326_),
    .B1(_01245_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .A2(_01239_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ));
 sg13g2_nand4_1 _09063_ (.B(_01321_),
    .C(_01325_),
    .A(_01319_),
    .Y(_01327_),
    .D(_01326_));
 sg13g2_nor2_2 _09064_ (.A(_01324_),
    .B(_01327_),
    .Y(_01328_));
 sg13g2_nor2_1 _09065_ (.A(_01217_),
    .B(_01328_),
    .Y(_01329_));
 sg13g2_a21oi_2 _09066_ (.B1(_01329_),
    .Y(_01330_),
    .A2(_01318_),
    .A1(_01217_));
 sg13g2_xnor2_1 _09067_ (.Y(_01331_),
    .A(_01214_),
    .B(_01330_));
 sg13g2_nor2_1 _09068_ (.A(_01312_),
    .B(_01331_),
    .Y(_01332_));
 sg13g2_a22oi_1 _09069_ (.Y(_01333_),
    .B1(_01177_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .A2(_01175_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ));
 sg13g2_a22oi_1 _09070_ (.Y(_01334_),
    .B1(_01264_),
    .B2(net2245),
    .A2(_01167_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ));
 sg13g2_a22oi_1 _09071_ (.Y(_01335_),
    .B1(_01173_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .A2(_01161_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_a22oi_1 _09072_ (.Y(_01336_),
    .B1(_01178_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .A2(_01158_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ));
 sg13g2_a22oi_1 _09073_ (.Y(_01337_),
    .B1(_01179_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .A2(_01176_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ));
 sg13g2_nand3_1 _09074_ (.B(_01336_),
    .C(_01337_),
    .A(_01335_),
    .Y(_01338_));
 sg13g2_a221oi_1 _09075_ (.B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .C1(_01338_),
    .B1(_01171_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .Y(_01339_),
    .A2(_01168_));
 sg13g2_a22oi_1 _09076_ (.Y(_01340_),
    .B1(_01174_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A2(_01170_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ));
 sg13g2_nand4_1 _09077_ (.B(_01334_),
    .C(_01339_),
    .A(_01333_),
    .Y(_01341_),
    .D(_01340_));
 sg13g2_a22oi_1 _09078_ (.Y(_01342_),
    .B1(_01265_),
    .B2(\i_tinyqv.cpu.instr_data_start[8] ),
    .A2(net2244),
    .A1(net2409));
 sg13g2_nor2_2 _09079_ (.A(net2375),
    .B(net2317),
    .Y(_01343_));
 sg13g2_nand2_2 _09080_ (.Y(_01344_),
    .A(net2336),
    .B(net2318));
 sg13g2_nand2_1 _09081_ (.Y(_01345_),
    .A(net2417),
    .B(_01343_));
 sg13g2_nor2_2 _09082_ (.A(net2378),
    .B(net2307),
    .Y(_01346_));
 sg13g2_a22oi_1 _09083_ (.Y(_01347_),
    .B1(_01346_),
    .B2(\i_tinyqv.cpu.instr_data_start[12] ),
    .A2(net2243),
    .A1(\i_tinyqv.cpu.instr_data_start[16] ));
 sg13g2_nand3_1 _09084_ (.B(_01345_),
    .C(_01347_),
    .A(_01342_),
    .Y(_01348_));
 sg13g2_mux2_1 _09085_ (.A0(_01348_),
    .A1(_01341_),
    .S(_01192_),
    .X(_01349_));
 sg13g2_nand2_1 _09086_ (.Y(_01350_),
    .A(net2323),
    .B(_01349_));
 sg13g2_inv_1 _09087_ (.Y(_01351_),
    .A(_01350_));
 sg13g2_a22oi_1 _09088_ (.Y(_01352_),
    .B1(_01245_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .A2(_01244_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ));
 sg13g2_a22oi_1 _09089_ (.Y(_01353_),
    .B1(_01240_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .A2(_01234_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ));
 sg13g2_a22oi_1 _09090_ (.Y(_01354_),
    .B1(_01243_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .A2(_01239_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ));
 sg13g2_a22oi_1 _09091_ (.Y(_01355_),
    .B1(_01235_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .A2(_01230_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ));
 sg13g2_a22oi_1 _09092_ (.Y(_01356_),
    .B1(_01242_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .A2(_01237_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ));
 sg13g2_a22oi_1 _09093_ (.Y(_01357_),
    .B1(_01236_),
    .B2(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .A2(_01227_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ));
 sg13g2_nand3_1 _09094_ (.B(_01356_),
    .C(_01357_),
    .A(_01355_),
    .Y(_01358_));
 sg13g2_a221oi_1 _09095_ (.B2(net2245),
    .C1(_01358_),
    .B1(_01283_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .Y(_01359_),
    .A2(_01241_));
 sg13g2_nand4_1 _09096_ (.B(_01353_),
    .C(_01354_),
    .A(_01352_),
    .Y(_01360_),
    .D(_01359_));
 sg13g2_a21oi_1 _09097_ (.A1(\i_tinyqv.cpu.imm[16] ),
    .A2(net2313),
    .Y(_01361_),
    .B1(net2336));
 sg13g2_nor2_1 _09098_ (.A(_01075_),
    .B(net2324),
    .Y(_01362_));
 sg13g2_a221oi_1 _09099_ (.B2(\i_tinyqv.cpu.imm[28] ),
    .C1(_01362_),
    .B1(net2310),
    .A1(\i_tinyqv.cpu.imm[20] ),
    .Y(_01363_),
    .A2(net2320));
 sg13g2_nand2_1 _09100_ (.Y(_01364_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .B(net2313));
 sg13g2_a21o_1 _09101_ (.A2(net2325),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .B1(net2376),
    .X(_01365_));
 sg13g2_a221oi_1 _09102_ (.B2(\i_tinyqv.cpu.imm[12] ),
    .C1(_01365_),
    .B1(net2308),
    .A1(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .Y(_01366_),
    .A2(net2318));
 sg13g2_a22oi_1 _09103_ (.Y(_01367_),
    .B1(_01364_),
    .B2(_01366_),
    .A2(_01363_),
    .A1(_01361_));
 sg13g2_mux2_1 _09104_ (.A0(_01360_),
    .A1(_01367_),
    .S(_01217_),
    .X(_01368_));
 sg13g2_xnor2_1 _09105_ (.Y(_01369_),
    .A(_01214_),
    .B(_01368_));
 sg13g2_xor2_1 _09106_ (.B(_01369_),
    .A(_01350_),
    .X(_01370_));
 sg13g2_nor2_1 _09107_ (.A(net2375),
    .B(_01199_),
    .Y(_01371_));
 sg13g2_nand2_1 _09108_ (.Y(_01372_),
    .A(net2337),
    .B(net2314));
 sg13g2_nand2_1 _09109_ (.Y(_01373_),
    .A(\i_tinyqv.cpu.i_core.cy ),
    .B(net2233));
 sg13g2_o21ai_1 _09110_ (.B1(_01373_),
    .Y(_01374_),
    .A1(_01214_),
    .A2(net2233));
 sg13g2_nor2b_1 _09111_ (.A(_01370_),
    .B_N(_01374_),
    .Y(_01375_));
 sg13g2_a21oi_1 _09112_ (.A1(_01351_),
    .A2(_01369_),
    .Y(_01376_),
    .B1(_01375_));
 sg13g2_xnor2_1 _09113_ (.Y(_01377_),
    .A(_01312_),
    .B(_01331_));
 sg13g2_nor2_1 _09114_ (.A(_01376_),
    .B(_01377_),
    .Y(_01378_));
 sg13g2_nor2_1 _09115_ (.A(_01332_),
    .B(_01378_),
    .Y(_01379_));
 sg13g2_xnor2_1 _09116_ (.Y(_01380_),
    .A(_01276_),
    .B(_01294_));
 sg13g2_nor2b_1 _09117_ (.A(_01379_),
    .B_N(_01380_),
    .Y(_01381_));
 sg13g2_a21oi_1 _09118_ (.A1(_01276_),
    .A2(_01295_),
    .Y(_01382_),
    .B1(_01381_));
 sg13g2_xnor2_1 _09119_ (.Y(_01383_),
    .A(_01212_),
    .B(_01257_));
 sg13g2_or2_1 _09120_ (.X(_01384_),
    .B(_01383_),
    .A(_01382_));
 sg13g2_o21ai_1 _09121_ (.B1(_01384_),
    .Y(\i_tinyqv.cpu.i_core.cy_out ),
    .A1(_01212_),
    .A2(_01257_));
 sg13g2_nor2_2 _09122_ (.A(net2337),
    .B(net2307),
    .Y(_01385_));
 sg13g2_nand2_1 _09123_ (.Y(_01386_),
    .A(net2377),
    .B(net2308));
 sg13g2_a21oi_1 _09124_ (.A1(_01212_),
    .A2(_01257_),
    .Y(_01387_),
    .B1(_01213_));
 sg13g2_o21ai_1 _09125_ (.B1(_01213_),
    .Y(_01388_),
    .A1(\i_tinyqv.cpu.i_core.cmp ),
    .A2(net2236));
 sg13g2_nor2_1 _09126_ (.A(_01276_),
    .B(_01293_),
    .Y(_01389_));
 sg13g2_nand2_1 _09127_ (.Y(_01390_),
    .A(_01276_),
    .B(_01293_));
 sg13g2_nor2b_1 _09128_ (.A(_01389_),
    .B_N(_01390_),
    .Y(_01391_));
 sg13g2_xnor2_1 _09129_ (.Y(_01392_),
    .A(_01212_),
    .B(_01255_));
 sg13g2_nor2_1 _09130_ (.A(_01351_),
    .B(_01368_),
    .Y(_01393_));
 sg13g2_nand2_1 _09131_ (.Y(_01394_),
    .A(_01351_),
    .B(_01368_));
 sg13g2_nand2b_1 _09132_ (.Y(_01395_),
    .B(_01394_),
    .A_N(_01393_));
 sg13g2_or2_1 _09133_ (.X(_01396_),
    .B(_01330_),
    .A(_01312_));
 sg13g2_xnor2_1 _09134_ (.Y(_01397_),
    .A(_01312_),
    .B(_01330_));
 sg13g2_nand2_1 _09135_ (.Y(_01398_),
    .A(_01395_),
    .B(_01397_));
 sg13g2_nor4_1 _09136_ (.A(_01388_),
    .B(_01391_),
    .C(_01392_),
    .D(_01398_),
    .Y(_01399_));
 sg13g2_a21o_1 _09137_ (.A2(_01387_),
    .A1(_01384_),
    .B1(_01399_),
    .X(_01400_));
 sg13g2_xor2_1 _09138_ (.B(_01400_),
    .A(net2373),
    .X(_01401_));
 sg13g2_nor3_1 _09139_ (.A(net2503),
    .B(_01195_),
    .C(_01401_),
    .Y(_01402_));
 sg13g2_and2_1 _09140_ (.A(net2356),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .X(_01403_));
 sg13g2_and2_1 _09141_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.no_write_in_progress ),
    .X(_01404_));
 sg13g2_nand2_2 _09142_ (.Y(_01405_),
    .A(net3442),
    .B(\i_tinyqv.cpu.no_write_in_progress ));
 sg13g2_nand2_2 _09143_ (.Y(_01406_),
    .A(net2357),
    .B(net2303));
 sg13g2_and2_1 _09144_ (.A(net2355),
    .B(net3825),
    .X(_01407_));
 sg13g2_o21ai_1 _09145_ (.B1(net2355),
    .Y(_01408_),
    .A1(\i_tinyqv.cpu.is_alu_reg ),
    .A2(\i_tinyqv.cpu.is_alu_imm ));
 sg13g2_nand2_1 _09146_ (.Y(_01409_),
    .A(net2354),
    .B(net2371));
 sg13g2_nand2b_2 _09147_ (.Y(_01410_),
    .B(net2374),
    .A_N(net2371));
 sg13g2_nand2_1 _09148_ (.Y(_01411_),
    .A(_01409_),
    .B(_01410_));
 sg13g2_xor2_1 _09149_ (.B(_01411_),
    .A(net2504),
    .X(_01412_));
 sg13g2_nand4_1 _09150_ (.B(\i_tinyqv.cpu.i_core.load_done ),
    .C(_01403_),
    .A(\i_tinyqv.cpu.is_load ),
    .Y(_01413_),
    .D(_01408_));
 sg13g2_o21ai_1 _09151_ (.B1(_01413_),
    .Y(_01414_),
    .A1(_01408_),
    .A2(_01412_));
 sg13g2_o21ai_1 _09152_ (.B1(_01406_),
    .Y(_01415_),
    .A1(_01194_),
    .A2(_01414_));
 sg13g2_nor2_2 _09153_ (.A(\i_tinyqv.cpu.is_store ),
    .B(\i_tinyqv.cpu.is_load ),
    .Y(_01416_));
 sg13g2_o21ai_1 _09154_ (.B1(net2356),
    .Y(_01417_),
    .A1(\i_tinyqv.cpu.no_write_in_progress ),
    .A2(_01416_));
 sg13g2_and2_1 _09155_ (.A(net2355),
    .B(\i_tinyqv.cpu.is_system ),
    .X(_01418_));
 sg13g2_nand2_2 _09156_ (.Y(_01419_),
    .A(net2355),
    .B(\i_tinyqv.cpu.is_system ));
 sg13g2_nor4_1 _09157_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(\i_tinyqv.cpu.is_branch ),
    .C(_01417_),
    .D(_01418_),
    .Y(_01420_));
 sg13g2_nor2b_1 _09158_ (.A(net2504),
    .B_N(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .Y(_01421_));
 sg13g2_a21oi_1 _09159_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A2(_01421_),
    .Y(_01422_),
    .B1(_01406_));
 sg13g2_a21oi_2 _09160_ (.B1(_00923_),
    .Y(_01423_),
    .A2(_00926_),
    .A1(_00925_));
 sg13g2_o21ai_1 _09161_ (.B1(net2356),
    .Y(_01424_),
    .A1(\i_tinyqv.cpu.is_jal ),
    .A2(\i_tinyqv.cpu.is_jalr ));
 sg13g2_and2_1 _09162_ (.A(net2355),
    .B(\i_tinyqv.cpu.is_lui ),
    .X(_01425_));
 sg13g2_nand2_2 _09163_ (.Y(_01426_),
    .A(net2356),
    .B(\i_tinyqv.cpu.is_lui ));
 sg13g2_and3_1 _09164_ (.X(_01427_),
    .A(_01191_),
    .B(_01424_),
    .C(_01426_));
 sg13g2_nand2_1 _09165_ (.Y(_01428_),
    .A(_01420_),
    .B(_01427_));
 sg13g2_nor2_1 _09166_ (.A(_01422_),
    .B(_01428_),
    .Y(_01429_));
 sg13g2_o21ai_1 _09167_ (.B1(_01429_),
    .Y(_01430_),
    .A1(_01402_),
    .A2(_01415_));
 sg13g2_and2_1 _09168_ (.A(net2231),
    .B(_01430_),
    .X(_01431_));
 sg13g2_inv_2 _09169_ (.Y(_01432_),
    .A(_01431_));
 sg13g2_nor2_2 _09170_ (.A(_01417_),
    .B(_01432_),
    .Y(_01433_));
 sg13g2_a21o_2 _09171_ (.A2(_01431_),
    .A1(net3476),
    .B1(_01433_),
    .X(_00020_));
 sg13g2_nand2b_1 _09172_ (.Y(_01434_),
    .B(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .A_N(\i_tinyqv.mem.data_txn_len[0] ));
 sg13g2_xor2_1 _09173_ (.B(\i_tinyqv.mem.data_txn_len[1] ),
    .A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .X(_01435_));
 sg13g2_a21oi_1 _09174_ (.A1(_00985_),
    .A2(\i_tinyqv.mem.data_txn_len[0] ),
    .Y(_01436_),
    .B1(_01435_));
 sg13g2_and2_1 _09175_ (.A(_01434_),
    .B(_01436_),
    .X(_01437_));
 sg13g2_and2_1 _09176_ (.A(net3423),
    .B(_01437_),
    .X(_00073_));
 sg13g2_and2_1 _09177_ (.A(net2503),
    .B(_01305_),
    .X(_01438_));
 sg13g2_nand2_1 _09178_ (.Y(_01439_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .B(net2004));
 sg13g2_and2_1 _09179_ (.A(net2503),
    .B(_01341_),
    .X(_01440_));
 sg13g2_nand3_1 _09180_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .C(net1962),
    .A(net2465),
    .Y(_01441_));
 sg13g2_a21o_1 _09181_ (.A2(net1962),
    .A1(net2465),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .X(_01442_));
 sg13g2_nand2_1 _09182_ (.Y(_01443_),
    .A(_01441_),
    .B(_01442_));
 sg13g2_xor2_1 _09183_ (.B(_01443_),
    .A(_01439_),
    .X(_01444_));
 sg13g2_nand3_1 _09184_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .C(net1962),
    .A(net2466),
    .Y(_01445_));
 sg13g2_and4_1 _09185_ (.A(net2466),
    .B(net4161),
    .C(net1964),
    .D(_01444_),
    .X(_01446_));
 sg13g2_nor2b_2 _09186_ (.A(_01269_),
    .B_N(net2503),
    .Y(_01447_));
 sg13g2_nand2_1 _09187_ (.Y(_01448_),
    .A(net2466),
    .B(net2002));
 sg13g2_o21ai_1 _09188_ (.B1(_01441_),
    .Y(_01449_),
    .A1(_01439_),
    .A2(_01443_));
 sg13g2_nand2_1 _09189_ (.Y(_01450_),
    .A(net2465),
    .B(net2004));
 sg13g2_nand3_1 _09190_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .C(net1964),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .Y(_01451_));
 sg13g2_a21o_1 _09191_ (.A2(net1962),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .X(_01452_));
 sg13g2_nand2_1 _09192_ (.Y(_01453_),
    .A(_01451_),
    .B(_01452_));
 sg13g2_xor2_1 _09193_ (.B(_01453_),
    .A(_01450_),
    .X(_01454_));
 sg13g2_nand2_1 _09194_ (.Y(_01455_),
    .A(_01449_),
    .B(_01454_));
 sg13g2_xnor2_1 _09195_ (.Y(_01456_),
    .A(_01449_),
    .B(_01454_));
 sg13g2_xor2_1 _09196_ (.B(_01456_),
    .A(_01448_),
    .X(_01457_));
 sg13g2_nand2_1 _09197_ (.Y(_01458_),
    .A(_01446_),
    .B(_01457_));
 sg13g2_and2_1 _09198_ (.A(net2503),
    .B(_01189_),
    .X(_01459_));
 sg13g2_nand2_1 _09199_ (.Y(_01460_),
    .A(net2466),
    .B(net2000));
 sg13g2_o21ai_1 _09200_ (.B1(_01455_),
    .Y(_01461_),
    .A1(_01448_),
    .A2(_01456_));
 sg13g2_nand2_1 _09201_ (.Y(_01462_),
    .A(net2465),
    .B(net2002));
 sg13g2_o21ai_1 _09202_ (.B1(_01451_),
    .Y(_01463_),
    .A1(_01450_),
    .A2(_01453_));
 sg13g2_nand2_1 _09203_ (.Y(_01464_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net2004));
 sg13g2_nand3_1 _09204_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .C(net1962),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .Y(_01465_));
 sg13g2_a21o_1 _09205_ (.A2(net1962),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .X(_01466_));
 sg13g2_nand2_1 _09206_ (.Y(_01467_),
    .A(_01465_),
    .B(_01466_));
 sg13g2_xor2_1 _09207_ (.B(_01467_),
    .A(_01464_),
    .X(_01468_));
 sg13g2_nand2_1 _09208_ (.Y(_01469_),
    .A(_01463_),
    .B(_01468_));
 sg13g2_xnor2_1 _09209_ (.Y(_01470_),
    .A(_01463_),
    .B(_01468_));
 sg13g2_xor2_1 _09210_ (.B(_01470_),
    .A(_01462_),
    .X(_01471_));
 sg13g2_nand2_1 _09211_ (.Y(_01472_),
    .A(_01461_),
    .B(_01471_));
 sg13g2_xnor2_1 _09212_ (.Y(_01473_),
    .A(_01461_),
    .B(_01471_));
 sg13g2_xnor2_1 _09213_ (.Y(_01474_),
    .A(_01460_),
    .B(_01473_));
 sg13g2_nor2_1 _09214_ (.A(_01458_),
    .B(_01474_),
    .Y(_01475_));
 sg13g2_nand2_1 _09215_ (.Y(_01476_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .B(net2000));
 sg13g2_o21ai_1 _09216_ (.B1(_01469_),
    .Y(_01477_),
    .A1(_01462_),
    .A2(_01470_));
 sg13g2_nand2_1 _09217_ (.Y(_01478_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net2002));
 sg13g2_o21ai_1 _09218_ (.B1(_01465_),
    .Y(_01479_),
    .A1(_01464_),
    .A2(_01467_));
 sg13g2_nand2_1 _09219_ (.Y(_01480_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net2004));
 sg13g2_nand3_1 _09220_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .C(net1962),
    .A(net2464),
    .Y(_01481_));
 sg13g2_a21o_1 _09221_ (.A2(net1962),
    .A1(net2464),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .X(_01482_));
 sg13g2_nand2_1 _09222_ (.Y(_01483_),
    .A(_01481_),
    .B(_01482_));
 sg13g2_xor2_1 _09223_ (.B(_01483_),
    .A(_01480_),
    .X(_01484_));
 sg13g2_nand2_1 _09224_ (.Y(_01485_),
    .A(_01479_),
    .B(_01484_));
 sg13g2_xnor2_1 _09225_ (.Y(_01486_),
    .A(_01479_),
    .B(_01484_));
 sg13g2_xor2_1 _09226_ (.B(_01486_),
    .A(_01478_),
    .X(_01487_));
 sg13g2_nand2_1 _09227_ (.Y(_01488_),
    .A(_01477_),
    .B(_01487_));
 sg13g2_xnor2_1 _09228_ (.Y(_01489_),
    .A(_01477_),
    .B(_01487_));
 sg13g2_xor2_1 _09229_ (.B(_01489_),
    .A(_01476_),
    .X(_01490_));
 sg13g2_o21ai_1 _09230_ (.B1(_01472_),
    .Y(_01491_),
    .A1(_01460_),
    .A2(_01473_));
 sg13g2_nand2_1 _09231_ (.Y(_01492_),
    .A(_01490_),
    .B(_01491_));
 sg13g2_xor2_1 _09232_ (.B(_01491_),
    .A(_01490_),
    .X(_01493_));
 sg13g2_nand2_1 _09233_ (.Y(_01494_),
    .A(_01475_),
    .B(_01493_));
 sg13g2_xor2_1 _09234_ (.B(_01493_),
    .A(_01475_),
    .X(_00007_));
 sg13g2_nand2_1 _09235_ (.Y(_01495_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .B(net2000));
 sg13g2_o21ai_1 _09236_ (.B1(_01485_),
    .Y(_01496_),
    .A1(_01478_),
    .A2(_01486_));
 sg13g2_nand2_1 _09237_ (.Y(_01497_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(_01447_));
 sg13g2_o21ai_1 _09238_ (.B1(_01481_),
    .Y(_01498_),
    .A1(_01480_),
    .A2(_01483_));
 sg13g2_nand2_1 _09239_ (.Y(_01499_),
    .A(net2464),
    .B(net2004));
 sg13g2_nand3_1 _09240_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .C(net1963),
    .A(net2463),
    .Y(_01500_));
 sg13g2_a21o_1 _09241_ (.A2(net1963),
    .A1(net2463),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .X(_01501_));
 sg13g2_nand2_1 _09242_ (.Y(_01502_),
    .A(_01500_),
    .B(_01501_));
 sg13g2_xor2_1 _09243_ (.B(_01502_),
    .A(_01499_),
    .X(_01503_));
 sg13g2_nand2_1 _09244_ (.Y(_01504_),
    .A(_01498_),
    .B(_01503_));
 sg13g2_xnor2_1 _09245_ (.Y(_01505_),
    .A(_01498_),
    .B(_01503_));
 sg13g2_xor2_1 _09246_ (.B(_01505_),
    .A(_01497_),
    .X(_01506_));
 sg13g2_nand2_1 _09247_ (.Y(_01507_),
    .A(_01496_),
    .B(_01506_));
 sg13g2_xnor2_1 _09248_ (.Y(_01508_),
    .A(_01496_),
    .B(_01506_));
 sg13g2_xor2_1 _09249_ (.B(_01508_),
    .A(_01495_),
    .X(_01509_));
 sg13g2_o21ai_1 _09250_ (.B1(_01488_),
    .Y(_01510_),
    .A1(_01476_),
    .A2(_01489_));
 sg13g2_nand2_1 _09251_ (.Y(_01511_),
    .A(_01509_),
    .B(_01510_));
 sg13g2_xnor2_1 _09252_ (.Y(_01512_),
    .A(_01509_),
    .B(_01510_));
 sg13g2_a21o_1 _09253_ (.A2(_01494_),
    .A1(_01492_),
    .B1(_01512_),
    .X(_01513_));
 sg13g2_nand3_1 _09254_ (.B(_01494_),
    .C(_01512_),
    .A(_01492_),
    .Y(_01514_));
 sg13g2_and2_1 _09255_ (.A(_01513_),
    .B(_01514_),
    .X(_00010_));
 sg13g2_nand2_1 _09256_ (.Y(_01515_),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .B(net2000));
 sg13g2_o21ai_1 _09257_ (.B1(_01504_),
    .Y(_01516_),
    .A1(_01497_),
    .A2(_01505_));
 sg13g2_nand2_1 _09258_ (.Y(_01517_),
    .A(net2464),
    .B(net2002));
 sg13g2_o21ai_1 _09259_ (.B1(_01500_),
    .Y(_01518_),
    .A1(_01499_),
    .A2(_01502_));
 sg13g2_nand2_1 _09260_ (.Y(_01519_),
    .A(net2463),
    .B(net2004));
 sg13g2_nand3_1 _09261_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .C(net1963),
    .A(net2461),
    .Y(_01520_));
 sg13g2_a21o_1 _09262_ (.A2(net1963),
    .A1(net2461),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .X(_01521_));
 sg13g2_nand2_1 _09263_ (.Y(_01522_),
    .A(_01520_),
    .B(_01521_));
 sg13g2_xor2_1 _09264_ (.B(_01522_),
    .A(_01519_),
    .X(_01523_));
 sg13g2_nand2_1 _09265_ (.Y(_01524_),
    .A(_01518_),
    .B(_01523_));
 sg13g2_xnor2_1 _09266_ (.Y(_01525_),
    .A(_01518_),
    .B(_01523_));
 sg13g2_xor2_1 _09267_ (.B(_01525_),
    .A(_01517_),
    .X(_01526_));
 sg13g2_nand2_1 _09268_ (.Y(_01527_),
    .A(_01516_),
    .B(_01526_));
 sg13g2_xnor2_1 _09269_ (.Y(_01528_),
    .A(_01516_),
    .B(_01526_));
 sg13g2_xor2_1 _09270_ (.B(_01528_),
    .A(_01515_),
    .X(_01529_));
 sg13g2_o21ai_1 _09271_ (.B1(_01507_),
    .Y(_01530_),
    .A1(_01495_),
    .A2(_01508_));
 sg13g2_nand2_1 _09272_ (.Y(_01531_),
    .A(_01529_),
    .B(_01530_));
 sg13g2_xnor2_1 _09273_ (.Y(_01532_),
    .A(_01529_),
    .B(_01530_));
 sg13g2_a21o_1 _09274_ (.A2(_01513_),
    .A1(_01511_),
    .B1(_01532_),
    .X(_01533_));
 sg13g2_nand3_1 _09275_ (.B(_01513_),
    .C(_01532_),
    .A(_01511_),
    .Y(_01534_));
 sg13g2_and2_1 _09276_ (.A(_01533_),
    .B(_01534_),
    .X(_00011_));
 sg13g2_nand2_1 _09277_ (.Y(_01535_),
    .A(net2464),
    .B(net2000));
 sg13g2_o21ai_1 _09278_ (.B1(_01524_),
    .Y(_01536_),
    .A1(_01517_),
    .A2(_01525_));
 sg13g2_nand2_1 _09279_ (.Y(_01537_),
    .A(net2463),
    .B(net2002));
 sg13g2_o21ai_1 _09280_ (.B1(_01520_),
    .Y(_01538_),
    .A1(_01519_),
    .A2(_01522_));
 sg13g2_nand2_1 _09281_ (.Y(_01539_),
    .A(net2461),
    .B(_01438_));
 sg13g2_nand3_1 _09282_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .C(net1963),
    .A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .Y(_01540_));
 sg13g2_a21o_1 _09283_ (.A2(net1963),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .X(_01541_));
 sg13g2_nand2_1 _09284_ (.Y(_01542_),
    .A(_01540_),
    .B(_01541_));
 sg13g2_xor2_1 _09285_ (.B(_01542_),
    .A(_01539_),
    .X(_01543_));
 sg13g2_nand2_1 _09286_ (.Y(_01544_),
    .A(_01538_),
    .B(_01543_));
 sg13g2_xnor2_1 _09287_ (.Y(_01545_),
    .A(_01538_),
    .B(_01543_));
 sg13g2_xor2_1 _09288_ (.B(_01545_),
    .A(_01537_),
    .X(_01546_));
 sg13g2_nand2_1 _09289_ (.Y(_01547_),
    .A(_01536_),
    .B(_01546_));
 sg13g2_xnor2_1 _09290_ (.Y(_01548_),
    .A(_01536_),
    .B(_01546_));
 sg13g2_xor2_1 _09291_ (.B(_01548_),
    .A(_01535_),
    .X(_01549_));
 sg13g2_o21ai_1 _09292_ (.B1(_01527_),
    .Y(_01550_),
    .A1(_01515_),
    .A2(_01528_));
 sg13g2_xnor2_1 _09293_ (.Y(_01551_),
    .A(_01549_),
    .B(_01550_));
 sg13g2_a21oi_1 _09294_ (.A1(_01531_),
    .A2(_01533_),
    .Y(_01552_),
    .B1(_01551_));
 sg13g2_nand3_1 _09295_ (.B(_01533_),
    .C(_01551_),
    .A(_01531_),
    .Y(_01553_));
 sg13g2_nor2b_1 _09296_ (.A(_01552_),
    .B_N(_01553_),
    .Y(_00012_));
 sg13g2_a21o_1 _09297_ (.A2(_01550_),
    .A1(_01549_),
    .B1(_01552_),
    .X(_01554_));
 sg13g2_o21ai_1 _09298_ (.B1(_01547_),
    .Y(_01555_),
    .A1(_01535_),
    .A2(_01548_));
 sg13g2_nand2_1 _09299_ (.Y(_01556_),
    .A(net2463),
    .B(net2000));
 sg13g2_o21ai_1 _09300_ (.B1(_01544_),
    .Y(_01557_),
    .A1(_01537_),
    .A2(_01545_));
 sg13g2_nand2_1 _09301_ (.Y(_01558_),
    .A(net2461),
    .B(net2002));
 sg13g2_o21ai_1 _09302_ (.B1(_01540_),
    .Y(_01559_),
    .A1(_01539_),
    .A2(_01542_));
 sg13g2_nand2_1 _09303_ (.Y(_01560_),
    .A(net2460),
    .B(net2003));
 sg13g2_nand3_1 _09304_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .C(net1961),
    .A(net2459),
    .Y(_01561_));
 sg13g2_a21o_1 _09305_ (.A2(net1961),
    .A1(net2459),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .X(_01562_));
 sg13g2_nand2_1 _09306_ (.Y(_01563_),
    .A(_01561_),
    .B(_01562_));
 sg13g2_xor2_1 _09307_ (.B(_01563_),
    .A(_01560_),
    .X(_01564_));
 sg13g2_nand2_1 _09308_ (.Y(_01565_),
    .A(_01559_),
    .B(_01564_));
 sg13g2_xnor2_1 _09309_ (.Y(_01566_),
    .A(_01559_),
    .B(_01564_));
 sg13g2_xor2_1 _09310_ (.B(_01566_),
    .A(_01558_),
    .X(_01567_));
 sg13g2_nand2_1 _09311_ (.Y(_01568_),
    .A(_01557_),
    .B(_01567_));
 sg13g2_xnor2_1 _09312_ (.Y(_01569_),
    .A(_01557_),
    .B(_01567_));
 sg13g2_xor2_1 _09313_ (.B(_01569_),
    .A(_01556_),
    .X(_01570_));
 sg13g2_nand2_1 _09314_ (.Y(_01571_),
    .A(_01555_),
    .B(_01570_));
 sg13g2_xnor2_1 _09315_ (.Y(_01572_),
    .A(_01555_),
    .B(_01570_));
 sg13g2_nand2b_1 _09316_ (.Y(_01573_),
    .B(_01554_),
    .A_N(_01572_));
 sg13g2_xnor2_1 _09317_ (.Y(_00013_),
    .A(_01554_),
    .B(_01572_));
 sg13g2_nand2_1 _09318_ (.Y(_01574_),
    .A(net2461),
    .B(_01459_));
 sg13g2_o21ai_1 _09319_ (.B1(_01565_),
    .Y(_01575_),
    .A1(_01558_),
    .A2(_01566_));
 sg13g2_nand2_1 _09320_ (.Y(_01576_),
    .A(net2460),
    .B(net2001));
 sg13g2_o21ai_1 _09321_ (.B1(_01561_),
    .Y(_01577_),
    .A1(_01560_),
    .A2(_01563_));
 sg13g2_nand2_1 _09322_ (.Y(_01578_),
    .A(net2459),
    .B(net2004));
 sg13g2_nand3_1 _09323_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .C(net1961),
    .A(net2458),
    .Y(_01579_));
 sg13g2_a21o_1 _09324_ (.A2(net1961),
    .A1(net2458),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .X(_01580_));
 sg13g2_nand2_1 _09325_ (.Y(_01581_),
    .A(_01579_),
    .B(_01580_));
 sg13g2_xor2_1 _09326_ (.B(_01581_),
    .A(_01578_),
    .X(_01582_));
 sg13g2_nand2_1 _09327_ (.Y(_01583_),
    .A(_01577_),
    .B(_01582_));
 sg13g2_xnor2_1 _09328_ (.Y(_01584_),
    .A(_01577_),
    .B(_01582_));
 sg13g2_xor2_1 _09329_ (.B(_01584_),
    .A(_01576_),
    .X(_01585_));
 sg13g2_nand2_1 _09330_ (.Y(_01586_),
    .A(_01575_),
    .B(_01585_));
 sg13g2_xnor2_1 _09331_ (.Y(_01587_),
    .A(_01575_),
    .B(_01585_));
 sg13g2_xor2_1 _09332_ (.B(_01587_),
    .A(_01574_),
    .X(_01588_));
 sg13g2_o21ai_1 _09333_ (.B1(_01568_),
    .Y(_01589_),
    .A1(_01556_),
    .A2(_01569_));
 sg13g2_nand2_1 _09334_ (.Y(_01590_),
    .A(_01588_),
    .B(_01589_));
 sg13g2_xnor2_1 _09335_ (.Y(_01591_),
    .A(_01588_),
    .B(_01589_));
 sg13g2_a21o_1 _09336_ (.A2(_01573_),
    .A1(_01571_),
    .B1(_01591_),
    .X(_01592_));
 sg13g2_nand3_1 _09337_ (.B(_01573_),
    .C(_01591_),
    .A(_01571_),
    .Y(_01593_));
 sg13g2_and2_1 _09338_ (.A(_01592_),
    .B(_01593_),
    .X(_00014_));
 sg13g2_nand2_1 _09339_ (.Y(_01594_),
    .A(net2460),
    .B(net1999));
 sg13g2_o21ai_1 _09340_ (.B1(_01583_),
    .Y(_01595_),
    .A1(_01576_),
    .A2(_01584_));
 sg13g2_nand2_1 _09341_ (.Y(_01596_),
    .A(net2459),
    .B(net2002));
 sg13g2_o21ai_1 _09342_ (.B1(_01579_),
    .Y(_01597_),
    .A1(_01578_),
    .A2(_01581_));
 sg13g2_nand2_1 _09343_ (.Y(_01598_),
    .A(net2458),
    .B(net2003));
 sg13g2_nand3_1 _09344_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .C(net1959),
    .A(net2457),
    .Y(_01599_));
 sg13g2_a21o_1 _09345_ (.A2(net1959),
    .A1(net2457),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .X(_01600_));
 sg13g2_nand2_1 _09346_ (.Y(_01601_),
    .A(_01599_),
    .B(_01600_));
 sg13g2_xor2_1 _09347_ (.B(_01601_),
    .A(_01598_),
    .X(_01602_));
 sg13g2_nand2_1 _09348_ (.Y(_01603_),
    .A(_01597_),
    .B(_01602_));
 sg13g2_xnor2_1 _09349_ (.Y(_01604_),
    .A(_01597_),
    .B(_01602_));
 sg13g2_xor2_1 _09350_ (.B(_01604_),
    .A(_01596_),
    .X(_01605_));
 sg13g2_nand2_1 _09351_ (.Y(_01606_),
    .A(_01595_),
    .B(_01605_));
 sg13g2_xnor2_1 _09352_ (.Y(_01607_),
    .A(_01595_),
    .B(_01605_));
 sg13g2_xor2_1 _09353_ (.B(_01607_),
    .A(_01594_),
    .X(_01608_));
 sg13g2_o21ai_1 _09354_ (.B1(_01586_),
    .Y(_01609_),
    .A1(_01574_),
    .A2(_01587_));
 sg13g2_xnor2_1 _09355_ (.Y(_01610_),
    .A(_01608_),
    .B(_01609_));
 sg13g2_a21oi_1 _09356_ (.A1(_01590_),
    .A2(_01592_),
    .Y(_01611_),
    .B1(_01610_));
 sg13g2_nand3_1 _09357_ (.B(_01592_),
    .C(_01610_),
    .A(_01590_),
    .Y(_01612_));
 sg13g2_nor2b_1 _09358_ (.A(_01611_),
    .B_N(_01612_),
    .Y(_00015_));
 sg13g2_a21o_1 _09359_ (.A2(_01609_),
    .A1(_01608_),
    .B1(_01611_),
    .X(_01613_));
 sg13g2_o21ai_1 _09360_ (.B1(_01606_),
    .Y(_01614_),
    .A1(_01594_),
    .A2(_01607_));
 sg13g2_nand2_1 _09361_ (.Y(_01615_),
    .A(net2459),
    .B(net2000));
 sg13g2_o21ai_1 _09362_ (.B1(_01603_),
    .Y(_01616_),
    .A1(_01596_),
    .A2(_01604_));
 sg13g2_nand2_1 _09363_ (.Y(_01617_),
    .A(net2458),
    .B(net2001));
 sg13g2_o21ai_1 _09364_ (.B1(_01599_),
    .Y(_01618_),
    .A1(_01598_),
    .A2(_01601_));
 sg13g2_nand2_1 _09365_ (.Y(_01619_),
    .A(net2457),
    .B(net2003));
 sg13g2_nand3_1 _09366_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .C(net1959),
    .A(net2456),
    .Y(_01620_));
 sg13g2_a21o_1 _09367_ (.A2(net1959),
    .A1(net2456),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .X(_01621_));
 sg13g2_nand2_1 _09368_ (.Y(_01622_),
    .A(_01620_),
    .B(_01621_));
 sg13g2_xor2_1 _09369_ (.B(_01622_),
    .A(_01619_),
    .X(_01623_));
 sg13g2_nand2_1 _09370_ (.Y(_01624_),
    .A(_01618_),
    .B(_01623_));
 sg13g2_xnor2_1 _09371_ (.Y(_01625_),
    .A(_01618_),
    .B(_01623_));
 sg13g2_xor2_1 _09372_ (.B(_01625_),
    .A(_01617_),
    .X(_01626_));
 sg13g2_nand2_1 _09373_ (.Y(_01627_),
    .A(_01616_),
    .B(_01626_));
 sg13g2_xnor2_1 _09374_ (.Y(_01628_),
    .A(_01616_),
    .B(_01626_));
 sg13g2_xor2_1 _09375_ (.B(_01628_),
    .A(_01615_),
    .X(_01629_));
 sg13g2_xnor2_1 _09376_ (.Y(_01630_),
    .A(_01614_),
    .B(_01629_));
 sg13g2_nor2b_1 _09377_ (.A(_01630_),
    .B_N(_01613_),
    .Y(_01631_));
 sg13g2_xnor2_1 _09378_ (.Y(_00016_),
    .A(_01613_),
    .B(_01630_));
 sg13g2_a21o_1 _09379_ (.A2(_01629_),
    .A1(_01614_),
    .B1(_01631_),
    .X(_01632_));
 sg13g2_o21ai_1 _09380_ (.B1(_01627_),
    .Y(_01633_),
    .A1(_01615_),
    .A2(_01628_));
 sg13g2_nand2_1 _09381_ (.Y(_01634_),
    .A(net2458),
    .B(net1999));
 sg13g2_o21ai_1 _09382_ (.B1(_01624_),
    .Y(_01635_),
    .A1(_01617_),
    .A2(_01625_));
 sg13g2_nand2_1 _09383_ (.Y(_01636_),
    .A(net2457),
    .B(net2001));
 sg13g2_o21ai_1 _09384_ (.B1(_01620_),
    .Y(_01637_),
    .A1(_01619_),
    .A2(_01622_));
 sg13g2_nand2_1 _09385_ (.Y(_01638_),
    .A(net2456),
    .B(net2003));
 sg13g2_nand3_1 _09386_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .C(net1959),
    .A(net2455),
    .Y(_01639_));
 sg13g2_a21o_1 _09387_ (.A2(net1959),
    .A1(net2455),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .X(_01640_));
 sg13g2_nand2_1 _09388_ (.Y(_01641_),
    .A(_01639_),
    .B(_01640_));
 sg13g2_xor2_1 _09389_ (.B(_01641_),
    .A(_01638_),
    .X(_01642_));
 sg13g2_nand2_1 _09390_ (.Y(_01643_),
    .A(_01637_),
    .B(_01642_));
 sg13g2_xnor2_1 _09391_ (.Y(_01644_),
    .A(_01637_),
    .B(_01642_));
 sg13g2_xor2_1 _09392_ (.B(_01644_),
    .A(_01636_),
    .X(_01645_));
 sg13g2_nand2_1 _09393_ (.Y(_01646_),
    .A(_01635_),
    .B(_01645_));
 sg13g2_xnor2_1 _09394_ (.Y(_01647_),
    .A(_01635_),
    .B(_01645_));
 sg13g2_xor2_1 _09395_ (.B(_01647_),
    .A(_01634_),
    .X(_01648_));
 sg13g2_xnor2_1 _09396_ (.Y(_01649_),
    .A(_01633_),
    .B(_01648_));
 sg13g2_nor2b_1 _09397_ (.A(_01649_),
    .B_N(_01632_),
    .Y(_01650_));
 sg13g2_xnor2_1 _09398_ (.Y(_00017_),
    .A(_01632_),
    .B(_01649_));
 sg13g2_a21o_1 _09399_ (.A2(_01648_),
    .A1(_01633_),
    .B1(_01650_),
    .X(_01651_));
 sg13g2_o21ai_1 _09400_ (.B1(_01646_),
    .Y(_01652_),
    .A1(_01634_),
    .A2(_01647_));
 sg13g2_nand2_1 _09401_ (.Y(_01653_),
    .A(net2457),
    .B(net1999));
 sg13g2_o21ai_1 _09402_ (.B1(_01643_),
    .Y(_01654_),
    .A1(_01636_),
    .A2(_01644_));
 sg13g2_nand2_1 _09403_ (.Y(_01655_),
    .A(net2456),
    .B(net2001));
 sg13g2_o21ai_1 _09404_ (.B1(_01639_),
    .Y(_01656_),
    .A1(_01638_),
    .A2(_01641_));
 sg13g2_nand2_1 _09405_ (.Y(_01657_),
    .A(net2455),
    .B(net2003));
 sg13g2_nand3_1 _09406_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .C(net1959),
    .A(net2454),
    .Y(_01658_));
 sg13g2_a21o_1 _09407_ (.A2(net1960),
    .A1(net2454),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .X(_01659_));
 sg13g2_nand2_1 _09408_ (.Y(_01660_),
    .A(_01658_),
    .B(_01659_));
 sg13g2_xor2_1 _09409_ (.B(_01660_),
    .A(_01657_),
    .X(_01661_));
 sg13g2_nand2_1 _09410_ (.Y(_01662_),
    .A(_01656_),
    .B(_01661_));
 sg13g2_xnor2_1 _09411_ (.Y(_01663_),
    .A(_01656_),
    .B(_01661_));
 sg13g2_xor2_1 _09412_ (.B(_01663_),
    .A(_01655_),
    .X(_01664_));
 sg13g2_nand2_1 _09413_ (.Y(_01665_),
    .A(_01654_),
    .B(_01664_));
 sg13g2_xnor2_1 _09414_ (.Y(_01666_),
    .A(_01654_),
    .B(_01664_));
 sg13g2_xor2_1 _09415_ (.B(_01666_),
    .A(_01653_),
    .X(_01667_));
 sg13g2_xnor2_1 _09416_ (.Y(_01668_),
    .A(_01652_),
    .B(_01667_));
 sg13g2_nor2b_1 _09417_ (.A(_01668_),
    .B_N(_01651_),
    .Y(_01669_));
 sg13g2_xnor2_1 _09418_ (.Y(_00018_),
    .A(_01651_),
    .B(_01668_));
 sg13g2_a21o_1 _09419_ (.A2(_01667_),
    .A1(_01652_),
    .B1(_01669_),
    .X(_01670_));
 sg13g2_o21ai_1 _09420_ (.B1(_01665_),
    .Y(_01671_),
    .A1(_01653_),
    .A2(_01666_));
 sg13g2_nand2_1 _09421_ (.Y(_01672_),
    .A(net2456),
    .B(net1999));
 sg13g2_o21ai_1 _09422_ (.B1(_01662_),
    .Y(_01673_),
    .A1(_01655_),
    .A2(_01663_));
 sg13g2_nand2_1 _09423_ (.Y(_01674_),
    .A(net2455),
    .B(net2001));
 sg13g2_o21ai_1 _09424_ (.B1(_01658_),
    .Y(_01675_),
    .A1(_01657_),
    .A2(_01660_));
 sg13g2_nand2_1 _09425_ (.Y(_01676_),
    .A(net2454),
    .B(net2003));
 sg13g2_nand3_1 _09426_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .C(net1959),
    .A(net2453),
    .Y(_01677_));
 sg13g2_a21o_1 _09427_ (.A2(net1960),
    .A1(net2453),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .X(_01678_));
 sg13g2_nand2_1 _09428_ (.Y(_01679_),
    .A(_01677_),
    .B(_01678_));
 sg13g2_xor2_1 _09429_ (.B(_01679_),
    .A(_01676_),
    .X(_01680_));
 sg13g2_nand2_1 _09430_ (.Y(_01681_),
    .A(_01675_),
    .B(_01680_));
 sg13g2_xnor2_1 _09431_ (.Y(_01682_),
    .A(_01675_),
    .B(_01680_));
 sg13g2_xor2_1 _09432_ (.B(_01682_),
    .A(_01674_),
    .X(_01683_));
 sg13g2_nand2_1 _09433_ (.Y(_01684_),
    .A(_01673_),
    .B(_01683_));
 sg13g2_xnor2_1 _09434_ (.Y(_01685_),
    .A(_01673_),
    .B(_01683_));
 sg13g2_xor2_1 _09435_ (.B(_01685_),
    .A(_01672_),
    .X(_01686_));
 sg13g2_nand2_1 _09436_ (.Y(_01687_),
    .A(_01671_),
    .B(_01686_));
 sg13g2_xnor2_1 _09437_ (.Y(_01688_),
    .A(_01671_),
    .B(_01686_));
 sg13g2_nand2b_1 _09438_ (.Y(_01689_),
    .B(_01670_),
    .A_N(_01688_));
 sg13g2_xnor2_1 _09439_ (.Y(_00008_),
    .A(_01670_),
    .B(_01688_));
 sg13g2_nand2_1 _09440_ (.Y(_01690_),
    .A(net2455),
    .B(net1999));
 sg13g2_o21ai_1 _09441_ (.B1(_01681_),
    .Y(_01691_),
    .A1(_01674_),
    .A2(_01682_));
 sg13g2_nand2_1 _09442_ (.Y(_01692_),
    .A(net2454),
    .B(net2001));
 sg13g2_o21ai_1 _09443_ (.B1(_01677_),
    .Y(_01693_),
    .A1(_01676_),
    .A2(_01679_));
 sg13g2_nand2_2 _09444_ (.Y(_01694_),
    .A(net2453),
    .B(net2003));
 sg13g2_nand3_1 _09445_ (.B(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .C(net1960),
    .A(net2452),
    .Y(_01695_));
 sg13g2_a21o_1 _09446_ (.A2(net1960),
    .A1(net2452),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .X(_01696_));
 sg13g2_nand2_1 _09447_ (.Y(_01697_),
    .A(_01695_),
    .B(_01696_));
 sg13g2_xor2_1 _09448_ (.B(_01697_),
    .A(_01694_),
    .X(_01698_));
 sg13g2_nand2_1 _09449_ (.Y(_01699_),
    .A(_01693_),
    .B(_01698_));
 sg13g2_xnor2_1 _09450_ (.Y(_01700_),
    .A(_01693_),
    .B(_01698_));
 sg13g2_xor2_1 _09451_ (.B(_01700_),
    .A(_01692_),
    .X(_01701_));
 sg13g2_nand2_1 _09452_ (.Y(_01702_),
    .A(_01691_),
    .B(_01701_));
 sg13g2_xnor2_1 _09453_ (.Y(_01703_),
    .A(_01691_),
    .B(_01701_));
 sg13g2_or2_1 _09454_ (.X(_01704_),
    .B(_01703_),
    .A(_01690_));
 sg13g2_xor2_1 _09455_ (.B(_01703_),
    .A(_01690_),
    .X(_01705_));
 sg13g2_o21ai_1 _09456_ (.B1(_01684_),
    .Y(_01706_),
    .A1(_01672_),
    .A2(_01685_));
 sg13g2_nand2_1 _09457_ (.Y(_01707_),
    .A(_01705_),
    .B(_01706_));
 sg13g2_xnor2_1 _09458_ (.Y(_01708_),
    .A(_01705_),
    .B(_01706_));
 sg13g2_a21o_1 _09459_ (.A2(_01689_),
    .A1(_01687_),
    .B1(_01708_),
    .X(_01709_));
 sg13g2_nand3_1 _09460_ (.B(_01689_),
    .C(_01708_),
    .A(_01687_),
    .Y(_01710_));
 sg13g2_and2_1 _09461_ (.A(_01709_),
    .B(_01710_),
    .X(_00009_));
 sg13g2_nand2_1 _09462_ (.Y(_01711_),
    .A(net2373),
    .B(net2323));
 sg13g2_nand2_1 _09463_ (.Y(_01712_),
    .A(_01400_),
    .B(_01711_));
 sg13g2_o21ai_1 _09464_ (.B1(_01712_),
    .Y(\i_tinyqv.cpu.i_core.cmp_out ),
    .A1(\i_tinyqv.cpu.i_core.cy_out ),
    .A2(_01711_));
 sg13g2_nand2_2 _09465_ (.Y(_01713_),
    .A(_01191_),
    .B(_01408_));
 sg13g2_and2_1 _09466_ (.A(net2367),
    .B(net2466),
    .X(_01714_));
 sg13g2_nor2b_2 _09467_ (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .B_N(net2503),
    .Y(_01715_));
 sg13g2_nand2b_2 _09468_ (.Y(_01716_),
    .B(net2503),
    .A_N(net3576));
 sg13g2_nor2_1 _09469_ (.A(_01193_),
    .B(_01716_),
    .Y(_01717_));
 sg13g2_nand2b_2 _09470_ (.Y(_01718_),
    .B(_01715_),
    .A_N(_01193_));
 sg13g2_nand2_1 _09471_ (.Y(_01719_),
    .A(_01714_),
    .B(_01717_));
 sg13g2_nand2_2 _09472_ (.Y(_01720_),
    .A(\i_tinyqv.cpu.alu_op[3] ),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[31] ));
 sg13g2_xnor2_1 _09473_ (.Y(_01721_),
    .A(net2368),
    .B(net2375));
 sg13g2_nor2_1 _09474_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_01721_),
    .Y(_01722_));
 sg13g2_nand2_1 _09475_ (.Y(_01723_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .B(_01721_));
 sg13g2_xor2_1 _09476_ (.B(net2381),
    .A(net2368),
    .X(_01724_));
 sg13g2_nor2_1 _09477_ (.A(_01122_),
    .B(_01724_),
    .Y(_01725_));
 sg13g2_xnor2_1 _09478_ (.Y(_01726_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .B(_01724_));
 sg13g2_xnor2_1 _09479_ (.Y(_01727_),
    .A(net2370),
    .B(net2384));
 sg13g2_and2_1 _09480_ (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_01727_),
    .X(_01728_));
 sg13g2_nand2_1 _09481_ (.Y(_01729_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_01727_));
 sg13g2_a21oi_1 _09482_ (.A1(_01726_),
    .A2(_01728_),
    .Y(_01730_),
    .B1(_01725_));
 sg13g2_o21ai_1 _09483_ (.B1(_01723_),
    .Y(_01731_),
    .A1(_01722_),
    .A2(_01730_));
 sg13g2_and2_1 _09484_ (.A(_01720_),
    .B(_01731_),
    .X(_01732_));
 sg13g2_nand2_1 _09485_ (.Y(_01733_),
    .A(_01720_),
    .B(_01731_));
 sg13g2_mux2_1 _09486_ (.A0(net2452),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net2363),
    .X(_01734_));
 sg13g2_or2_1 _09487_ (.X(_01735_),
    .B(net2453),
    .A(net2363));
 sg13g2_o21ai_1 _09488_ (.B1(_01735_),
    .Y(_01736_),
    .A1(net2353),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[17] ));
 sg13g2_nor2_1 _09489_ (.A(net2473),
    .B(_01734_),
    .Y(_01737_));
 sg13g2_a21oi_1 _09490_ (.A1(net2472),
    .A2(_01736_),
    .Y(_01738_),
    .B1(_01737_));
 sg13g2_xor2_1 _09491_ (.B(_01727_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .X(_01739_));
 sg13g2_xnor2_1 _09492_ (.Y(_01740_),
    .A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .B(_01727_));
 sg13g2_mux2_1 _09493_ (.A0(net2454),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(net2364),
    .X(_01741_));
 sg13g2_mux2_1 _09494_ (.A0(net2455),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(net2364),
    .X(_01742_));
 sg13g2_mux2_1 _09495_ (.A0(_01741_),
    .A1(_01742_),
    .S(net2473),
    .X(_01743_));
 sg13g2_xnor2_1 _09496_ (.Y(_01744_),
    .A(_01726_),
    .B(_01729_));
 sg13g2_xnor2_1 _09497_ (.Y(_01745_),
    .A(_01726_),
    .B(_01728_));
 sg13g2_or2_1 _09498_ (.X(_01746_),
    .B(net2456),
    .A(net2363));
 sg13g2_o21ai_1 _09499_ (.B1(_01746_),
    .Y(_01747_),
    .A1(net2353),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[20] ));
 sg13g2_mux2_1 _09500_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(net2363),
    .X(_01748_));
 sg13g2_nand2_1 _09501_ (.Y(_01749_),
    .A(net2473),
    .B(_01748_));
 sg13g2_o21ai_1 _09502_ (.B1(_01749_),
    .Y(_01750_),
    .A1(net2472),
    .A2(_01747_));
 sg13g2_mux4_1 _09503_ (.S0(net2363),
    .A0(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S1(net2474),
    .X(_01751_));
 sg13g2_nand2b_1 _09504_ (.Y(_01752_),
    .B(_01723_),
    .A_N(_01722_));
 sg13g2_and2_1 _09505_ (.A(_01730_),
    .B(_01752_),
    .X(_01753_));
 sg13g2_nand2_2 _09506_ (.Y(_01754_),
    .A(_01730_),
    .B(_01752_));
 sg13g2_nand2_1 _09507_ (.Y(_01755_),
    .A(net2362),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[25] ));
 sg13g2_nand2_1 _09508_ (.Y(_01756_),
    .A(net2353),
    .B(net2461));
 sg13g2_mux4_1 _09509_ (.S0(net2365),
    .A0(net2460),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A2(net2462),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S1(net2480),
    .X(_01757_));
 sg13g2_inv_1 _09510_ (.Y(_01758_),
    .A(_01757_));
 sg13g2_mux2_1 _09511_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(net2366),
    .X(_01759_));
 sg13g2_mux2_1 _09512_ (.A0(net2464),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(net2366),
    .X(_01760_));
 sg13g2_mux2_1 _09513_ (.A0(_01759_),
    .A1(_01760_),
    .S(net2476),
    .X(_01761_));
 sg13g2_inv_1 _09514_ (.Y(_01762_),
    .A(_01761_));
 sg13g2_a21oi_1 _09515_ (.A1(net2470),
    .A2(_01762_),
    .Y(_01763_),
    .B1(net2227));
 sg13g2_o21ai_1 _09516_ (.B1(_01763_),
    .Y(_01764_),
    .A1(net2470),
    .A2(_01757_));
 sg13g2_mux2_1 _09517_ (.A0(net2465),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .S(net2366),
    .X(_01765_));
 sg13g2_mux2_1 _09518_ (.A0(net2466),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .S(net2367),
    .X(_01766_));
 sg13g2_mux2_1 _09519_ (.A0(_01765_),
    .A1(_01766_),
    .S(net2477),
    .X(_01767_));
 sg13g2_inv_1 _09520_ (.Y(_01768_),
    .A(_01767_));
 sg13g2_or2_1 _09521_ (.X(_01769_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .A(net2367));
 sg13g2_o21ai_1 _09522_ (.B1(_01769_),
    .Y(_01770_),
    .A1(net2353),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[28] ));
 sg13g2_mux2_1 _09523_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .S(net2370),
    .X(_01771_));
 sg13g2_nand2_1 _09524_ (.Y(_01772_),
    .A(net2478),
    .B(_01771_));
 sg13g2_o21ai_1 _09525_ (.B1(_01772_),
    .Y(_01773_),
    .A1(net2477),
    .A2(_01770_));
 sg13g2_a21oi_1 _09526_ (.A1(net2469),
    .A2(_01768_),
    .Y(_01774_),
    .B1(net2226));
 sg13g2_o21ai_1 _09527_ (.B1(_01774_),
    .Y(_01775_),
    .A1(net2469),
    .A2(_01773_));
 sg13g2_mux2_1 _09528_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(net2462),
    .S(net2362),
    .X(_01776_));
 sg13g2_or2_1 _09529_ (.X(_01777_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .A(net2362));
 sg13g2_o21ai_1 _09530_ (.B1(_01777_),
    .Y(_01778_),
    .A1(net2353),
    .A2(net2460));
 sg13g2_nor2_1 _09531_ (.A(net2476),
    .B(_01776_),
    .Y(_01779_));
 sg13g2_a21oi_1 _09532_ (.A1(net2476),
    .A2(_01778_),
    .Y(_01780_),
    .B1(_01779_));
 sg13g2_or2_1 _09533_ (.X(_01781_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A(net2366));
 sg13g2_o21ai_1 _09534_ (.B1(_01781_),
    .Y(_01782_),
    .A1(net2353),
    .A2(net2464));
 sg13g2_nor2_1 _09535_ (.A(net2477),
    .B(_01782_),
    .Y(_01783_));
 sg13g2_mux2_1 _09536_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .S(net2366),
    .X(_01784_));
 sg13g2_a21oi_1 _09537_ (.A1(net2477),
    .A2(_01784_),
    .Y(_01785_),
    .B1(_01783_));
 sg13g2_nand2_1 _09538_ (.Y(_01786_),
    .A(net2367),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[2] ));
 sg13g2_nand2_1 _09539_ (.Y(_01787_),
    .A(net2354),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[29] ));
 sg13g2_and2_1 _09540_ (.A(_01786_),
    .B(_01787_),
    .X(_01788_));
 sg13g2_nand2_1 _09541_ (.Y(_01789_),
    .A(net2367),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[3] ));
 sg13g2_o21ai_1 _09542_ (.B1(_01789_),
    .Y(_01790_),
    .A1(net2367),
    .A2(_01119_));
 sg13g2_nand2_1 _09543_ (.Y(_01791_),
    .A(net2479),
    .B(_01790_));
 sg13g2_o21ai_1 _09544_ (.B1(_01791_),
    .Y(_01792_),
    .A1(net2479),
    .A2(_01788_));
 sg13g2_mux2_1 _09545_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A1(net2465),
    .S(net2367),
    .X(_01793_));
 sg13g2_nand2_1 _09546_ (.Y(_01794_),
    .A(net2479),
    .B(_01793_));
 sg13g2_a21oi_1 _09547_ (.A1(net2354),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .Y(_01795_),
    .B1(_01714_));
 sg13g2_o21ai_1 _09548_ (.B1(_01794_),
    .Y(_01796_),
    .A1(net2479),
    .A2(_01795_));
 sg13g2_mux2_1 _09549_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(net2457),
    .S(net2362),
    .X(_01797_));
 sg13g2_mux2_1 _09550_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .S(net2364),
    .X(_01798_));
 sg13g2_mux2_1 _09551_ (.A0(_01797_),
    .A1(_01798_),
    .S(net2474),
    .X(_01799_));
 sg13g2_nor2_1 _09552_ (.A(net2331),
    .B(_01799_),
    .Y(_01800_));
 sg13g2_mux2_1 _09553_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .S(net2362),
    .X(_01801_));
 sg13g2_or2_1 _09554_ (.X(_01802_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A(net2362));
 sg13g2_o21ai_1 _09555_ (.B1(_01802_),
    .Y(_01803_),
    .A1(net2353),
    .A2(\i_tinyqv.cpu.i_core.i_shift.a[9] ));
 sg13g2_nor2_1 _09556_ (.A(net2475),
    .B(_01801_),
    .Y(_01804_));
 sg13g2_a21oi_1 _09557_ (.A1(net2475),
    .A2(_01803_),
    .Y(_01805_),
    .B1(_01804_));
 sg13g2_inv_1 _09558_ (.Y(_01806_),
    .A(_01805_));
 sg13g2_a21oi_1 _09559_ (.A1(net2332),
    .A2(_01806_),
    .Y(_01807_),
    .B1(_01800_));
 sg13g2_or2_1 _09560_ (.X(_01808_),
    .B(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A(net2364));
 sg13g2_o21ai_1 _09561_ (.B1(_01808_),
    .Y(_01809_),
    .A1(net2353),
    .A2(net2455));
 sg13g2_mux2_1 _09562_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .S(net2364),
    .X(_01810_));
 sg13g2_nand2_1 _09563_ (.Y(_01811_),
    .A(net2472),
    .B(_01810_));
 sg13g2_o21ai_1 _09564_ (.B1(_01811_),
    .Y(_01812_),
    .A1(net2472),
    .A2(_01809_));
 sg13g2_mux2_1 _09565_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(net2453),
    .S(net2363),
    .X(_01813_));
 sg13g2_mux2_1 _09566_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(net2452),
    .S(net2363),
    .X(_01814_));
 sg13g2_mux2_1 _09567_ (.A0(_01813_),
    .A1(_01814_),
    .S(net2473),
    .X(_01815_));
 sg13g2_inv_1 _09568_ (.Y(_01816_),
    .A(_01815_));
 sg13g2_a21oi_1 _09569_ (.A1(net2467),
    .A2(_01816_),
    .Y(_01817_),
    .B1(net2224));
 sg13g2_o21ai_1 _09570_ (.B1(_01817_),
    .Y(_01818_),
    .A1(net2471),
    .A2(_01812_));
 sg13g2_nand3_1 _09571_ (.B(_01764_),
    .C(_01775_),
    .A(_01754_),
    .Y(_01819_));
 sg13g2_a21oi_1 _09572_ (.A1(net2224),
    .A2(_01807_),
    .Y(_01820_),
    .B1(net2147));
 sg13g2_a21oi_1 _09573_ (.A1(_01818_),
    .A2(_01820_),
    .Y(_01821_),
    .B1(_01745_));
 sg13g2_mux4_1 _09574_ (.S0(net2467),
    .A0(_01738_),
    .A1(_01743_),
    .A2(_01750_),
    .A3(_01751_),
    .S1(net2227),
    .X(_01822_));
 sg13g2_nand2b_1 _09575_ (.Y(_01823_),
    .B(net2147),
    .A_N(_01822_));
 sg13g2_o21ai_1 _09576_ (.B1(net2227),
    .Y(_01824_),
    .A1(net2333),
    .A2(_01780_));
 sg13g2_a21o_1 _09577_ (.A2(_01785_),
    .A1(net2333),
    .B1(_01824_),
    .X(_01825_));
 sg13g2_mux2_1 _09578_ (.A0(_01792_),
    .A1(_01796_),
    .S(net2334),
    .X(_01826_));
 sg13g2_a21oi_1 _09579_ (.A1(net2226),
    .A2(_01826_),
    .Y(_01827_),
    .B1(net2147));
 sg13g2_a21oi_1 _09580_ (.A1(_01825_),
    .A2(_01827_),
    .Y(_01828_),
    .B1(_01744_));
 sg13g2_a221oi_1 _09581_ (.B2(_01828_),
    .C1(_01731_),
    .B1(_01823_),
    .A1(_01819_),
    .Y(_01829_),
    .A2(_01821_));
 sg13g2_nor2_1 _09582_ (.A(_01732_),
    .B(_01829_),
    .Y(_01830_));
 sg13g2_nor2_1 _09583_ (.A(net2354),
    .B(_01830_),
    .Y(_01831_));
 sg13g2_nand2b_2 _09584_ (.Y(_01832_),
    .B(_01715_),
    .A_N(_01410_));
 sg13g2_mux4_1 _09585_ (.S0(net2362),
    .A0(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A2(net2460),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S1(net2475),
    .X(_01833_));
 sg13g2_a21oi_1 _09586_ (.A1(_01755_),
    .A2(_01756_),
    .Y(_01834_),
    .B1(net2475));
 sg13g2_a21oi_1 _09587_ (.A1(net2480),
    .A2(_01759_),
    .Y(_01835_),
    .B1(_01834_));
 sg13g2_a21oi_1 _09588_ (.A1(net2468),
    .A2(_01835_),
    .Y(_01836_),
    .B1(net2224));
 sg13g2_o21ai_1 _09589_ (.B1(_01836_),
    .Y(_01837_),
    .A1(net2468),
    .A2(_01833_));
 sg13g2_nor2_1 _09590_ (.A(net2473),
    .B(_01742_),
    .Y(_01838_));
 sg13g2_a21oi_1 _09591_ (.A1(net2472),
    .A2(_01747_),
    .Y(_01839_),
    .B1(_01838_));
 sg13g2_mux4_1 _09592_ (.S0(net2363),
    .A0(net2457),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A2(net2458),
    .A3(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S1(net2474),
    .X(_01840_));
 sg13g2_mux2_1 _09593_ (.A0(_01839_),
    .A1(_01840_),
    .S(net2467),
    .X(_01841_));
 sg13g2_a21oi_1 _09594_ (.A1(net2225),
    .A2(_01841_),
    .Y(_01842_),
    .B1(_01753_));
 sg13g2_nand2_1 _09595_ (.Y(_01843_),
    .A(net2475),
    .B(_01801_));
 sg13g2_o21ai_1 _09596_ (.B1(_01843_),
    .Y(_01844_),
    .A1(net2475),
    .A2(_01778_));
 sg13g2_nor2_1 _09597_ (.A(net2475),
    .B(_01803_),
    .Y(_01845_));
 sg13g2_a21oi_1 _09598_ (.A1(net2475),
    .A2(_01797_),
    .Y(_01846_),
    .B1(_01845_));
 sg13g2_a21oi_1 _09599_ (.A1(net2468),
    .A2(_01846_),
    .Y(_01847_),
    .B1(net2224));
 sg13g2_o21ai_1 _09600_ (.B1(_01847_),
    .Y(_01848_),
    .A1(net2468),
    .A2(_01844_));
 sg13g2_nor2_1 _09601_ (.A(net2478),
    .B(_01790_),
    .Y(_01849_));
 sg13g2_a21oi_1 _09602_ (.A1(net2477),
    .A2(_01782_),
    .Y(_01850_),
    .B1(_01849_));
 sg13g2_and2_1 _09603_ (.A(net2480),
    .B(_01776_),
    .X(_01851_));
 sg13g2_a21oi_1 _09604_ (.A1(_01120_),
    .A2(_01784_),
    .Y(_01852_),
    .B1(_01851_));
 sg13g2_a21oi_1 _09605_ (.A1(net2470),
    .A2(_01852_),
    .Y(_01853_),
    .B1(net2227));
 sg13g2_o21ai_1 _09606_ (.B1(_01853_),
    .Y(_01854_),
    .A1(net2470),
    .A2(_01850_));
 sg13g2_nand3_1 _09607_ (.B(_01848_),
    .C(_01854_),
    .A(_01753_),
    .Y(_01855_));
 sg13g2_a21oi_1 _09608_ (.A1(_01837_),
    .A2(_01842_),
    .Y(_01856_),
    .B1(_01744_));
 sg13g2_nand2_1 _09609_ (.Y(_01857_),
    .A(_01855_),
    .B(_01856_));
 sg13g2_nand2b_1 _09610_ (.Y(_01858_),
    .B(net2477),
    .A_N(_01765_));
 sg13g2_o21ai_1 _09611_ (.B1(_01858_),
    .Y(_01859_),
    .A1(net2477),
    .A2(_01771_));
 sg13g2_nor2_1 _09612_ (.A(net2476),
    .B(_01760_),
    .Y(_01860_));
 sg13g2_a21oi_1 _09613_ (.A1(net2477),
    .A2(_01770_),
    .Y(_01861_),
    .B1(_01860_));
 sg13g2_a21oi_1 _09614_ (.A1(net2469),
    .A2(_01859_),
    .Y(_01862_),
    .B1(net2227));
 sg13g2_o21ai_1 _09615_ (.B1(_01862_),
    .Y(_01863_),
    .A1(net2470),
    .A2(_01861_));
 sg13g2_a21oi_1 _09616_ (.A1(net2469),
    .A2(_01720_),
    .Y(_01864_),
    .B1(net2226));
 sg13g2_nor2_1 _09617_ (.A(net2478),
    .B(_01766_),
    .Y(_01865_));
 sg13g2_a21oi_1 _09618_ (.A1(net2478),
    .A2(_01720_),
    .Y(_01866_),
    .B1(_01865_));
 sg13g2_o21ai_1 _09619_ (.B1(_01864_),
    .Y(_01867_),
    .A1(net2469),
    .A2(_01866_));
 sg13g2_nand3_1 _09620_ (.B(_01863_),
    .C(_01867_),
    .A(_01754_),
    .Y(_01868_));
 sg13g2_mux2_1 _09621_ (.A0(_01810_),
    .A1(_01813_),
    .S(net2473),
    .X(_01869_));
 sg13g2_nor2_1 _09622_ (.A(net2472),
    .B(_01798_),
    .Y(_01870_));
 sg13g2_a21oi_1 _09623_ (.A1(net2476),
    .A2(_01809_),
    .Y(_01871_),
    .B1(_01870_));
 sg13g2_mux2_1 _09624_ (.A0(_01869_),
    .A1(_01871_),
    .S(net2331),
    .X(_01872_));
 sg13g2_mux2_1 _09625_ (.A0(_01814_),
    .A1(_01734_),
    .S(net2473),
    .X(_01873_));
 sg13g2_nand2_1 _09626_ (.Y(_01874_),
    .A(net2472),
    .B(_01741_));
 sg13g2_o21ai_1 _09627_ (.B1(_01874_),
    .Y(_01875_),
    .A1(net2472),
    .A2(_01736_));
 sg13g2_inv_1 _09628_ (.Y(_01876_),
    .A(_01875_));
 sg13g2_a21oi_1 _09629_ (.A1(net2467),
    .A2(_01876_),
    .Y(_01877_),
    .B1(net2224));
 sg13g2_o21ai_1 _09630_ (.B1(_01877_),
    .Y(_01878_),
    .A1(net2467),
    .A2(_01873_));
 sg13g2_a21oi_1 _09631_ (.A1(net2225),
    .A2(_01872_),
    .Y(_01879_),
    .B1(net2147));
 sg13g2_a21oi_1 _09632_ (.A1(_01878_),
    .A2(_01879_),
    .Y(_01880_),
    .B1(_01745_));
 sg13g2_a21oi_1 _09633_ (.A1(_01868_),
    .A2(_01880_),
    .Y(_01881_),
    .B1(_01731_));
 sg13g2_a21oi_1 _09634_ (.A1(_01857_),
    .A2(_01881_),
    .Y(_01882_),
    .B1(_01732_));
 sg13g2_nor2_1 _09635_ (.A(net2368),
    .B(_01882_),
    .Y(_01883_));
 sg13g2_nor3_1 _09636_ (.A(_01831_),
    .B(_01832_),
    .C(_01883_),
    .Y(_01884_));
 sg13g2_nand2b_1 _09637_ (.Y(_01885_),
    .B(_01370_),
    .A_N(_01374_));
 sg13g2_nor2_1 _09638_ (.A(net2372),
    .B(net2374),
    .Y(_01886_));
 sg13g2_nor3_1 _09639_ (.A(net2369),
    .B(net2372),
    .C(net2374),
    .Y(_01887_));
 sg13g2_nand2_2 _09640_ (.Y(_01888_),
    .A(net2354),
    .B(_01886_));
 sg13g2_nand3b_1 _09641_ (.B(_01885_),
    .C(_01887_),
    .Y(_01889_),
    .A_N(_01375_));
 sg13g2_a21o_2 _09642_ (.A2(_01886_),
    .A1(net2369),
    .B1(_01194_),
    .X(_01890_));
 sg13g2_nand3_1 _09643_ (.B(net2371),
    .C(_01195_),
    .A(net2369),
    .Y(_01891_));
 sg13g2_a21oi_1 _09644_ (.A1(net2373),
    .A2(_01394_),
    .Y(_01892_),
    .B1(_01891_));
 sg13g2_a21oi_1 _09645_ (.A1(_01394_),
    .A2(_01890_),
    .Y(_01893_),
    .B1(_01892_));
 sg13g2_o21ai_1 _09646_ (.B1(_01889_),
    .Y(_01894_),
    .A1(_01393_),
    .A2(_01893_));
 sg13g2_a21oi_1 _09647_ (.A1(net2466),
    .A2(net1963),
    .Y(_01895_),
    .B1(\i_tinyqv.cpu.i_core.multiplier.accum[0] ));
 sg13g2_nor2_2 _09648_ (.A(net2369),
    .B(_01193_),
    .Y(_01896_));
 sg13g2_nand2_1 _09649_ (.Y(_01897_),
    .A(_01445_),
    .B(_01896_));
 sg13g2_nor4_1 _09650_ (.A(\i_tinyqv.cpu.alu_op[3] ),
    .B(net2233),
    .C(_01409_),
    .D(_01716_),
    .Y(_01898_));
 sg13g2_inv_1 _09651_ (.Y(_01899_),
    .A(_01898_));
 sg13g2_o21ai_1 _09652_ (.B1(_01899_),
    .Y(_01900_),
    .A1(_01895_),
    .A2(_01897_));
 sg13g2_nor3_1 _09653_ (.A(_01884_),
    .B(_01894_),
    .C(_01900_),
    .Y(_01901_));
 sg13g2_o21ai_1 _09654_ (.B1(net2323),
    .Y(_01902_),
    .A1(\i_tinyqv.cpu.i_core.cmp ),
    .A2(_01899_));
 sg13g2_o21ai_1 _09655_ (.B1(_01719_),
    .Y(_01903_),
    .A1(_01901_),
    .A2(_01902_));
 sg13g2_nor3_2 _09656_ (.A(\addr[27] ),
    .B(\addr[26] ),
    .C(\addr[25] ),
    .Y(_01904_));
 sg13g2_or3_1 _09657_ (.A(\addr[27] ),
    .B(\addr[26] ),
    .C(\addr[25] ),
    .X(_01905_));
 sg13g2_nand2_1 _09658_ (.Y(_01906_),
    .A(net2435),
    .B(_01437_));
 sg13g2_and2_1 _09659_ (.A(\i_tinyqv.cpu.data_write_n[1] ),
    .B(\i_tinyqv.cpu.data_write_n[0] ),
    .X(_01907_));
 sg13g2_nand2_2 _09660_ (.Y(_01908_),
    .A(\i_tinyqv.cpu.data_write_n[1] ),
    .B(\i_tinyqv.cpu.data_write_n[0] ));
 sg13g2_nor2_1 _09661_ (.A(net2300),
    .B(_01907_),
    .Y(_01909_));
 sg13g2_nor2_2 _09662_ (.A(net2426),
    .B(net2427),
    .Y(_01910_));
 sg13g2_nor3_2 _09663_ (.A(net2424),
    .B(net2426),
    .C(net2428),
    .Y(_01911_));
 sg13g2_nand2b_2 _09664_ (.Y(_01912_),
    .B(_01910_),
    .A_N(net2424));
 sg13g2_nor2_2 _09665_ (.A(net4137),
    .B(_01912_),
    .Y(_01913_));
 sg13g2_nand2_1 _09666_ (.Y(_01914_),
    .A(\i_tinyqv.cpu.data_read_n[1] ),
    .B(\i_tinyqv.cpu.data_read_n[0] ));
 sg13g2_and4_1 _09667_ (.A(\i_tinyqv.cpu.data_read_n[1] ),
    .B(\i_tinyqv.cpu.data_read_n[0] ),
    .C(_01909_),
    .D(_01913_),
    .X(_01915_));
 sg13g2_nor2_1 _09668_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .Y(_01916_));
 sg13g2_nand3_1 _09669_ (.B(_01909_),
    .C(_01916_),
    .A(\i_tinyqv.mem.data_stall ),
    .Y(_01917_));
 sg13g2_nor2b_1 _09670_ (.A(_01915_),
    .B_N(_01917_),
    .Y(_01918_));
 sg13g2_a21oi_1 _09671_ (.A1(_01906_),
    .A2(_01918_),
    .Y(_01919_),
    .B1(net2438));
 sg13g2_inv_1 _09672_ (.Y(_01920_),
    .A(net1998));
 sg13g2_nor2_2 _09673_ (.A(\addr[1] ),
    .B(\addr[0] ),
    .Y(_01921_));
 sg13g2_nor2_1 _09674_ (.A(\addr[7] ),
    .B(\addr[6] ),
    .Y(_01922_));
 sg13g2_nor4_1 _09675_ (.A(\addr[11] ),
    .B(\addr[10] ),
    .C(\addr[9] ),
    .D(\addr[8] ),
    .Y(_01923_));
 sg13g2_nand3_1 _09676_ (.B(_01922_),
    .C(_01923_),
    .A(_01921_),
    .Y(_01924_));
 sg13g2_nor2_1 _09677_ (.A(net2388),
    .B(_01924_),
    .Y(_01925_));
 sg13g2_inv_1 _09678_ (.Y(_01926_),
    .A(_01925_));
 sg13g2_nand3b_1 _09679_ (.B(_00928_),
    .C(\addr[27] ),
    .Y(_01927_),
    .A_N(\addr[24] ));
 sg13g2_nor4_1 _09680_ (.A(\addr[26] ),
    .B(\addr[25] ),
    .C(\addr[22] ),
    .D(_01927_),
    .Y(_01928_));
 sg13g2_nor3_1 _09681_ (.A(\addr[13] ),
    .B(\addr[12] ),
    .C(\addr[11] ),
    .Y(_01929_));
 sg13g2_nor4_1 _09682_ (.A(\addr[17] ),
    .B(\addr[16] ),
    .C(\addr[15] ),
    .D(\addr[14] ),
    .Y(_01930_));
 sg13g2_nor4_1 _09683_ (.A(\addr[21] ),
    .B(\addr[20] ),
    .C(\addr[19] ),
    .D(\addr[18] ),
    .Y(_01931_));
 sg13g2_and4_1 _09684_ (.A(_01928_),
    .B(_01929_),
    .C(_01930_),
    .D(_01931_),
    .X(_01932_));
 sg13g2_o21ai_1 _09685_ (.B1(_01932_),
    .Y(_01933_),
    .A1(net2386),
    .A2(_01924_));
 sg13g2_or2_1 _09686_ (.X(_01934_),
    .B(_01933_),
    .A(_01925_));
 sg13g2_nor2_1 _09687_ (.A(\addr[5] ),
    .B(_01924_),
    .Y(_01935_));
 sg13g2_o21ai_1 _09688_ (.B1(_01932_),
    .Y(_01936_),
    .A1(net2385),
    .A2(_01924_));
 sg13g2_inv_1 _09689_ (.Y(_01937_),
    .A(_01936_));
 sg13g2_or2_1 _09690_ (.X(_01938_),
    .B(_01936_),
    .A(_01935_));
 sg13g2_inv_1 _09691_ (.Y(_01939_),
    .A(_01938_));
 sg13g2_nor2_2 _09692_ (.A(_01934_),
    .B(_01938_),
    .Y(_01940_));
 sg13g2_or2_1 _09693_ (.X(_01941_),
    .B(_01938_),
    .A(_01934_));
 sg13g2_or4_1 _09694_ (.A(\i_peripherals.data_ready_r ),
    .B(net2302),
    .C(_01908_),
    .D(net1958),
    .X(_01942_));
 sg13g2_o21ai_1 _09695_ (.B1(_01942_),
    .Y(_01943_),
    .A1(net2300),
    .A2(net1998));
 sg13g2_a21oi_2 _09696_ (.B1(_01943_),
    .Y(_01944_),
    .A2(\addr[26] ),
    .A1(\addr[27] ));
 sg13g2_or2_1 _09697_ (.X(_01945_),
    .B(_01944_),
    .A(net3689));
 sg13g2_nand2_1 _09698_ (.Y(_01946_),
    .A(\addr[11] ),
    .B(\addr[8] ));
 sg13g2_nand4_1 _09699_ (.B(\addr[18] ),
    .C(\addr[17] ),
    .A(\addr[19] ),
    .Y(_01947_),
    .D(\addr[16] ));
 sg13g2_nand4_1 _09700_ (.B(\addr[14] ),
    .C(\addr[13] ),
    .A(\addr[15] ),
    .Y(_01948_),
    .D(\addr[12] ));
 sg13g2_nor4_2 _09701_ (.A(net2386),
    .B(_01946_),
    .C(_01947_),
    .Y(_01949_),
    .D(_01948_));
 sg13g2_nor2_2 _09702_ (.A(\addr[5] ),
    .B(\addr[4] ),
    .Y(_01950_));
 sg13g2_nand4_1 _09703_ (.B(\addr[9] ),
    .C(_01922_),
    .A(\addr[10] ),
    .Y(_01951_),
    .D(_01950_));
 sg13g2_nand4_1 _09704_ (.B(\addr[22] ),
    .C(\addr[21] ),
    .A(\addr[23] ),
    .Y(_01952_),
    .D(\addr[20] ));
 sg13g2_nand4_1 _09705_ (.B(\addr[26] ),
    .C(\addr[25] ),
    .A(\addr[27] ),
    .Y(_01953_),
    .D(\addr[24] ));
 sg13g2_nor3_1 _09706_ (.A(_01951_),
    .B(_01952_),
    .C(_01953_),
    .Y(_01954_));
 sg13g2_and2_1 _09707_ (.A(_01949_),
    .B(_01954_),
    .X(_01955_));
 sg13g2_nand2_2 _09708_ (.Y(_01956_),
    .A(_01949_),
    .B(_01954_));
 sg13g2_nor3_1 _09709_ (.A(net2234),
    .B(_01945_),
    .C(_01955_),
    .Y(_01957_));
 sg13g2_nor2_1 _09710_ (.A(net3732),
    .B(net2237),
    .Y(_01958_));
 sg13g2_nor2_1 _09711_ (.A(_01957_),
    .B(_01958_),
    .Y(_01959_));
 sg13g2_nand3_1 _09712_ (.B(_01403_),
    .C(_01959_),
    .A(\i_tinyqv.cpu.is_load ),
    .Y(_01960_));
 sg13g2_nand2_1 _09713_ (.Y(_01961_),
    .A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ));
 sg13g2_xnor2_1 _09714_ (.Y(_01962_),
    .A(\i_tinyqv.cpu.instr_len[2] ),
    .B(\i_tinyqv.cpu.pc[2] ));
 sg13g2_nand2_1 _09715_ (.Y(_01963_),
    .A(\i_tinyqv.cpu.instr_len[1] ),
    .B(\i_tinyqv.cpu.pc[1] ));
 sg13g2_o21ai_1 _09716_ (.B1(_01961_),
    .Y(_01964_),
    .A1(_01962_),
    .A2(_01963_));
 sg13g2_nand3_1 _09717_ (.B(net2418),
    .C(_01964_),
    .A(\i_tinyqv.cpu.instr_data_start[4] ),
    .Y(_01965_));
 sg13g2_nand4_1 _09718_ (.B(net2417),
    .C(net2418),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .Y(_01966_),
    .D(_01964_));
 sg13g2_nor2_2 _09719_ (.A(_00981_),
    .B(_01966_),
    .Y(_01967_));
 sg13g2_nand3_1 _09720_ (.B(net2416),
    .C(_01967_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .Y(_01968_));
 sg13g2_nor2_1 _09721_ (.A(_00980_),
    .B(_01968_),
    .Y(_01969_));
 sg13g2_nand3_1 _09722_ (.B(net2415),
    .C(_01969_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .Y(_01970_));
 sg13g2_nor2_1 _09723_ (.A(_00979_),
    .B(_01970_),
    .Y(_01971_));
 sg13g2_nand3_1 _09724_ (.B(net2414),
    .C(_01971_),
    .A(net2413),
    .Y(_01972_));
 sg13g2_nor2_1 _09725_ (.A(_00978_),
    .B(_01972_),
    .Y(_01973_));
 sg13g2_nand3_1 _09726_ (.B(net2412),
    .C(_01973_),
    .A(net2411),
    .Y(_01974_));
 sg13g2_nor2_1 _09727_ (.A(_00977_),
    .B(_01974_),
    .Y(_01975_));
 sg13g2_nand3_1 _09728_ (.B(net2410),
    .C(_01975_),
    .A(net2409),
    .Y(_01976_));
 sg13g2_a21o_1 _09729_ (.A2(_01975_),
    .A1(net2410),
    .B1(net2409),
    .X(_01977_));
 sg13g2_nand2_1 _09730_ (.Y(_01978_),
    .A(_01976_),
    .B(_01977_));
 sg13g2_xor2_1 _09731_ (.B(_01973_),
    .A(net2412),
    .X(_01979_));
 sg13g2_xnor2_1 _09732_ (.Y(_01980_),
    .A(\i_tinyqv.cpu.instr_data_start[12] ),
    .B(_01970_));
 sg13g2_a21o_1 _09733_ (.A2(_01967_),
    .A1(net2416),
    .B1(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(_01981_));
 sg13g2_and2_1 _09734_ (.A(_01968_),
    .B(_01981_),
    .X(_01982_));
 sg13g2_a21o_1 _09735_ (.A2(_01964_),
    .A1(net2418),
    .B1(net2417),
    .X(_01983_));
 sg13g2_and2_1 _09736_ (.A(_01965_),
    .B(_01983_),
    .X(_01984_));
 sg13g2_a22oi_1 _09737_ (.Y(_01985_),
    .B1(_01984_),
    .B2(net2318),
    .A2(_01982_),
    .A1(net2326));
 sg13g2_nor2_1 _09738_ (.A(net2375),
    .B(_01985_),
    .Y(_01986_));
 sg13g2_a221oi_1 _09739_ (.B2(_01346_),
    .C1(_01986_),
    .B1(_01980_),
    .A1(net2243),
    .Y(_01987_),
    .A2(_01979_));
 sg13g2_o21ai_1 _09740_ (.B1(_01987_),
    .Y(_01988_),
    .A1(_01207_),
    .A2(_01978_));
 sg13g2_nand2_1 _09741_ (.Y(_01989_),
    .A(_01423_),
    .B(_01988_));
 sg13g2_nand2b_2 _09742_ (.Y(_01990_),
    .B(_01418_),
    .A_N(_01886_));
 sg13g2_nor3_2 _09743_ (.A(\i_tinyqv.cpu.is_jal ),
    .B(\i_tinyqv.cpu.is_jalr ),
    .C(_01990_),
    .Y(_01991_));
 sg13g2_nor2_1 _09744_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .Y(_01992_));
 sg13g2_nand3b_1 _09745_ (.B(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .C(_01992_),
    .Y(_01993_),
    .A_N(net2439));
 sg13g2_inv_1 _09746_ (.Y(_01994_),
    .A(_01993_));
 sg13g2_nor3_1 _09747_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .Y(_01995_));
 sg13g2_nand2_2 _09748_ (.Y(_01996_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_nor3_1 _09749_ (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .C(_01996_),
    .Y(_01997_));
 sg13g2_nand2_1 _09750_ (.Y(_01998_),
    .A(_01995_),
    .B(_01997_));
 sg13g2_nand3_1 _09751_ (.B(_01995_),
    .C(_01997_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .Y(_01999_));
 sg13g2_or2_1 _09752_ (.X(_02000_),
    .B(_01999_),
    .A(_01993_));
 sg13g2_nand2_2 _09753_ (.Y(_02001_),
    .A(net2378),
    .B(_01199_));
 sg13g2_nor2_2 _09754_ (.A(net2319),
    .B(_02001_),
    .Y(_02002_));
 sg13g2_nand2_1 _09755_ (.Y(_02003_),
    .A(net2381),
    .B(net2375));
 sg13g2_nor2_2 _09756_ (.A(_02000_),
    .B(_02002_),
    .Y(_02004_));
 sg13g2_nand2_1 _09757_ (.Y(_02005_),
    .A(\i_tinyqv.cpu.i_core.mepc[0] ),
    .B(_02004_));
 sg13g2_nor4_1 _09758_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(_01070_),
    .C(net2439),
    .D(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .Y(_02006_));
 sg13g2_nor2b_2 _09759_ (.A(_01999_),
    .B_N(_02006_),
    .Y(_02007_));
 sg13g2_and2_1 _09760_ (.A(net2242),
    .B(_02007_),
    .X(_02008_));
 sg13g2_nand3b_1 _09761_ (.B(_01992_),
    .C(net2439),
    .Y(_02009_),
    .A_N(\i_tinyqv.cpu.i_core.imm_lo[0] ));
 sg13g2_nor2_1 _09762_ (.A(_01999_),
    .B(_02009_),
    .Y(_02010_));
 sg13g2_nor3_2 _09763_ (.A(net2233),
    .B(_01999_),
    .C(_02009_),
    .Y(_02011_));
 sg13g2_a22oi_1 _09764_ (.Y(_02012_),
    .B1(_02011_),
    .B2(\i_tinyqv.cpu.i_core.mcause[0] ),
    .A2(_02008_),
    .A1(\i_tinyqv.cpu.i_core.mip[0] ));
 sg13g2_nand2_1 _09765_ (.Y(_02013_),
    .A(_02005_),
    .B(_02012_));
 sg13g2_a22oi_1 _09766_ (.Y(_02014_),
    .B1(net2231),
    .B2(\i_tinyqv.cpu.i_core.mie[12] ),
    .A2(net2245),
    .A1(\i_tinyqv.cpu.i_core.mie[8] ));
 sg13g2_a22oi_1 _09767_ (.Y(_02015_),
    .B1(_01207_),
    .B2(_02014_),
    .A2(_01205_),
    .A1(_01020_));
 sg13g2_a21oi_1 _09768_ (.A1(\i_tinyqv.cpu.i_core.mie[0] ),
    .A2(net2242),
    .Y(_02016_),
    .B1(_02015_));
 sg13g2_nor2_2 _09769_ (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .B(_01998_),
    .Y(_02017_));
 sg13g2_nand2_2 _09770_ (.Y(_02018_),
    .A(_02006_),
    .B(_02017_));
 sg13g2_inv_1 _09771_ (.Y(_02019_),
    .A(_02018_));
 sg13g2_or2_1 _09772_ (.X(_02020_),
    .B(_02018_),
    .A(_02016_));
 sg13g2_nand2_1 _09773_ (.Y(_02021_),
    .A(_01994_),
    .B(_02017_));
 sg13g2_a22oi_1 _09774_ (.Y(_02022_),
    .B1(_02017_),
    .B2(_01994_),
    .A2(_02010_),
    .A1(\i_tinyqv.cpu.i_core.mcause[4] ));
 sg13g2_nand2b_1 _09775_ (.Y(_02023_),
    .B(_01343_),
    .A_N(_02022_));
 sg13g2_nand3b_1 _09776_ (.B(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .C(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .Y(_02024_),
    .A_N(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_nor3_1 _09777_ (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .C(_02024_),
    .Y(_02025_));
 sg13g2_nand2_2 _09778_ (.Y(_02026_),
    .A(_01995_),
    .B(_02025_));
 sg13g2_nor2_2 _09779_ (.A(_02009_),
    .B(_02026_),
    .Y(_02027_));
 sg13g2_nor3_1 _09780_ (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .C(_01996_),
    .Y(_02028_));
 sg13g2_nand2_1 _09781_ (.Y(_02029_),
    .A(_01992_),
    .B(_02028_));
 sg13g2_nand3_1 _09782_ (.B(net2439),
    .C(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .A(net2338),
    .Y(_02030_));
 sg13g2_nor4_1 _09783_ (.A(_01364_),
    .B(_02024_),
    .C(_02029_),
    .D(_02030_),
    .Y(_02031_));
 sg13g2_a21oi_1 _09784_ (.A1(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .A2(_02027_),
    .Y(_02032_),
    .B1(_02031_));
 sg13g2_nor2_2 _09785_ (.A(_01993_),
    .B(_02026_),
    .Y(_02033_));
 sg13g2_nor4_1 _09786_ (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .C(net2439),
    .D(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .Y(_02034_));
 sg13g2_nor2b_2 _09787_ (.A(_02026_),
    .B_N(_02034_),
    .Y(_02035_));
 sg13g2_a22oi_1 _09788_ (.Y(_02036_),
    .B1(_02035_),
    .B2(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .A2(_02033_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[3] ));
 sg13g2_nand4_1 _09789_ (.B(_02023_),
    .C(_02032_),
    .A(_02020_),
    .Y(_02037_),
    .D(_02036_));
 sg13g2_o21ai_1 _09790_ (.B1(_01991_),
    .Y(_02038_),
    .A1(_02013_),
    .A2(_02037_));
 sg13g2_nand3_1 _09791_ (.B(_01989_),
    .C(_02038_),
    .A(_01426_),
    .Y(_02039_));
 sg13g2_o21ai_1 _09792_ (.B1(_02039_),
    .Y(_02040_),
    .A1(_01367_),
    .A2(_01426_));
 sg13g2_a21oi_1 _09793_ (.A1(_00946_),
    .A2(net2380),
    .Y(_02041_),
    .B1(net2376));
 sg13g2_nor2_2 _09794_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(_02041_),
    .Y(_02042_));
 sg13g2_or2_1 _09795_ (.X(_02043_),
    .B(_02041_),
    .A(\i_tinyqv.cpu.i_core.mem_op[1] ));
 sg13g2_a21oi_2 _09796_ (.B1(_01960_),
    .Y(_02044_),
    .A2(_02042_),
    .A1(\i_tinyqv.cpu.i_core.load_top_bit ));
 sg13g2_nand2b_1 _09797_ (.Y(_02045_),
    .B(net3945),
    .A_N(net3882));
 sg13g2_or2_1 _09798_ (.X(_02046_),
    .B(_02045_),
    .A(_01920_));
 sg13g2_nand2b_1 _09799_ (.Y(_02047_),
    .B(net1954),
    .A_N(\i_tinyqv.mem.qspi_data_buf[8] ));
 sg13g2_o21ai_1 _09800_ (.B1(_02047_),
    .Y(_02048_),
    .A1(net2423),
    .A2(net1953));
 sg13g2_mux2_1 _09801_ (.A0(net2420),
    .A1(\i_tinyqv.mem.qspi_data_buf[12] ),
    .S(net1953),
    .X(_02049_));
 sg13g2_a21oi_1 _09802_ (.A1(net2382),
    .A2(_02049_),
    .Y(_02050_),
    .B1(net2301));
 sg13g2_o21ai_1 _09803_ (.B1(_02050_),
    .Y(_02051_),
    .A1(net2382),
    .A2(_02048_));
 sg13g2_a21oi_1 _09804_ (.A1(\addr[5] ),
    .A2(_01932_),
    .Y(_02052_),
    .B1(_01937_));
 sg13g2_nand4_1 _09805_ (.B(_01925_),
    .C(_01932_),
    .A(net2386),
    .Y(_02053_),
    .D(_02052_));
 sg13g2_nand2_2 _09806_ (.Y(_02054_),
    .A(_01934_),
    .B(_02053_));
 sg13g2_inv_2 _09807_ (.Y(_02055_),
    .A(_02054_));
 sg13g2_nor2b_1 _09808_ (.A(net2382),
    .B_N(\i_peripherals.data_out[8] ),
    .Y(_02056_));
 sg13g2_a21oi_1 _09809_ (.A1(\i_peripherals.data_out[12] ),
    .A2(net2383),
    .Y(_02057_),
    .B1(_02056_));
 sg13g2_o21ai_1 _09810_ (.B1(_02054_),
    .Y(_02058_),
    .A1(net1958),
    .A2(_02057_));
 sg13g2_nand3_1 _09811_ (.B(_02051_),
    .C(_02058_),
    .A(net2379),
    .Y(_02059_));
 sg13g2_nor3_1 _09812_ (.A(\i_tinyqv.mem.data_txn_len[1] ),
    .B(\i_tinyqv.mem.data_txn_len[0] ),
    .C(_01920_),
    .Y(_02060_));
 sg13g2_a21oi_1 _09813_ (.A1(net2423),
    .A2(net1952),
    .Y(_02061_),
    .B1(net2300));
 sg13g2_o21ai_1 _09814_ (.B1(_02061_),
    .Y(_02062_),
    .A1(_01117_),
    .A2(net1952));
 sg13g2_nand3_1 _09815_ (.B(_01932_),
    .C(_01936_),
    .A(\addr[5] ),
    .Y(_02063_));
 sg13g2_or3_1 _09816_ (.A(net3365),
    .B(\i_debug_uart_tx.fsm_state[2] ),
    .C(net3182),
    .X(_02064_));
 sg13g2_nor2_2 _09817_ (.A(net3988),
    .B(_02064_),
    .Y(_02065_));
 sg13g2_nand2b_2 _09818_ (.Y(_02066_),
    .B(_01023_),
    .A_N(_02064_));
 sg13g2_nand4_1 _09819_ (.B(_01932_),
    .C(_01935_),
    .A(net2385),
    .Y(_02067_),
    .D(_02066_));
 sg13g2_nand3b_1 _09820_ (.B(_02063_),
    .C(_02067_),
    .Y(_02068_),
    .A_N(_01934_));
 sg13g2_a21oi_1 _09821_ (.A1(\i_peripherals.data_out[0] ),
    .A2(_01939_),
    .Y(_02069_),
    .B1(_02068_));
 sg13g2_nor2_1 _09822_ (.A(_01199_),
    .B(_02069_),
    .Y(_02070_));
 sg13g2_a21oi_1 _09823_ (.A1(net2420),
    .A2(net1952),
    .Y(_02071_),
    .B1(net2301));
 sg13g2_o21ai_1 _09824_ (.B1(_02071_),
    .Y(_02072_),
    .A1(_01118_),
    .A2(net1952));
 sg13g2_nor2_2 _09825_ (.A(_01934_),
    .B(_02063_),
    .Y(_02073_));
 sg13g2_a221oi_1 _09826_ (.B2(\time_limit[4] ),
    .C1(_02055_),
    .B1(_02073_),
    .A1(\i_peripherals.data_out[4] ),
    .Y(_02074_),
    .A2(_01940_));
 sg13g2_nor2_1 _09827_ (.A(net2317),
    .B(_02074_),
    .Y(_02075_));
 sg13g2_a22oi_1 _09828_ (.Y(_02076_),
    .B1(_02072_),
    .B2(_02075_),
    .A2(_02070_),
    .A1(_02062_));
 sg13g2_a21oi_1 _09829_ (.A1(_02059_),
    .A2(_02076_),
    .Y(_02077_),
    .B1(net2376));
 sg13g2_mux2_1 _09830_ (.A0(\i_tinyqv.mem.qspi_data_buf[24] ),
    .A1(net2422),
    .S(net1997),
    .X(_02078_));
 sg13g2_mux2_1 _09831_ (.A0(\i_tinyqv.mem.qspi_data_buf[28] ),
    .A1(net2420),
    .S(net1997),
    .X(_02079_));
 sg13g2_a22oi_1 _09832_ (.Y(_02080_),
    .B1(net2314),
    .B2(\i_tinyqv.mem.data_from_read[16] ),
    .A2(net2322),
    .A1(\i_tinyqv.mem.data_from_read[20] ));
 sg13g2_nand2_1 _09833_ (.Y(_02081_),
    .A(net2302),
    .B(_02080_));
 sg13g2_a221oi_1 _09834_ (.B2(net2310),
    .C1(_02081_),
    .B1(_02079_),
    .A1(net2327),
    .Y(_02082_),
    .A2(_02078_));
 sg13g2_a22oi_1 _09835_ (.Y(_02083_),
    .B1(net2316),
    .B2(\i_peripherals.data_out[16] ),
    .A2(net2327),
    .A1(\i_peripherals.data_out[24] ));
 sg13g2_a22oi_1 _09836_ (.Y(_02084_),
    .B1(net2310),
    .B2(\i_peripherals.data_out[28] ),
    .A2(net2322),
    .A1(\i_peripherals.data_out[20] ));
 sg13g2_a21oi_2 _09837_ (.B1(net1958),
    .Y(_02085_),
    .A2(_02084_),
    .A1(_02083_));
 sg13g2_o21ai_1 _09838_ (.B1(net2377),
    .Y(_02086_),
    .A1(_02055_),
    .A2(_02085_));
 sg13g2_nor2_1 _09839_ (.A(_02082_),
    .B(_02086_),
    .Y(_02087_));
 sg13g2_nor2_1 _09840_ (.A(net2387),
    .B(_01113_),
    .Y(_02088_));
 sg13g2_a21oi_2 _09841_ (.B1(_02088_),
    .Y(_02089_),
    .A2(\i_tinyqv.cpu.i_timer.mtimecmp[4] ),
    .A1(\addr[2] ));
 sg13g2_a21oi_1 _09842_ (.A1(_01955_),
    .A2(_02089_),
    .Y(_02090_),
    .B1(_02042_));
 sg13g2_o21ai_1 _09843_ (.B1(_02090_),
    .Y(_02091_),
    .A1(_02077_),
    .A2(_02087_));
 sg13g2_a22oi_1 _09844_ (.Y(_02092_),
    .B1(_02044_),
    .B2(_02091_),
    .A2(_02040_),
    .A1(_01960_));
 sg13g2_mux2_1 _09845_ (.A0(_02092_),
    .A1(_01903_),
    .S(_01713_),
    .X(\debug_rd[0] ));
 sg13g2_and3_1 _09846_ (.X(_02093_),
    .A(_01408_),
    .B(_01427_),
    .C(_01990_));
 sg13g2_nor3_1 _09847_ (.A(net2370),
    .B(net2504),
    .C(_01193_),
    .Y(_02094_));
 sg13g2_a22oi_1 _09848_ (.Y(_02095_),
    .B1(_02094_),
    .B2(_01713_),
    .A2(_02093_),
    .A1(_01960_));
 sg13g2_and3_2 _09849_ (.X(_02096_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(net2502),
    .C(net2501));
 sg13g2_nand3_1 _09850_ (.B(net1891),
    .C(_02096_),
    .A(net2500),
    .Y(_02097_));
 sg13g2_mux2_1 _09851_ (.A0(net1874),
    .A1(net3650),
    .S(_02097_),
    .X(_00041_));
 sg13g2_a21o_1 _09852_ (.A2(_01377_),
    .A1(_01376_),
    .B1(_01888_),
    .X(_02098_));
 sg13g2_a21oi_1 _09853_ (.A1(net2373),
    .A2(_01396_),
    .Y(_02099_),
    .B1(_01891_));
 sg13g2_a21oi_1 _09854_ (.A1(_01396_),
    .A2(_01890_),
    .Y(_02100_),
    .B1(_02099_));
 sg13g2_a21o_1 _09855_ (.A2(_01330_),
    .A1(_01312_),
    .B1(_02100_),
    .X(_02101_));
 sg13g2_o21ai_1 _09856_ (.B1(_02101_),
    .Y(_02102_),
    .A1(_01378_),
    .A2(_02098_));
 sg13g2_nor2_2 _09857_ (.A(_01194_),
    .B(_01898_),
    .Y(_02103_));
 sg13g2_mux2_1 _09858_ (.A0(_01743_),
    .A1(_01750_),
    .S(net2467),
    .X(_02104_));
 sg13g2_nand2b_1 _09859_ (.Y(_02105_),
    .B(net2331),
    .A_N(_01751_));
 sg13g2_a21oi_1 _09860_ (.A1(net2471),
    .A2(_01758_),
    .Y(_02106_),
    .B1(net2224));
 sg13g2_a221oi_1 _09861_ (.B2(_02106_),
    .C1(_01753_),
    .B1(_02105_),
    .A1(net2225),
    .Y(_02107_),
    .A2(_02104_));
 sg13g2_o21ai_1 _09862_ (.B1(net2226),
    .Y(_02108_),
    .A1(net2469),
    .A2(_01792_));
 sg13g2_a21oi_1 _09863_ (.A1(net2470),
    .A2(_01785_),
    .Y(_02109_),
    .B1(_02108_));
 sg13g2_o21ai_1 _09864_ (.B1(net2227),
    .Y(_02110_),
    .A1(net2468),
    .A2(_01780_));
 sg13g2_a21oi_1 _09865_ (.A1(net2468),
    .A2(_01806_),
    .Y(_02111_),
    .B1(_02110_));
 sg13g2_nor3_1 _09866_ (.A(net2147),
    .B(_02109_),
    .C(_02111_),
    .Y(_02112_));
 sg13g2_nor3_1 _09867_ (.A(_01744_),
    .B(_02107_),
    .C(_02112_),
    .Y(_02113_));
 sg13g2_o21ai_1 _09868_ (.B1(net2226),
    .Y(_02114_),
    .A1(net2334),
    .A2(_01773_));
 sg13g2_a21o_1 _09869_ (.A2(_01762_),
    .A1(net2334),
    .B1(_02114_),
    .X(_02115_));
 sg13g2_o21ai_1 _09870_ (.B1(_01864_),
    .Y(_02116_),
    .A1(net2469),
    .A2(_01767_));
 sg13g2_nand3_1 _09871_ (.B(_02115_),
    .C(_02116_),
    .A(_01754_),
    .Y(_02117_));
 sg13g2_nor2_1 _09872_ (.A(net2467),
    .B(_01799_),
    .Y(_02118_));
 sg13g2_nor2_1 _09873_ (.A(net2227),
    .B(_02118_),
    .Y(_02119_));
 sg13g2_o21ai_1 _09874_ (.B1(_02119_),
    .Y(_02120_),
    .A1(net2332),
    .A2(_01812_));
 sg13g2_nor2_1 _09875_ (.A(net2332),
    .B(_01738_),
    .Y(_02121_));
 sg13g2_a21oi_1 _09876_ (.A1(net2331),
    .A2(_01816_),
    .Y(_02122_),
    .B1(_02121_));
 sg13g2_a21oi_1 _09877_ (.A1(net2227),
    .A2(_02122_),
    .Y(_02123_),
    .B1(net2147));
 sg13g2_a21oi_1 _09878_ (.A1(_02120_),
    .A2(_02123_),
    .Y(_02124_),
    .B1(_01745_));
 sg13g2_a21o_1 _09879_ (.A2(_02124_),
    .A1(_02117_),
    .B1(_01731_),
    .X(_02125_));
 sg13g2_o21ai_1 _09880_ (.B1(_01733_),
    .Y(_02126_),
    .A1(_02113_),
    .A2(_02125_));
 sg13g2_o21ai_1 _09881_ (.B1(_01739_),
    .Y(_02127_),
    .A1(net2334),
    .A2(_01866_));
 sg13g2_a21o_1 _09882_ (.A2(_01859_),
    .A1(net2334),
    .B1(_02127_),
    .X(_02128_));
 sg13g2_nor2_1 _09883_ (.A(net2333),
    .B(_01861_),
    .Y(_02129_));
 sg13g2_a21oi_1 _09884_ (.A1(net2333),
    .A2(_01835_),
    .Y(_02130_),
    .B1(_02129_));
 sg13g2_nand2_1 _09885_ (.Y(_02131_),
    .A(net2469),
    .B(_01850_));
 sg13g2_nand2_1 _09886_ (.Y(_02132_),
    .A(net2480),
    .B(_01788_));
 sg13g2_o21ai_1 _09887_ (.B1(_02132_),
    .Y(_02133_),
    .A1(net2479),
    .A2(_01793_));
 sg13g2_nor2_1 _09888_ (.A(net2331),
    .B(_01871_),
    .Y(_02134_));
 sg13g2_a21oi_1 _09889_ (.A1(net2331),
    .A2(_01846_),
    .Y(_02135_),
    .B1(_02134_));
 sg13g2_nor2_1 _09890_ (.A(net2467),
    .B(_01869_),
    .Y(_02136_));
 sg13g2_nor2_1 _09891_ (.A(net2224),
    .B(_02136_),
    .Y(_02137_));
 sg13g2_o21ai_1 _09892_ (.B1(_02137_),
    .Y(_02138_),
    .A1(net2331),
    .A2(_01873_));
 sg13g2_a21oi_1 _09893_ (.A1(_01740_),
    .A2(_02130_),
    .Y(_02139_),
    .B1(_01753_));
 sg13g2_a21oi_1 _09894_ (.A1(net2225),
    .A2(_02135_),
    .Y(_02140_),
    .B1(net2147));
 sg13g2_a221oi_1 _09895_ (.B2(_02138_),
    .C1(_01745_),
    .B1(_02140_),
    .A1(_02128_),
    .Y(_02141_),
    .A2(_02139_));
 sg13g2_mux4_1 _09896_ (.S0(net2224),
    .A0(_01833_),
    .A1(_01839_),
    .A2(_01840_),
    .A3(_01875_),
    .S1(net2331),
    .X(_02142_));
 sg13g2_a21oi_1 _09897_ (.A1(net2333),
    .A2(_01852_),
    .Y(_02143_),
    .B1(net2225));
 sg13g2_o21ai_1 _09898_ (.B1(_02143_),
    .Y(_02144_),
    .A1(net2333),
    .A2(_01844_));
 sg13g2_o21ai_1 _09899_ (.B1(_02131_),
    .Y(_02145_),
    .A1(net2470),
    .A2(_02133_));
 sg13g2_a21oi_1 _09900_ (.A1(net2226),
    .A2(_02145_),
    .Y(_02146_),
    .B1(net2147));
 sg13g2_a21oi_1 _09901_ (.A1(_02144_),
    .A2(_02146_),
    .Y(_02147_),
    .B1(_01744_));
 sg13g2_o21ai_1 _09902_ (.B1(_02147_),
    .Y(_02148_),
    .A1(_01753_),
    .A2(_02142_));
 sg13g2_nand2b_1 _09903_ (.Y(_02149_),
    .B(_02148_),
    .A_N(_01731_));
 sg13g2_o21ai_1 _09904_ (.B1(_01733_),
    .Y(_02150_),
    .A1(_02141_),
    .A2(_02149_));
 sg13g2_a21o_1 _09905_ (.A2(_02150_),
    .A1(net2368),
    .B1(_01832_),
    .X(_02151_));
 sg13g2_a21oi_1 _09906_ (.A1(net2354),
    .A2(_02126_),
    .Y(_02152_),
    .B1(_02151_));
 sg13g2_xor2_1 _09907_ (.B(_01445_),
    .A(_01444_),
    .X(_02153_));
 sg13g2_nor2_1 _09908_ (.A(_01896_),
    .B(_02102_),
    .Y(_02154_));
 sg13g2_a21oi_1 _09909_ (.A1(_01896_),
    .A2(_02153_),
    .Y(_02155_),
    .B1(_02154_));
 sg13g2_o21ai_1 _09910_ (.B1(_02103_),
    .Y(_02156_),
    .A1(_02152_),
    .A2(_02155_));
 sg13g2_nand3_1 _09911_ (.B(net2465),
    .C(_01717_),
    .A(net2368),
    .Y(_02157_));
 sg13g2_and2_1 _09912_ (.A(_02156_),
    .B(_02157_),
    .X(_02158_));
 sg13g2_or2_1 _09913_ (.X(_02159_),
    .B(_01976_),
    .A(_00976_));
 sg13g2_xnor2_1 _09914_ (.Y(_02160_),
    .A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(_01976_));
 sg13g2_a21o_1 _09915_ (.A2(_01973_),
    .A1(net2412),
    .B1(net2411),
    .X(_02161_));
 sg13g2_nand2_1 _09916_ (.Y(_02162_),
    .A(_01974_),
    .B(_02161_));
 sg13g2_inv_1 _09917_ (.Y(_02163_),
    .A(_02162_));
 sg13g2_xnor2_1 _09918_ (.Y(_02164_),
    .A(net2414),
    .B(_01971_));
 sg13g2_xnor2_1 _09919_ (.Y(_02165_),
    .A(_00980_),
    .B(_01968_));
 sg13g2_xor2_1 _09920_ (.B(_01965_),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(_02166_));
 sg13g2_xnor2_1 _09921_ (.Y(_02167_),
    .A(\i_tinyqv.cpu.instr_len[1] ),
    .B(\i_tinyqv.cpu.pc[1] ));
 sg13g2_a22oi_1 _09922_ (.Y(_02168_),
    .B1(_02167_),
    .B2(net2313),
    .A2(_02166_),
    .A1(net2318));
 sg13g2_nand2_1 _09923_ (.Y(_02169_),
    .A(net2336),
    .B(_02168_));
 sg13g2_a221oi_1 _09924_ (.B2(net2326),
    .C1(_02169_),
    .B1(_02165_),
    .A1(net2309),
    .Y(_02170_),
    .A2(_02164_));
 sg13g2_a221oi_1 _09925_ (.B2(net2243),
    .C1(_02170_),
    .B1(_02163_),
    .A1(net2244),
    .Y(_02171_),
    .A2(_02160_));
 sg13g2_a21oi_1 _09926_ (.A1(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .A2(_02035_),
    .Y(_02172_),
    .B1(_02031_));
 sg13g2_mux2_1 _09927_ (.A0(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .S(net2228),
    .X(_02173_));
 sg13g2_a22oi_1 _09928_ (.Y(_02174_),
    .B1(_02033_),
    .B2(_02173_),
    .A2(_02027_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[1] ));
 sg13g2_a22oi_1 _09929_ (.Y(_02175_),
    .B1(_02011_),
    .B2(\i_tinyqv.cpu.i_core.mcause[1] ),
    .A2(_02004_),
    .A1(\i_tinyqv.cpu.i_core.mepc[1] ));
 sg13g2_a221oi_1 _09930_ (.B2(\i_tinyqv.cpu.i_core.mie[13] ),
    .C1(_01205_),
    .B1(net2231),
    .A1(\i_tinyqv.cpu.i_core.mie[9] ),
    .Y(_02176_),
    .A2(net2245));
 sg13g2_nand2b_1 _09931_ (.Y(_02177_),
    .B(net2241),
    .A_N(\i_tinyqv.cpu.i_core.mie[1] ));
 sg13g2_o21ai_1 _09932_ (.B1(_02177_),
    .Y(_02178_),
    .A1(\i_tinyqv.cpu.i_core.mie[5] ),
    .A2(_01207_));
 sg13g2_nor3_1 _09933_ (.A(_02018_),
    .B(_02176_),
    .C(_02178_),
    .Y(_02179_));
 sg13g2_a21oi_1 _09934_ (.A1(\i_tinyqv.cpu.i_core.mip[1] ),
    .A2(_02008_),
    .Y(_02180_),
    .B1(_02179_));
 sg13g2_nand4_1 _09935_ (.B(_02174_),
    .C(_02175_),
    .A(_02172_),
    .Y(_02181_),
    .D(_02180_));
 sg13g2_a21oi_1 _09936_ (.A1(_01991_),
    .A2(_02181_),
    .Y(_02182_),
    .B1(_01425_));
 sg13g2_o21ai_1 _09937_ (.B1(_02182_),
    .Y(_02183_),
    .A1(_01424_),
    .A2(_02171_));
 sg13g2_o21ai_1 _09938_ (.B1(_02183_),
    .Y(_02184_),
    .A1(_01318_),
    .A2(_01426_));
 sg13g2_nand2_1 _09939_ (.Y(_02185_),
    .A(_01960_),
    .B(_02184_));
 sg13g2_o21ai_1 _09940_ (.B1(net2314),
    .Y(_02186_),
    .A1(\i_tinyqv.cpu.instr_data_in[1] ),
    .A2(net1952));
 sg13g2_a21oi_1 _09941_ (.A1(_01124_),
    .A2(net1951),
    .Y(_02187_),
    .B1(_02186_));
 sg13g2_o21ai_1 _09942_ (.B1(net2320),
    .Y(_02188_),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .A2(net1952));
 sg13g2_a21oi_1 _09943_ (.A1(_01125_),
    .A2(net1952),
    .Y(_02189_),
    .B1(_02188_));
 sg13g2_o21ai_1 _09944_ (.B1(net2325),
    .Y(_02190_),
    .A1(\i_tinyqv.cpu.instr_data_in[9] ),
    .A2(net1954));
 sg13g2_a21oi_1 _09945_ (.A1(_01126_),
    .A2(net1954),
    .Y(_02191_),
    .B1(_02190_));
 sg13g2_o21ai_1 _09946_ (.B1(net2310),
    .Y(_02192_),
    .A1(\i_tinyqv.cpu.instr_data_in[13] ),
    .A2(net1954));
 sg13g2_a21oi_1 _09947_ (.A1(_01127_),
    .A2(net1954),
    .Y(_02193_),
    .B1(_02192_));
 sg13g2_nor3_1 _09948_ (.A(_02187_),
    .B(_02189_),
    .C(_02191_),
    .Y(_02194_));
 sg13g2_nor2_1 _09949_ (.A(net2301),
    .B(_02193_),
    .Y(_02195_));
 sg13g2_mux2_1 _09950_ (.A0(\i_peripherals.data_out[1] ),
    .A1(\i_peripherals.data_out[5] ),
    .S(net2383),
    .X(_02196_));
 sg13g2_nand2_1 _09951_ (.Y(_02197_),
    .A(net2383),
    .B(_01109_));
 sg13g2_a22oi_1 _09952_ (.Y(_02198_),
    .B1(_02197_),
    .B2(_02073_),
    .A2(_02196_),
    .A1(_01940_));
 sg13g2_nor2_1 _09953_ (.A(net2379),
    .B(_02198_),
    .Y(_02199_));
 sg13g2_a22oi_1 _09954_ (.Y(_02200_),
    .B1(net2310),
    .B2(\i_peripherals.data_out[13] ),
    .A2(net2327),
    .A1(\i_peripherals.data_out[9] ));
 sg13g2_o21ai_1 _09955_ (.B1(_02054_),
    .Y(_02201_),
    .A1(net1958),
    .A2(_02200_));
 sg13g2_o21ai_1 _09956_ (.B1(net2337),
    .Y(_02202_),
    .A1(_02199_),
    .A2(_02201_));
 sg13g2_a21oi_1 _09957_ (.A1(_02194_),
    .A2(_02195_),
    .Y(_02203_),
    .B1(_02202_));
 sg13g2_a21oi_1 _09958_ (.A1(_01125_),
    .A2(net1996),
    .Y(_02204_),
    .B1(net2307));
 sg13g2_o21ai_1 _09959_ (.B1(_02204_),
    .Y(_02205_),
    .A1(\i_tinyqv.mem.qspi_data_buf[29] ),
    .A2(net1996));
 sg13g2_a21oi_1 _09960_ (.A1(_01124_),
    .A2(net1996),
    .Y(_02206_),
    .B1(net2324));
 sg13g2_o21ai_1 _09961_ (.B1(_02206_),
    .Y(_02207_),
    .A1(\i_tinyqv.mem.qspi_data_buf[25] ),
    .A2(net1996));
 sg13g2_a22oi_1 _09962_ (.Y(_02208_),
    .B1(net2316),
    .B2(\i_tinyqv.mem.data_from_read[17] ),
    .A2(net2322),
    .A1(\i_tinyqv.mem.data_from_read[21] ));
 sg13g2_nand4_1 _09963_ (.B(_02205_),
    .C(_02207_),
    .A(net2302),
    .Y(_02209_),
    .D(_02208_));
 sg13g2_a22oi_1 _09964_ (.Y(_02210_),
    .B1(net2322),
    .B2(\i_peripherals.data_out[21] ),
    .A2(net2327),
    .A1(\i_peripherals.data_out[25] ));
 sg13g2_a22oi_1 _09965_ (.Y(_02211_),
    .B1(net2310),
    .B2(\i_peripherals.data_out[29] ),
    .A2(net2316),
    .A1(\i_peripherals.data_out[17] ));
 sg13g2_a21oi_1 _09966_ (.A1(_02210_),
    .A2(_02211_),
    .Y(_02212_),
    .B1(net1958));
 sg13g2_o21ai_1 _09967_ (.B1(net2377),
    .Y(_02213_),
    .A1(_02055_),
    .A2(_02212_));
 sg13g2_nor2b_1 _09968_ (.A(_02213_),
    .B_N(_02209_),
    .Y(_02214_));
 sg13g2_nor3_2 _09969_ (.A(_01955_),
    .B(_02203_),
    .C(_02214_),
    .Y(_02215_));
 sg13g2_nand2_1 _09970_ (.Y(_02216_),
    .A(net2387),
    .B(\i_tinyqv.cpu.i_timer.mtimecmp[5] ));
 sg13g2_o21ai_1 _09971_ (.B1(_02216_),
    .Y(_02217_),
    .A1(net2387),
    .A2(_01112_));
 sg13g2_o21ai_1 _09972_ (.B1(_02043_),
    .Y(_02218_),
    .A1(_01956_),
    .A2(_02217_));
 sg13g2_o21ai_1 _09973_ (.B1(_02044_),
    .Y(_02219_),
    .A1(_02215_),
    .A2(_02218_));
 sg13g2_a21oi_1 _09974_ (.A1(_02185_),
    .A2(_02219_),
    .Y(_02220_),
    .B1(_01713_));
 sg13g2_a21oi_2 _09975_ (.B1(_02220_),
    .Y(\debug_rd[1] ),
    .A2(_02158_),
    .A1(_01713_));
 sg13g2_mux2_1 _09976_ (.A0(net1872),
    .A1(net3755),
    .S(_02097_),
    .X(_00042_));
 sg13g2_nor3_1 _09977_ (.A(_01332_),
    .B(_01378_),
    .C(_01380_),
    .Y(_02221_));
 sg13g2_nor3_1 _09978_ (.A(_01381_),
    .B(_01888_),
    .C(_02221_),
    .Y(_02222_));
 sg13g2_nand2_1 _09979_ (.Y(_02223_),
    .A(net2373),
    .B(_01390_));
 sg13g2_nor2_1 _09980_ (.A(_01389_),
    .B(_01891_),
    .Y(_02224_));
 sg13g2_a221oi_1 _09981_ (.B2(_02224_),
    .C1(_02222_),
    .B1(_02223_),
    .A1(_01391_),
    .Y(_02225_),
    .A2(_01890_));
 sg13g2_or2_1 _09982_ (.X(_02226_),
    .B(_01457_),
    .A(_01446_));
 sg13g2_nand3_1 _09983_ (.B(_01896_),
    .C(_02226_),
    .A(_01458_),
    .Y(_02227_));
 sg13g2_nand3_1 _09984_ (.B(_02225_),
    .C(_02227_),
    .A(_01832_),
    .Y(_02228_));
 sg13g2_and2_1 _09985_ (.A(net2368),
    .B(_02126_),
    .X(_02229_));
 sg13g2_a21oi_1 _09986_ (.A1(_00924_),
    .A2(_02150_),
    .Y(_02230_),
    .B1(_02229_));
 sg13g2_o21ai_1 _09987_ (.B1(_02103_),
    .Y(_02231_),
    .A1(_01832_),
    .A2(_02230_));
 sg13g2_nand2b_1 _09988_ (.Y(_02232_),
    .B(_02228_),
    .A_N(_02231_));
 sg13g2_o21ai_1 _09989_ (.B1(_02232_),
    .Y(_02233_),
    .A1(_01718_),
    .A2(_01786_));
 sg13g2_nor2_1 _09990_ (.A(_00975_),
    .B(_02159_),
    .Y(_02234_));
 sg13g2_xnor2_1 _09991_ (.Y(_02235_),
    .A(_00975_),
    .B(_02159_));
 sg13g2_xnor2_1 _09992_ (.Y(_02236_),
    .A(\i_tinyqv.cpu.instr_data_start[18] ),
    .B(_01974_));
 sg13g2_a21o_1 _09993_ (.A2(_01971_),
    .A1(net2414),
    .B1(net4136),
    .X(_02237_));
 sg13g2_nand2_2 _09994_ (.Y(_02238_),
    .A(_01972_),
    .B(_02237_));
 sg13g2_xor2_1 _09995_ (.B(_01969_),
    .A(net2415),
    .X(_02239_));
 sg13g2_xnor2_1 _09996_ (.Y(_02240_),
    .A(_00981_),
    .B(_01966_));
 sg13g2_xnor2_1 _09997_ (.Y(_02241_),
    .A(_01962_),
    .B(_01963_));
 sg13g2_or2_1 _09998_ (.X(_02242_),
    .B(_02241_),
    .A(_01199_));
 sg13g2_o21ai_1 _09999_ (.B1(_02242_),
    .Y(_02243_),
    .A1(net2317),
    .A2(_02240_));
 sg13g2_a21oi_1 _10000_ (.A1(net2326),
    .A2(_02239_),
    .Y(_02244_),
    .B1(_02243_));
 sg13g2_o21ai_1 _10001_ (.B1(_02244_),
    .Y(_02245_),
    .A1(net2307),
    .A2(_02238_));
 sg13g2_a22oi_1 _10002_ (.Y(_02246_),
    .B1(_02245_),
    .B2(net2337),
    .A2(_02236_),
    .A1(net2243));
 sg13g2_o21ai_1 _10003_ (.B1(_02246_),
    .Y(_02247_),
    .A1(_01207_),
    .A2(_02235_));
 sg13g2_nand2_2 _10004_ (.Y(_02248_),
    .A(_02017_),
    .B(_02034_));
 sg13g2_inv_1 _10005_ (.Y(_02249_),
    .A(_02248_));
 sg13g2_nor2_1 _10006_ (.A(net2233),
    .B(_02248_),
    .Y(_02250_));
 sg13g2_nor3_1 _10007_ (.A(_00074_),
    .B(net2233),
    .C(_02248_),
    .Y(_02251_));
 sg13g2_a221oi_1 _10008_ (.B2(\i_tinyqv.cpu.i_core.mcause[2] ),
    .C1(_02251_),
    .B1(_02011_),
    .A1(\i_peripherals.i_uart.uart_rx_buffered ),
    .Y(_02252_),
    .A2(_02008_));
 sg13g2_a21oi_1 _10009_ (.A1(net2233),
    .A2(net2228),
    .Y(_02253_),
    .B1(_02021_));
 sg13g2_a21oi_1 _10010_ (.A1(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .A2(_02027_),
    .Y(_02254_),
    .B1(_02253_));
 sg13g2_mux2_1 _10011_ (.A0(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .A1(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .S(net2228),
    .X(_02255_));
 sg13g2_a22oi_1 _10012_ (.Y(_02256_),
    .B1(_02255_),
    .B2(_02033_),
    .A2(_02035_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[2] ));
 sg13g2_a221oi_1 _10013_ (.B2(\i_tinyqv.cpu.i_core.mie[14] ),
    .C1(_01205_),
    .B1(net2231),
    .A1(\i_tinyqv.cpu.i_core.mie[10] ),
    .Y(_02257_),
    .A2(net2245));
 sg13g2_nand2b_1 _10014_ (.Y(_02258_),
    .B(net2241),
    .A_N(\i_tinyqv.cpu.i_core.mie[2] ));
 sg13g2_o21ai_1 _10015_ (.B1(_02258_),
    .Y(_02259_),
    .A1(\i_tinyqv.cpu.i_core.mie[6] ),
    .A2(_01207_));
 sg13g2_nor3_1 _10016_ (.A(_02018_),
    .B(_02257_),
    .C(_02259_),
    .Y(_02260_));
 sg13g2_a21oi_1 _10017_ (.A1(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A2(_02004_),
    .Y(_02261_),
    .B1(_02260_));
 sg13g2_nand4_1 _10018_ (.B(_02254_),
    .C(_02256_),
    .A(_02252_),
    .Y(_02262_),
    .D(_02261_));
 sg13g2_a22oi_1 _10019_ (.Y(_02263_),
    .B1(_02262_),
    .B2(_01991_),
    .A2(_02247_),
    .A1(_01423_));
 sg13g2_nand2_1 _10020_ (.Y(_02264_),
    .A(_01426_),
    .B(_02263_));
 sg13g2_o21ai_1 _10021_ (.B1(_02264_),
    .Y(_02265_),
    .A1(_01282_),
    .A2(_01426_));
 sg13g2_mux2_1 _10022_ (.A0(\i_tinyqv.cpu.instr_data_in[14] ),
    .A1(\i_tinyqv.mem.qspi_data_buf[14] ),
    .S(net1954),
    .X(_02266_));
 sg13g2_a21oi_1 _10023_ (.A1(net2310),
    .A2(_02266_),
    .Y(_02267_),
    .B1(net2300));
 sg13g2_o21ai_1 _10024_ (.B1(net2328),
    .Y(_02268_),
    .A1(\i_tinyqv.cpu.instr_data_in[10] ),
    .A2(net1953));
 sg13g2_a21oi_1 _10025_ (.A1(_01130_),
    .A2(net1953),
    .Y(_02269_),
    .B1(_02268_));
 sg13g2_o21ai_1 _10026_ (.B1(net2321),
    .Y(_02270_),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .A2(net1951));
 sg13g2_a21oi_1 _10027_ (.A1(_01129_),
    .A2(net1951),
    .Y(_02271_),
    .B1(_02270_));
 sg13g2_o21ai_1 _10028_ (.B1(net2315),
    .Y(_02272_),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .A2(net1951));
 sg13g2_a21oi_1 _10029_ (.A1(net2330),
    .A2(net1951),
    .Y(_02273_),
    .B1(_02272_));
 sg13g2_nor3_1 _10030_ (.A(_02269_),
    .B(_02271_),
    .C(_02273_),
    .Y(_02274_));
 sg13g2_nand2_1 _10031_ (.Y(_02275_),
    .A(\i_peripherals.data_out[6] ),
    .B(_01940_));
 sg13g2_nor2b_2 _10032_ (.A(_01934_),
    .B_N(_02052_),
    .Y(_02276_));
 sg13g2_a22oi_1 _10033_ (.Y(_02277_),
    .B1(_02276_),
    .B2(\gpio_out_sel[6] ),
    .A2(_02073_),
    .A1(\time_limit[6] ));
 sg13g2_nand3_1 _10034_ (.B(_02275_),
    .C(_02277_),
    .A(_02053_),
    .Y(_02278_));
 sg13g2_nand2_1 _10035_ (.Y(_02279_),
    .A(net2319),
    .B(_02278_));
 sg13g2_a22oi_1 _10036_ (.Y(_02280_),
    .B1(_02073_),
    .B2(\time_limit[2] ),
    .A2(_01940_),
    .A1(\i_peripherals.data_out[2] ));
 sg13g2_inv_1 _10037_ (.Y(_02281_),
    .A(_02280_));
 sg13g2_a22oi_1 _10038_ (.Y(_02282_),
    .B1(net2311),
    .B2(\i_peripherals.data_out[14] ),
    .A2(net2327),
    .A1(\i_peripherals.data_out[10] ));
 sg13g2_o21ai_1 _10039_ (.B1(_02054_),
    .Y(_02283_),
    .A1(net1958),
    .A2(_02282_));
 sg13g2_a21oi_1 _10040_ (.A1(net2314),
    .A2(_02281_),
    .Y(_02284_),
    .B1(_02283_));
 sg13g2_a221oi_1 _10041_ (.B2(_02284_),
    .C1(net2376),
    .B1(_02279_),
    .A1(_02267_),
    .Y(_02285_),
    .A2(_02274_));
 sg13g2_a21oi_1 _10042_ (.A1(net2330),
    .A2(net1996),
    .Y(_02286_),
    .B1(net2324));
 sg13g2_o21ai_1 _10043_ (.B1(_02286_),
    .Y(_02287_),
    .A1(\i_tinyqv.mem.qspi_data_buf[26] ),
    .A2(net1996));
 sg13g2_a21oi_1 _10044_ (.A1(_01129_),
    .A2(net1996),
    .Y(_02288_),
    .B1(net2307));
 sg13g2_o21ai_1 _10045_ (.B1(_02288_),
    .Y(_02289_),
    .A1(\i_tinyqv.mem.qspi_data_buf[30] ),
    .A2(net1996));
 sg13g2_a22oi_1 _10046_ (.Y(_02290_),
    .B1(net2316),
    .B2(\i_tinyqv.mem.data_from_read[18] ),
    .A2(net2322),
    .A1(\i_tinyqv.mem.data_from_read[22] ));
 sg13g2_nand4_1 _10047_ (.B(_02287_),
    .C(_02289_),
    .A(net2302),
    .Y(_02291_),
    .D(_02290_));
 sg13g2_a22oi_1 _10048_ (.Y(_02292_),
    .B1(net2322),
    .B2(\i_peripherals.data_out[22] ),
    .A2(net2327),
    .A1(\i_peripherals.data_out[26] ));
 sg13g2_a22oi_1 _10049_ (.Y(_02293_),
    .B1(net2311),
    .B2(\i_peripherals.data_out[30] ),
    .A2(net2316),
    .A1(\i_peripherals.data_out[18] ));
 sg13g2_and2_1 _10050_ (.A(_02292_),
    .B(_02293_),
    .X(_02294_));
 sg13g2_o21ai_1 _10051_ (.B1(_02054_),
    .Y(_02295_),
    .A1(net1958),
    .A2(_02294_));
 sg13g2_nand3_1 _10052_ (.B(_02291_),
    .C(_02295_),
    .A(net2377),
    .Y(_02296_));
 sg13g2_nand2_1 _10053_ (.Y(_02297_),
    .A(_01956_),
    .B(_02296_));
 sg13g2_nor2b_1 _10054_ (.A(net2387),
    .B_N(\i_tinyqv.cpu.i_timer.i_mtime.data[2] ),
    .Y(_02298_));
 sg13g2_a21oi_2 _10055_ (.B1(_02298_),
    .Y(_02299_),
    .A2(\i_tinyqv.cpu.i_timer.mtimecmp[6] ),
    .A1(net2387));
 sg13g2_a21oi_1 _10056_ (.A1(_01955_),
    .A2(_02299_),
    .Y(_02300_),
    .B1(_02042_));
 sg13g2_o21ai_1 _10057_ (.B1(_02300_),
    .Y(_02301_),
    .A1(_02285_),
    .A2(_02297_));
 sg13g2_a221oi_1 _10058_ (.B2(_02044_),
    .C1(_01713_),
    .B1(_02301_),
    .A1(_01960_),
    .Y(_02302_),
    .A2(_02265_));
 sg13g2_a21o_2 _10059_ (.A2(_02233_),
    .A1(_01713_),
    .B1(_02302_),
    .X(\debug_rd[2] ));
 sg13g2_mux2_1 _10060_ (.A0(net1867),
    .A1(net4017),
    .S(_02097_),
    .X(_00043_));
 sg13g2_o21ai_1 _10061_ (.B1(net2309),
    .Y(_02303_),
    .A1(net2419),
    .A2(net1953));
 sg13g2_a21oi_1 _10062_ (.A1(_01136_),
    .A2(net1953),
    .Y(_02304_),
    .B1(_02303_));
 sg13g2_o21ai_1 _10063_ (.B1(net2315),
    .Y(_02305_),
    .A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .A2(net1951));
 sg13g2_a21oi_1 _10064_ (.A1(_01133_),
    .A2(net1951),
    .Y(_02306_),
    .B1(_02305_));
 sg13g2_mux2_1 _10065_ (.A0(\i_tinyqv.cpu.instr_data_in[7] ),
    .A1(net2419),
    .S(net1951),
    .X(_02307_));
 sg13g2_a21oi_1 _10066_ (.A1(net2321),
    .A2(_02307_),
    .Y(_02308_),
    .B1(_02306_));
 sg13g2_o21ai_1 _10067_ (.B1(net2328),
    .Y(_02309_),
    .A1(\i_tinyqv.cpu.instr_data_in[11] ),
    .A2(net1953));
 sg13g2_a21oi_1 _10068_ (.A1(_01135_),
    .A2(net1953),
    .Y(_02310_),
    .B1(_02309_));
 sg13g2_nor3_1 _10069_ (.A(net2301),
    .B(_02304_),
    .C(_02310_),
    .Y(_02311_));
 sg13g2_a22oi_1 _10070_ (.Y(_02312_),
    .B1(_02276_),
    .B2(\gpio_out_sel[7] ),
    .A2(_01940_),
    .A1(\i_peripherals.data_out[7] ));
 sg13g2_nor2_1 _10071_ (.A(net2317),
    .B(_02312_),
    .Y(_02313_));
 sg13g2_nand3_1 _10072_ (.B(net2315),
    .C(_02073_),
    .A(\time_limit[3] ),
    .Y(_02314_));
 sg13g2_nand2_1 _10073_ (.Y(_02315_),
    .A(\i_peripherals.data_out[15] ),
    .B(net2311));
 sg13g2_a22oi_1 _10074_ (.Y(_02316_),
    .B1(net2316),
    .B2(\i_peripherals.data_out[3] ),
    .A2(net2328),
    .A1(\i_peripherals.data_out[11] ));
 sg13g2_a21o_1 _10075_ (.A2(_02316_),
    .A1(_02315_),
    .B1(net1958),
    .X(_02317_));
 sg13g2_nand3_1 _10076_ (.B(_02314_),
    .C(_02317_),
    .A(_02054_),
    .Y(_02318_));
 sg13g2_o21ai_1 _10077_ (.B1(net2337),
    .Y(_02319_),
    .A1(_02313_),
    .A2(_02318_));
 sg13g2_a21o_1 _10078_ (.A2(_02311_),
    .A1(_02308_),
    .B1(_02319_),
    .X(_02320_));
 sg13g2_mux2_1 _10079_ (.A0(\i_tinyqv.mem.qspi_data_buf[31] ),
    .A1(net2419),
    .S(net1997),
    .X(_02321_));
 sg13g2_o21ai_1 _10080_ (.B1(net2327),
    .Y(_02322_),
    .A1(\i_tinyqv.mem.qspi_data_buf[27] ),
    .A2(net1998));
 sg13g2_a21oi_1 _10081_ (.A1(_01133_),
    .A2(net1997),
    .Y(_02323_),
    .B1(_02322_));
 sg13g2_a221oi_1 _10082_ (.B2(\i_tinyqv.mem.data_from_read[19] ),
    .C1(net2300),
    .B1(net2314),
    .A1(\i_tinyqv.mem.data_from_read[23] ),
    .Y(_02324_),
    .A2(net2321));
 sg13g2_a21oi_1 _10083_ (.A1(net2310),
    .A2(_02321_),
    .Y(_02325_),
    .B1(_02323_));
 sg13g2_a22oi_1 _10084_ (.Y(_02326_),
    .B1(net2311),
    .B2(\i_peripherals.data_out[31] ),
    .A2(net2327),
    .A1(\i_peripherals.data_out[27] ));
 sg13g2_a22oi_1 _10085_ (.Y(_02327_),
    .B1(net2316),
    .B2(\i_peripherals.data_out[19] ),
    .A2(net2322),
    .A1(\i_peripherals.data_out[23] ));
 sg13g2_a21oi_1 _10086_ (.A1(_02326_),
    .A2(_02327_),
    .Y(_02328_),
    .B1(_01941_));
 sg13g2_o21ai_1 _10087_ (.B1(net2377),
    .Y(_02329_),
    .A1(_02055_),
    .A2(_02328_));
 sg13g2_a21oi_1 _10088_ (.A1(_02324_),
    .A2(_02325_),
    .Y(_02330_),
    .B1(_02329_));
 sg13g2_nor2_1 _10089_ (.A(_01955_),
    .B(_02330_),
    .Y(_02331_));
 sg13g2_nor2b_1 _10090_ (.A(net2387),
    .B_N(\i_tinyqv.cpu.i_timer.i_mtime.data[3] ),
    .Y(_02332_));
 sg13g2_a21oi_2 _10091_ (.B1(_02332_),
    .Y(_02333_),
    .A2(\i_tinyqv.cpu.i_timer.mtimecmp[7] ),
    .A1(net2387));
 sg13g2_a22oi_1 _10092_ (.Y(_02334_),
    .B1(_02333_),
    .B2(_01955_),
    .A2(_02331_),
    .A1(_02320_));
 sg13g2_nand2_1 _10093_ (.Y(_02335_),
    .A(_02043_),
    .B(_02334_));
 sg13g2_xnor2_1 _10094_ (.Y(_02336_),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .B(_02234_));
 sg13g2_xor2_1 _10095_ (.B(_01975_),
    .A(net2410),
    .X(_02337_));
 sg13g2_xnor2_1 _10096_ (.Y(_02338_),
    .A(_00978_),
    .B(_01972_));
 sg13g2_xor2_1 _10097_ (.B(_01967_),
    .A(net2416),
    .X(_02339_));
 sg13g2_inv_1 _10098_ (.Y(_02340_),
    .A(_02339_));
 sg13g2_xor2_1 _10099_ (.B(_01964_),
    .A(net4149),
    .X(_02341_));
 sg13g2_o21ai_1 _10100_ (.B1(net2336),
    .Y(_02342_),
    .A1(_01199_),
    .A2(_02341_));
 sg13g2_a21oi_1 _10101_ (.A1(net2318),
    .A2(_02340_),
    .Y(_02343_),
    .B1(_02342_));
 sg13g2_a21o_1 _10102_ (.A2(_01969_),
    .A1(net2415),
    .B1(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(_02344_));
 sg13g2_nand2_1 _10103_ (.Y(_02345_),
    .A(_01970_),
    .B(_02344_));
 sg13g2_a22oi_1 _10104_ (.Y(_02346_),
    .B1(_02345_),
    .B2(net2326),
    .A2(_02338_),
    .A1(net2309));
 sg13g2_a22oi_1 _10105_ (.Y(_02347_),
    .B1(_02343_),
    .B2(_02346_),
    .A2(_02337_),
    .A1(net2243));
 sg13g2_o21ai_1 _10106_ (.B1(_02347_),
    .Y(_02348_),
    .A1(_01207_),
    .A2(_02336_));
 sg13g2_nand2_1 _10107_ (.Y(_02349_),
    .A(_01423_),
    .B(_02348_));
 sg13g2_a22oi_1 _10108_ (.Y(_02350_),
    .B1(net2231),
    .B2(\i_tinyqv.cpu.i_core.mie[15] ),
    .A2(net2245),
    .A1(\i_tinyqv.cpu.i_core.mie[11] ));
 sg13g2_a22oi_1 _10109_ (.Y(_02351_),
    .B1(_01207_),
    .B2(_02350_),
    .A2(_01205_),
    .A1(_01021_));
 sg13g2_a21oi_1 _10110_ (.A1(\i_tinyqv.cpu.i_core.mie[3] ),
    .A2(net2242),
    .Y(_02352_),
    .B1(_02351_));
 sg13g2_o21ai_1 _10111_ (.B1(_02019_),
    .Y(_02353_),
    .A1(\i_tinyqv.cpu.i_core.mie[16] ),
    .A2(_01344_));
 sg13g2_a22oi_1 _10112_ (.Y(_02354_),
    .B1(_02249_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .A2(_02007_),
    .A1(\i_tinyqv.cpu.i_core.mip[16] ));
 sg13g2_nand2b_1 _10113_ (.Y(_02355_),
    .B(_01343_),
    .A_N(_02354_));
 sg13g2_a22oi_1 _10114_ (.Y(_02356_),
    .B1(_02353_),
    .B2(_02355_),
    .A2(_02352_),
    .A1(_01344_));
 sg13g2_and2_1 _10115_ (.A(\i_tinyqv.cpu.i_core.mcause[5] ),
    .B(net2231),
    .X(_02357_));
 sg13g2_a22oi_1 _10116_ (.Y(_02358_),
    .B1(_02357_),
    .B2(_02010_),
    .A2(_02035_),
    .A1(\i_tinyqv.cpu.i_core.cycle_count[3] ));
 sg13g2_nand2_1 _10117_ (.Y(_02359_),
    .A(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .B(net2228));
 sg13g2_o21ai_1 _10118_ (.B1(_02359_),
    .Y(_02360_),
    .A1(_01066_),
    .A2(net2228));
 sg13g2_a22oi_1 _10119_ (.Y(_02361_),
    .B1(_02033_),
    .B2(_02360_),
    .A2(_02027_),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.data[3] ));
 sg13g2_or3_1 _10120_ (.A(net3982),
    .B(net3532),
    .C(net2884),
    .X(_02362_));
 sg13g2_nor2_2 _10121_ (.A(\i_peripherals.i_uart.i_uart_tx.fsm_state[0] ),
    .B(_02362_),
    .Y(_02363_));
 sg13g2_nand2b_2 _10122_ (.Y(_02364_),
    .B(_01039_),
    .A_N(_02362_));
 sg13g2_a22oi_1 _10123_ (.Y(_02365_),
    .B1(_02008_),
    .B2(_02363_),
    .A2(_02004_),
    .A1(\i_tinyqv.cpu.i_core.mepc[3] ));
 sg13g2_a22oi_1 _10124_ (.Y(_02366_),
    .B1(_02250_),
    .B2(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .A2(_02011_),
    .A1(\i_tinyqv.cpu.i_core.mcause[3] ));
 sg13g2_nand4_1 _10125_ (.B(_02361_),
    .C(_02365_),
    .A(_02358_),
    .Y(_02367_),
    .D(_02366_));
 sg13g2_o21ai_1 _10126_ (.B1(_01991_),
    .Y(_02368_),
    .A1(_02356_),
    .A2(_02367_));
 sg13g2_nand3_1 _10127_ (.B(_02349_),
    .C(_02368_),
    .A(_01426_),
    .Y(_02369_));
 sg13g2_o21ai_1 _10128_ (.B1(_02369_),
    .Y(_02370_),
    .A1(_01223_),
    .A2(_01426_));
 sg13g2_a22oi_1 _10129_ (.Y(_02371_),
    .B1(_02370_),
    .B2(_01960_),
    .A2(_02335_),
    .A1(_02044_));
 sg13g2_nand2_1 _10130_ (.Y(_02372_),
    .A(_01458_),
    .B(_01474_));
 sg13g2_nand3b_1 _10131_ (.B(_01896_),
    .C(_02372_),
    .Y(_02373_),
    .A_N(_01475_));
 sg13g2_nand2_1 _10132_ (.Y(_02374_),
    .A(_01384_),
    .B(_01887_));
 sg13g2_a21oi_1 _10133_ (.A1(_01382_),
    .A2(_01383_),
    .Y(_02375_),
    .B1(_02374_));
 sg13g2_o21ai_1 _10134_ (.B1(net2373),
    .Y(_02376_),
    .A1(_01212_),
    .A2(_01256_));
 sg13g2_a21oi_1 _10135_ (.A1(_01212_),
    .A2(_01256_),
    .Y(_02377_),
    .B1(_01891_));
 sg13g2_a221oi_1 _10136_ (.B2(_02377_),
    .C1(_02375_),
    .B1(_02376_),
    .A1(_01392_),
    .Y(_02378_),
    .A2(_01890_));
 sg13g2_nand3_1 _10137_ (.B(_02373_),
    .C(_02378_),
    .A(_01832_),
    .Y(_02379_));
 sg13g2_a21o_1 _10138_ (.A2(_01882_),
    .A1(net2368),
    .B1(_01832_),
    .X(_02380_));
 sg13g2_a21o_1 _10139_ (.A2(_01830_),
    .A1(_00924_),
    .B1(_02380_),
    .X(_02381_));
 sg13g2_nand3_1 _10140_ (.B(_02379_),
    .C(_02381_),
    .A(_02103_),
    .Y(_02382_));
 sg13g2_o21ai_1 _10141_ (.B1(_02382_),
    .Y(_02383_),
    .A1(_01718_),
    .A2(_01789_));
 sg13g2_mux2_1 _10142_ (.A0(_02371_),
    .A1(_02383_),
    .S(_01713_),
    .X(\debug_rd[3] ));
 sg13g2_mux2_1 _10143_ (.A0(net1853),
    .A1(net3999),
    .S(_02097_),
    .X(_00044_));
 sg13g2_nor2b_2 _10144_ (.A(net2502),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .Y(_02384_));
 sg13g2_nand4_1 _10145_ (.B(net2500),
    .C(net1891),
    .A(net2501),
    .Y(_02385_),
    .D(_02384_));
 sg13g2_mux2_1 _10146_ (.A0(net1874),
    .A1(net3620),
    .S(_02385_),
    .X(_00037_));
 sg13g2_mux2_1 _10147_ (.A0(net1873),
    .A1(net3795),
    .S(_02385_),
    .X(_00038_));
 sg13g2_mux2_1 _10148_ (.A0(net1867),
    .A1(net3771),
    .S(_02385_),
    .X(_00039_));
 sg13g2_mux2_1 _10149_ (.A0(net1853),
    .A1(net3746),
    .S(_02385_),
    .X(_00040_));
 sg13g2_nor2b_2 _10150_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B_N(net2502),
    .Y(_02386_));
 sg13g2_nand4_1 _10151_ (.B(net2500),
    .C(net1891),
    .A(net2501),
    .Y(_02387_),
    .D(_02386_));
 sg13g2_mux2_1 _10152_ (.A0(net1875),
    .A1(net3902),
    .S(_02387_),
    .X(_00033_));
 sg13g2_mux2_1 _10153_ (.A0(net1872),
    .A1(net4065),
    .S(_02387_),
    .X(_00034_));
 sg13g2_mux2_1 _10154_ (.A0(net1867),
    .A1(net3936),
    .S(_02387_),
    .X(_00035_));
 sg13g2_mux2_1 _10155_ (.A0(net1854),
    .A1(net3633),
    .S(_02387_),
    .X(_00036_));
 sg13g2_nor2_1 _10156_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(net2502),
    .Y(_02388_));
 sg13g2_and4_1 _10157_ (.A(net2501),
    .B(net2500),
    .C(net1891),
    .D(_02388_),
    .X(_02389_));
 sg13g2_mux2_1 _10158_ (.A0(net3596),
    .A1(net1874),
    .S(_02389_),
    .X(_00029_));
 sg13g2_mux2_1 _10159_ (.A0(net3682),
    .A1(net1872),
    .S(_02389_),
    .X(_00030_));
 sg13g2_mux2_1 _10160_ (.A0(net3670),
    .A1(net1867),
    .S(_02389_),
    .X(_00031_));
 sg13g2_mux2_1 _10161_ (.A0(net3725),
    .A1(net1853),
    .S(_02389_),
    .X(_00032_));
 sg13g2_nand2_1 _10162_ (.Y(_02390_),
    .A(net2500),
    .B(net1891));
 sg13g2_nor2_2 _10163_ (.A(net2501),
    .B(_02390_),
    .Y(_02391_));
 sg13g2_nand3_1 _10164_ (.B(net2502),
    .C(_02391_),
    .A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .Y(_02392_));
 sg13g2_mux2_1 _10165_ (.A0(net1874),
    .A1(net3802),
    .S(_02392_),
    .X(_00025_));
 sg13g2_mux2_1 _10166_ (.A0(net1872),
    .A1(net4026),
    .S(_02392_),
    .X(_00026_));
 sg13g2_mux2_1 _10167_ (.A0(net1867),
    .A1(net4025),
    .S(_02392_),
    .X(_00027_));
 sg13g2_mux2_1 _10168_ (.A0(net1853),
    .A1(net3928),
    .S(_02392_),
    .X(_00028_));
 sg13g2_nand2_2 _10169_ (.Y(_02393_),
    .A(_02384_),
    .B(_02391_));
 sg13g2_mux2_1 _10170_ (.A0(net1874),
    .A1(net3542),
    .S(_02393_),
    .X(_00021_));
 sg13g2_mux2_1 _10171_ (.A0(net1873),
    .A1(net3971),
    .S(_02393_),
    .X(_00022_));
 sg13g2_mux2_1 _10172_ (.A0(net1868),
    .A1(net3826),
    .S(_02393_),
    .X(_00023_));
 sg13g2_mux2_1 _10173_ (.A0(net1853),
    .A1(net4001),
    .S(_02393_),
    .X(_00024_));
 sg13g2_nand2_2 _10174_ (.Y(_02394_),
    .A(_02386_),
    .B(_02391_));
 sg13g2_mux2_1 _10175_ (.A0(net1874),
    .A1(net3737),
    .S(_02394_),
    .X(_00069_));
 sg13g2_mux2_1 _10176_ (.A0(net1873),
    .A1(net3909),
    .S(_02394_),
    .X(_00070_));
 sg13g2_mux2_1 _10177_ (.A0(net1868),
    .A1(net3816),
    .S(_02394_),
    .X(_00071_));
 sg13g2_mux2_1 _10178_ (.A0(net1853),
    .A1(net3885),
    .S(_02394_),
    .X(_00072_));
 sg13g2_or4_1 _10179_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .B(net2502),
    .C(net2501),
    .D(_02390_),
    .X(_02395_));
 sg13g2_mux2_1 _10180_ (.A0(net1874),
    .A1(net3894),
    .S(_02395_),
    .X(_00065_));
 sg13g2_mux2_1 _10181_ (.A0(net1873),
    .A1(net3757),
    .S(_02395_),
    .X(_00066_));
 sg13g2_mux2_1 _10182_ (.A0(net1868),
    .A1(net3915),
    .S(_02395_),
    .X(_00067_));
 sg13g2_mux2_1 _10183_ (.A0(net1854),
    .A1(net4040),
    .S(_02395_),
    .X(_00068_));
 sg13g2_nand3b_1 _10184_ (.B(net1892),
    .C(_02096_),
    .Y(_02396_),
    .A_N(net2500));
 sg13g2_mux2_1 _10185_ (.A0(net1874),
    .A1(net3726),
    .S(_02396_),
    .X(_00061_));
 sg13g2_mux2_1 _10186_ (.A0(net1873),
    .A1(net3818),
    .S(_02396_),
    .X(_00062_));
 sg13g2_mux2_1 _10187_ (.A0(net1868),
    .A1(net3817),
    .S(_02396_),
    .X(_00063_));
 sg13g2_mux2_1 _10188_ (.A0(net1853),
    .A1(net3881),
    .S(_02396_),
    .X(_00064_));
 sg13g2_nor2b_1 _10189_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .B_N(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .Y(_02397_));
 sg13g2_nand3_1 _10190_ (.B(_02384_),
    .C(_02397_),
    .A(net1892),
    .Y(_02398_));
 sg13g2_mux2_1 _10191_ (.A0(net1875),
    .A1(net3622),
    .S(_02398_),
    .X(_00057_));
 sg13g2_mux2_1 _10192_ (.A0(net1872),
    .A1(net3567),
    .S(_02398_),
    .X(_00058_));
 sg13g2_mux2_1 _10193_ (.A0(net1868),
    .A1(net3570),
    .S(_02398_),
    .X(_00059_));
 sg13g2_mux2_1 _10194_ (.A0(net1853),
    .A1(net3779),
    .S(_02398_),
    .X(_00060_));
 sg13g2_nand3_1 _10195_ (.B(_02386_),
    .C(_02397_),
    .A(net1891),
    .Y(_02399_));
 sg13g2_mux2_1 _10196_ (.A0(net1875),
    .A1(net4006),
    .S(_02399_),
    .X(_00053_));
 sg13g2_mux2_1 _10197_ (.A0(net1872),
    .A1(net3678),
    .S(_02399_),
    .X(_00054_));
 sg13g2_mux2_1 _10198_ (.A0(net1867),
    .A1(net3969),
    .S(_02399_),
    .X(_00055_));
 sg13g2_mux2_1 _10199_ (.A0(net1854),
    .A1(net3829),
    .S(_02399_),
    .X(_00056_));
 sg13g2_nor2_1 _10200_ (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .B(net4166),
    .Y(_02400_));
 sg13g2_nand3_1 _10201_ (.B(_02384_),
    .C(_02400_),
    .A(net1891),
    .Y(_02401_));
 sg13g2_mux2_1 _10202_ (.A0(net1875),
    .A1(net3962),
    .S(_02401_),
    .X(_00049_));
 sg13g2_mux2_1 _10203_ (.A0(net1872),
    .A1(net4059),
    .S(_02401_),
    .X(_00050_));
 sg13g2_mux2_1 _10204_ (.A0(net1867),
    .A1(net4027),
    .S(_02401_),
    .X(_00051_));
 sg13g2_mux2_1 _10205_ (.A0(net1854),
    .A1(net4010),
    .S(_02401_),
    .X(_00052_));
 sg13g2_nand3_1 _10206_ (.B(_02386_),
    .C(net4167),
    .A(net1891),
    .Y(_02402_));
 sg13g2_mux2_1 _10207_ (.A0(net1875),
    .A1(net3838),
    .S(_02402_),
    .X(_00045_));
 sg13g2_mux2_1 _10208_ (.A0(net1872),
    .A1(net3640),
    .S(_02402_),
    .X(_00046_));
 sg13g2_mux2_1 _10209_ (.A0(net1867),
    .A1(net3854),
    .S(_02402_),
    .X(_00047_));
 sg13g2_mux2_1 _10210_ (.A0(net1854),
    .A1(net3806),
    .S(_02402_),
    .X(_00048_));
 sg13g2_and3_1 _10211_ (.X(_02403_),
    .A(_01025_),
    .B(_01027_),
    .C(\i_peripherals.func_sel[1] ));
 sg13g2_and4_1 _10212_ (.A(_01026_),
    .B(_01028_),
    .C(_01029_),
    .D(_02403_),
    .X(_02404_));
 sg13g2_nor2_1 _10213_ (.A(\i_peripherals.gpio_out[0] ),
    .B(_02404_),
    .Y(_02405_));
 sg13g2_nor3_1 _10214_ (.A(_01026_),
    .B(_01028_),
    .C(_01029_),
    .Y(_02406_));
 sg13g2_a221oi_1 _10215_ (.B2(_02403_),
    .C1(_02405_),
    .B1(_02406_),
    .A1(_01149_),
    .Y(uo_out[0]),
    .A2(_02404_));
 sg13g2_nand3_1 _10216_ (.B(_00993_),
    .C(\i_peripherals.func_sel[7] ),
    .A(_00991_),
    .Y(_02407_));
 sg13g2_nor4_1 _10217_ (.A(\i_peripherals.func_sel[10] ),
    .B(\i_peripherals.func_sel[8] ),
    .C(\i_peripherals.func_sel[6] ),
    .D(_02407_),
    .Y(_02408_));
 sg13g2_nor2_1 _10218_ (.A(\i_peripherals.gpio_out[1] ),
    .B(_02408_),
    .Y(_02409_));
 sg13g2_nor2b_1 _10219_ (.A(\i_peripherals.i_uart.i_uart_rx.uart_rts ),
    .B_N(_02408_),
    .Y(_02410_));
 sg13g2_nor4_1 _10220_ (.A(_00992_),
    .B(_00994_),
    .C(_00995_),
    .D(_02407_),
    .Y(_02411_));
 sg13g2_nor3_1 _10221_ (.A(_02409_),
    .B(_02410_),
    .C(_02411_),
    .Y(uo_out[1]));
 sg13g2_nor2b_1 _10222_ (.A(net2426),
    .B_N(net2427),
    .Y(_02412_));
 sg13g2_nand2b_2 _10223_ (.Y(_02413_),
    .B(net2427),
    .A_N(net2426));
 sg13g2_nor3_1 _10224_ (.A(net2424),
    .B(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .C(_02413_),
    .Y(_02414_));
 sg13g2_nand2_1 _10225_ (.Y(_02415_),
    .A(net2350),
    .B(_02414_));
 sg13g2_and2_1 _10226_ (.A(net2424),
    .B(_02412_),
    .X(_02416_));
 sg13g2_nor2b_2 _10227_ (.A(net2425),
    .B_N(net2426),
    .Y(_02417_));
 sg13g2_nor2b_1 _10228_ (.A(net2428),
    .B_N(_02417_),
    .Y(_02418_));
 sg13g2_nand2b_1 _10229_ (.Y(_02419_),
    .B(_02417_),
    .A_N(net2427));
 sg13g2_nand2_1 _10230_ (.Y(_02420_),
    .A(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .B(_02418_));
 sg13g2_o21ai_1 _10231_ (.B1(_02416_),
    .Y(_02421_),
    .A1(net2350),
    .A2(net2421));
 sg13g2_nand3_1 _10232_ (.B(_02420_),
    .C(_02421_),
    .A(_02415_),
    .Y(uio_out[1]));
 sg13g2_o21ai_1 _10233_ (.B1(_02413_),
    .Y(_02422_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .A2(_02419_));
 sg13g2_o21ai_1 _10234_ (.B1(_02416_),
    .Y(_02423_),
    .A1(net2350),
    .A2(\i_tinyqv.cpu.instr_data_in[13] ));
 sg13g2_nand3b_1 _10235_ (.B(_02422_),
    .C(_02423_),
    .Y(uio_out[2]),
    .A_N(_02414_));
 sg13g2_nand2_1 _10236_ (.Y(_02424_),
    .A(net2436),
    .B(_01129_));
 sg13g2_a22oi_1 _10237_ (.Y(_02425_),
    .B1(_02424_),
    .B2(_02416_),
    .A2(_02418_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[22] ));
 sg13g2_inv_2 _10238_ (.Y(uio_out[4]),
    .A(_02425_));
 sg13g2_o21ai_1 _10239_ (.B1(_02413_),
    .Y(_02426_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .A2(_02419_));
 sg13g2_o21ai_1 _10240_ (.B1(_02416_),
    .Y(_02427_),
    .A1(net2350),
    .A2(\i_tinyqv.cpu.instr_data_in[15] ));
 sg13g2_nand3_1 _10241_ (.B(_02426_),
    .C(_02427_),
    .A(_02415_),
    .Y(uio_out[5]));
 sg13g2_nand2b_1 _10242_ (.Y(_02428_),
    .B(net2271),
    .A_N(net4119));
 sg13g2_nor2_2 _10243_ (.A(net2302),
    .B(_01907_),
    .Y(_02429_));
 sg13g2_nand2_2 _10244_ (.Y(_02430_),
    .A(net2300),
    .B(_01908_));
 sg13g2_nand2_2 _10245_ (.Y(_02431_),
    .A(_02073_),
    .B(_02429_));
 sg13g2_mux2_1 _10246_ (.A0(net2396),
    .A1(_02428_),
    .S(_02431_),
    .X(_00002_));
 sg13g2_nand2b_1 _10247_ (.Y(_02432_),
    .B(net2271),
    .A_N(\time_limit[3] ));
 sg13g2_mux2_1 _10248_ (.A0(net2394),
    .A1(_02432_),
    .S(_02431_),
    .X(_00003_));
 sg13g2_nand2b_1 _10249_ (.Y(_02433_),
    .B(net2271),
    .A_N(net4122));
 sg13g2_mux2_1 _10250_ (.A0(net2392),
    .A1(_02433_),
    .S(_02431_),
    .X(_00004_));
 sg13g2_nand2_1 _10251_ (.Y(_02434_),
    .A(net2271),
    .B(_01109_));
 sg13g2_mux2_1 _10252_ (.A0(net2390),
    .A1(_02434_),
    .S(_02431_),
    .X(_00005_));
 sg13g2_a22oi_1 _10253_ (.Y(_02435_),
    .B1(_02073_),
    .B2(_02429_),
    .A2(net3782),
    .A1(net2270));
 sg13g2_nor2_2 _10254_ (.A(\data_to_write[6] ),
    .B(_02430_),
    .Y(_02436_));
 sg13g2_a21oi_1 _10255_ (.A1(_02073_),
    .A2(_02436_),
    .Y(_00006_),
    .B1(_02435_));
 sg13g2_nand2_1 _10256_ (.Y(_02437_),
    .A(_02276_),
    .B(_02429_));
 sg13g2_a22oi_1 _10257_ (.Y(_02438_),
    .B1(_02276_),
    .B2(_02429_),
    .A2(net3879),
    .A1(net2270));
 sg13g2_a21oi_1 _10258_ (.A1(_02276_),
    .A2(_02436_),
    .Y(_00000_),
    .B1(_02438_));
 sg13g2_nand2_1 _10259_ (.Y(_02439_),
    .A(net2270),
    .B(net4130));
 sg13g2_o21ai_1 _10260_ (.B1(_02439_),
    .Y(_02440_),
    .A1(net2270),
    .A2(net2));
 sg13g2_mux2_1 _10261_ (.A0(\data_to_write[7] ),
    .A1(_02440_),
    .S(_02437_),
    .X(_00001_));
 sg13g2_and2_1 _10262_ (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .B(net1),
    .X(uio_oe[5]));
 sg13g2_nand3_1 _10263_ (.B(_00998_),
    .C(\i_peripherals.func_sel[13] ),
    .A(_00996_),
    .Y(_02441_));
 sg13g2_nand3_1 _10264_ (.B(\i_peripherals.func_sel[14] ),
    .C(\i_peripherals.func_sel[12] ),
    .A(\i_peripherals.func_sel[16] ),
    .Y(_02442_));
 sg13g2_nor4_1 _10265_ (.A(\i_peripherals.func_sel[16] ),
    .B(\i_peripherals.func_sel[14] ),
    .C(\i_peripherals.func_sel[12] ),
    .D(_02441_),
    .Y(_02443_));
 sg13g2_or2_1 _10266_ (.X(_02444_),
    .B(_02443_),
    .A(\i_peripherals.gpio_out[2] ));
 sg13g2_o21ai_1 _10267_ (.B1(_02444_),
    .Y(_02445_),
    .A1(_02441_),
    .A2(_02442_));
 sg13g2_a21oi_1 _10268_ (.A1(_01149_),
    .A2(_02443_),
    .Y(_02446_),
    .B1(_02445_));
 sg13g2_mux2_1 _10269_ (.A0(_02446_),
    .A1(\debug_rd_r[0] ),
    .S(debug_register_data),
    .X(uo_out[2]));
 sg13g2_nand3_1 _10270_ (.B(_01003_),
    .C(\i_peripherals.func_sel[19] ),
    .A(_01001_),
    .Y(_02447_));
 sg13g2_nor4_1 _10271_ (.A(\i_peripherals.func_sel[22] ),
    .B(\i_peripherals.func_sel[20] ),
    .C(\i_peripherals.func_sel[18] ),
    .D(_02447_),
    .Y(_02448_));
 sg13g2_nor2_1 _10272_ (.A(\i_peripherals.gpio_out[3] ),
    .B(_02448_),
    .Y(_02449_));
 sg13g2_nor2b_1 _10273_ (.A(\i_peripherals.i_uart.i_uart_rx.uart_rts ),
    .B_N(_02448_),
    .Y(_02450_));
 sg13g2_nand3_1 _10274_ (.B(\i_peripherals.func_sel[20] ),
    .C(\i_peripherals.func_sel[18] ),
    .A(\i_peripherals.func_sel[22] ),
    .Y(_02451_));
 sg13g2_nor2_1 _10275_ (.A(_02447_),
    .B(_02451_),
    .Y(_02452_));
 sg13g2_nor3_1 _10276_ (.A(_02449_),
    .B(_02450_),
    .C(_02452_),
    .Y(_02453_));
 sg13g2_mux2_1 _10277_ (.A0(_02453_),
    .A1(\debug_rd_r[1] ),
    .S(debug_register_data),
    .X(uo_out[3]));
 sg13g2_nand3_1 _10278_ (.B(_01008_),
    .C(\i_peripherals.func_sel[25] ),
    .A(_01006_),
    .Y(_02454_));
 sg13g2_nor4_1 _10279_ (.A(\i_peripherals.func_sel[28] ),
    .B(\i_peripherals.func_sel[26] ),
    .C(\i_peripherals.func_sel[24] ),
    .D(_02454_),
    .Y(_02455_));
 sg13g2_or2_1 _10280_ (.X(_02456_),
    .B(_02455_),
    .A(\i_peripherals.gpio_out[4] ));
 sg13g2_nand3_1 _10281_ (.B(\i_peripherals.func_sel[26] ),
    .C(\i_peripherals.func_sel[24] ),
    .A(\i_peripherals.func_sel[28] ),
    .Y(_02457_));
 sg13g2_o21ai_1 _10282_ (.B1(_02456_),
    .Y(_02458_),
    .A1(_02454_),
    .A2(_02457_));
 sg13g2_a21oi_1 _10283_ (.A1(_01149_),
    .A2(_02455_),
    .Y(_02459_),
    .B1(_02458_));
 sg13g2_mux2_1 _10284_ (.A0(_02459_),
    .A1(\debug_rd_r[2] ),
    .S(debug_register_data),
    .X(uo_out[4]));
 sg13g2_nand3_1 _10285_ (.B(_01013_),
    .C(\i_peripherals.func_sel[31] ),
    .A(_01011_),
    .Y(_02460_));
 sg13g2_nand3_1 _10286_ (.B(\i_peripherals.func_sel[32] ),
    .C(\i_peripherals.func_sel[30] ),
    .A(\i_peripherals.func_sel[34] ),
    .Y(_02461_));
 sg13g2_nor4_1 _10287_ (.A(\i_peripherals.func_sel[34] ),
    .B(\i_peripherals.func_sel[32] ),
    .C(\i_peripherals.func_sel[30] ),
    .D(_02460_),
    .Y(_02462_));
 sg13g2_nor2_1 _10288_ (.A(\i_peripherals.gpio_out[5] ),
    .B(_02462_),
    .Y(_02463_));
 sg13g2_nor2b_1 _10289_ (.A(\i_peripherals.i_uart.i_uart_rx.uart_rts ),
    .B_N(_02462_),
    .Y(_02464_));
 sg13g2_nor2_1 _10290_ (.A(_02460_),
    .B(_02461_),
    .Y(_02465_));
 sg13g2_nor3_1 _10291_ (.A(_02463_),
    .B(_02464_),
    .C(_02465_),
    .Y(_02466_));
 sg13g2_mux2_1 _10292_ (.A0(_02466_),
    .A1(\debug_rd_r[3] ),
    .S(debug_register_data),
    .X(uo_out[5]));
 sg13g2_nor2b_1 _10293_ (.A(\gpio_out_sel[6] ),
    .B_N(debug_uart_txd),
    .Y(_02467_));
 sg13g2_or3_1 _10294_ (.A(\i_peripherals.func_sel[41] ),
    .B(\i_peripherals.func_sel[39] ),
    .C(_01018_),
    .X(_02468_));
 sg13g2_nor4_1 _10295_ (.A(\i_peripherals.func_sel[40] ),
    .B(\i_peripherals.func_sel[38] ),
    .C(\i_peripherals.func_sel[36] ),
    .D(_02468_),
    .Y(_02469_));
 sg13g2_nand3_1 _10296_ (.B(\i_peripherals.func_sel[38] ),
    .C(\i_peripherals.func_sel[36] ),
    .A(\i_peripherals.func_sel[40] ),
    .Y(_02470_));
 sg13g2_or2_1 _10297_ (.X(_02471_),
    .B(_02470_),
    .A(_02468_));
 sg13g2_o21ai_1 _10298_ (.B1(\gpio_out_sel[6] ),
    .Y(_02472_),
    .A1(\i_peripherals.gpio_out[6] ),
    .A2(_02469_));
 sg13g2_a21oi_1 _10299_ (.A1(_01149_),
    .A2(_02469_),
    .Y(_02473_),
    .B1(_02472_));
 sg13g2_a21o_2 _10300_ (.A2(_02473_),
    .A1(_02471_),
    .B1(_02467_),
    .X(uo_out[6]));
 sg13g2_nor3_2 _10301_ (.A(net2857),
    .B(net3839),
    .C(net4012),
    .Y(_02474_));
 sg13g2_and2_1 _10302_ (.A(_01433_),
    .B(_02474_),
    .X(_02475_));
 sg13g2_nand2_2 _10303_ (.Y(_02476_),
    .A(_01433_),
    .B(_02474_));
 sg13g2_o21ai_1 _10304_ (.B1(_02476_),
    .Y(_02477_),
    .A1(net2357),
    .A2(net2229));
 sg13g2_inv_1 _10305_ (.Y(_02478_),
    .A(_02477_));
 sg13g2_nor3_1 _10306_ (.A(_01417_),
    .B(_01432_),
    .C(_02474_),
    .Y(_02479_));
 sg13g2_nand2b_2 _10307_ (.Y(_02480_),
    .B(_01433_),
    .A_N(_02474_));
 sg13g2_a21oi_1 _10308_ (.A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(\i_tinyqv.cpu.i_core.cmp_out ),
    .Y(_02481_),
    .B1(net2306));
 sg13g2_o21ai_1 _10309_ (.B1(_02481_),
    .Y(_02482_),
    .A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(\i_tinyqv.cpu.i_core.cmp_out ));
 sg13g2_nor4_1 _10310_ (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .C(_01419_),
    .D(_01888_),
    .Y(_02483_));
 sg13g2_or2_1 _10311_ (.X(_02484_),
    .B(_02483_),
    .A(\i_tinyqv.cpu.i_core.is_interrupt ));
 sg13g2_nor3_2 _10312_ (.A(_01419_),
    .B(_01888_),
    .C(_01996_),
    .Y(_02485_));
 sg13g2_nand4_1 _10313_ (.B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .C(_01418_),
    .A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .Y(_02486_),
    .D(_01887_));
 sg13g2_nor3_1 _10314_ (.A(_01423_),
    .B(net2146),
    .C(_02485_),
    .Y(_02487_));
 sg13g2_a21oi_2 _10315_ (.B1(net2228),
    .Y(_02488_),
    .A2(_02487_),
    .A1(_02482_));
 sg13g2_a21o_2 _10316_ (.A2(_02487_),
    .A1(_02482_),
    .B1(net2228),
    .X(_02489_));
 sg13g2_nor2_1 _10317_ (.A(net2357),
    .B(\i_tinyqv.cpu.pc[2] ),
    .Y(_02490_));
 sg13g2_a21o_2 _10318_ (.A2(_02241_),
    .A1(net2357),
    .B1(_02490_),
    .X(_02491_));
 sg13g2_a21oi_1 _10319_ (.A1(net2357),
    .A2(_02241_),
    .Y(_02492_),
    .B1(_02490_));
 sg13g2_nor2_1 _10320_ (.A(net2357),
    .B(\i_tinyqv.cpu.pc[1] ),
    .Y(_02493_));
 sg13g2_a21o_2 _10321_ (.A2(_02167_),
    .A1(net2357),
    .B1(_02493_),
    .X(_02494_));
 sg13g2_a21oi_1 _10322_ (.A1(net2358),
    .A2(_02167_),
    .Y(_02495_),
    .B1(_02493_));
 sg13g2_mux4_1 _10323_ (.S0(net2218),
    .A0(\i_tinyqv.cpu.instr_data[1][0] ),
    .A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .A2(\i_tinyqv.cpu.instr_data[3][0] ),
    .A3(\i_tinyqv.cpu.instr_data[2][0] ),
    .S1(net2180),
    .X(_02496_));
 sg13g2_mux4_1 _10324_ (.S0(_02494_),
    .A0(\i_tinyqv.cpu.instr_data[1][1] ),
    .A1(\i_tinyqv.cpu.instr_data[0][1] ),
    .A2(\i_tinyqv.cpu.instr_data[3][1] ),
    .A3(\i_tinyqv.cpu.instr_data[2][1] ),
    .S1(net2181),
    .X(_02497_));
 sg13g2_inv_4 _10325_ (.A(net2143),
    .Y(_02498_));
 sg13g2_and2_1 _10326_ (.A(_02496_),
    .B(net2144),
    .X(_02499_));
 sg13g2_nand2_2 _10327_ (.Y(_02500_),
    .A(_02496_),
    .B(_02497_));
 sg13g2_nand2_1 _10328_ (.Y(_02501_),
    .A(_01076_),
    .B(net2185));
 sg13g2_nor2_1 _10329_ (.A(_01077_),
    .B(net2216),
    .Y(_02502_));
 sg13g2_nor2_1 _10330_ (.A(_01076_),
    .B(net2185),
    .Y(_02503_));
 sg13g2_xnor2_1 _10331_ (.Y(_02504_),
    .A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_02491_));
 sg13g2_o21ai_1 _10332_ (.B1(net2066),
    .Y(_02505_),
    .A1(_02502_),
    .A2(_02504_));
 sg13g2_nand2_1 _10333_ (.Y(_02506_),
    .A(net2358),
    .B(_01964_));
 sg13g2_xnor2_1 _10334_ (.Y(_02507_),
    .A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .B(_02506_));
 sg13g2_nand2_1 _10335_ (.Y(_02508_),
    .A(_01077_),
    .B(net2216));
 sg13g2_nor3_1 _10336_ (.A(_02503_),
    .B(_02507_),
    .C(_02508_),
    .Y(_02509_));
 sg13g2_a221oi_1 _10337_ (.B2(_02504_),
    .C1(_02509_),
    .B1(_02508_),
    .A1(_02501_),
    .Y(_02510_),
    .A2(_02507_));
 sg13g2_a21oi_1 _10338_ (.A1(_02505_),
    .A2(_02510_),
    .Y(_02511_),
    .B1(net2406));
 sg13g2_nand2_1 _10339_ (.Y(_02512_),
    .A(net1855),
    .B(_02511_));
 sg13g2_nand2_1 _10340_ (.Y(_02513_),
    .A(\i_tinyqv.cpu.i_core.mie[3] ),
    .B(_02363_));
 sg13g2_nand2_1 _10341_ (.Y(_02514_),
    .A(net3122),
    .B(\i_tinyqv.cpu.i_core.mie[1] ));
 sg13g2_a22oi_1 _10342_ (.Y(_02515_),
    .B1(\i_tinyqv.cpu.i_core.mie[1] ),
    .B2(net3122),
    .A2(net3310),
    .A1(net3409));
 sg13g2_and2_1 _10343_ (.A(\i_tinyqv.cpu.i_core.mie[16] ),
    .B(\i_tinyqv.cpu.i_core.mip[16] ),
    .X(_02516_));
 sg13g2_nand2_1 _10344_ (.Y(_02517_),
    .A(\i_tinyqv.cpu.i_core.mie[16] ),
    .B(\i_tinyqv.cpu.i_core.mip[16] ));
 sg13g2_nand2_1 _10345_ (.Y(_02518_),
    .A(\i_tinyqv.cpu.i_core.mie[2] ),
    .B(\i_peripherals.i_uart.uart_rx_buffered ));
 sg13g2_nand4_1 _10346_ (.B(_02515_),
    .C(_02517_),
    .A(_02513_),
    .Y(_02519_),
    .D(_02518_));
 sg13g2_nand2_2 _10347_ (.Y(_02520_),
    .A(net3903),
    .B(_02519_));
 sg13g2_o21ai_1 _10348_ (.B1(net2490),
    .Y(_02521_),
    .A1(_01432_),
    .A2(_02520_));
 sg13g2_nor4_2 _10349_ (.A(_02478_),
    .B(net1852),
    .C(_02512_),
    .Y(_02522_),
    .D(_02521_));
 sg13g2_mux4_1 _10350_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][13] ),
    .A1(\i_tinyqv.cpu.instr_data[0][13] ),
    .A2(\i_tinyqv.cpu.instr_data[3][13] ),
    .A3(\i_tinyqv.cpu.instr_data[2][13] ),
    .S1(net2183),
    .X(_02523_));
 sg13g2_mux4_1 _10351_ (.S0(net2218),
    .A0(\i_tinyqv.cpu.instr_data[1][14] ),
    .A1(\i_tinyqv.cpu.instr_data[0][14] ),
    .A2(\i_tinyqv.cpu.instr_data[3][14] ),
    .A3(\i_tinyqv.cpu.instr_data[2][14] ),
    .S1(net2185),
    .X(_02524_));
 sg13g2_inv_4 _10352_ (.A(net2139),
    .Y(_02525_));
 sg13g2_nor2_2 _10353_ (.A(net2141),
    .B(net2139),
    .Y(_02526_));
 sg13g2_or2_1 _10354_ (.X(_02527_),
    .B(net2139),
    .A(net2141));
 sg13g2_mux4_1 _10355_ (.S0(net2218),
    .A0(\i_tinyqv.cpu.instr_data[1][15] ),
    .A1(\i_tinyqv.cpu.instr_data[0][15] ),
    .A2(\i_tinyqv.cpu.instr_data[3][15] ),
    .A3(\i_tinyqv.cpu.instr_data[2][15] ),
    .S1(net2181),
    .X(_02528_));
 sg13g2_nand2b_2 _10356_ (.Y(_02529_),
    .B(_02528_),
    .A_N(_02496_));
 sg13g2_nor2_1 _10357_ (.A(_02498_),
    .B(_02529_),
    .Y(_02530_));
 sg13g2_nand2b_2 _10358_ (.Y(_02531_),
    .B(net2143),
    .A_N(_02529_));
 sg13g2_nor2_2 _10359_ (.A(_02527_),
    .B(_02531_),
    .Y(_02532_));
 sg13g2_nand2_1 _10360_ (.Y(_02533_),
    .A(_02526_),
    .B(_02530_));
 sg13g2_mux4_1 _10361_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][4] ),
    .A1(\i_tinyqv.cpu.instr_data[0][4] ),
    .A2(\i_tinyqv.cpu.instr_data[3][4] ),
    .A3(\i_tinyqv.cpu.instr_data[2][4] ),
    .S1(net2184),
    .X(_02534_));
 sg13g2_mux4_1 _10362_ (.S0(net2218),
    .A0(\i_tinyqv.cpu.instr_data[1][3] ),
    .A1(\i_tinyqv.cpu.instr_data[0][3] ),
    .A2(\i_tinyqv.cpu.instr_data[3][3] ),
    .A3(\i_tinyqv.cpu.instr_data[2][3] ),
    .S1(net2181),
    .X(_02535_));
 sg13g2_mux4_1 _10363_ (.S0(net2218),
    .A0(\i_tinyqv.cpu.instr_data[1][2] ),
    .A1(\i_tinyqv.cpu.instr_data[0][2] ),
    .A2(\i_tinyqv.cpu.instr_data[3][2] ),
    .A3(\i_tinyqv.cpu.instr_data[2][2] ),
    .S1(net2180),
    .X(_02536_));
 sg13g2_inv_2 _10364_ (.Y(_02537_),
    .A(_02536_));
 sg13g2_nor3_2 _10365_ (.A(net2138),
    .B(net2136),
    .C(_02536_),
    .Y(_02538_));
 sg13g2_inv_1 _10366_ (.Y(_02539_),
    .A(_02538_));
 sg13g2_mux4_1 _10367_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][5] ),
    .A1(\i_tinyqv.cpu.instr_data[0][5] ),
    .A2(\i_tinyqv.cpu.instr_data[3][5] ),
    .A3(\i_tinyqv.cpu.instr_data[2][5] ),
    .S1(net2183),
    .X(_02540_));
 sg13g2_mux4_1 _10368_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][6] ),
    .A1(\i_tinyqv.cpu.instr_data[0][6] ),
    .A2(\i_tinyqv.cpu.instr_data[3][6] ),
    .A3(\i_tinyqv.cpu.instr_data[2][6] ),
    .S1(net2182),
    .X(_02541_));
 sg13g2_nor2_1 _10369_ (.A(net2134),
    .B(net2131),
    .Y(_02542_));
 sg13g2_nor2_1 _10370_ (.A(_02539_),
    .B(net2131),
    .Y(_02543_));
 sg13g2_and2_1 _10371_ (.A(_02538_),
    .B(_02542_),
    .X(_02544_));
 sg13g2_and2_1 _10372_ (.A(_02532_),
    .B(_02544_),
    .X(_02545_));
 sg13g2_nand2_1 _10373_ (.Y(_02546_),
    .A(_02532_),
    .B(_02544_));
 sg13g2_mux4_1 _10374_ (.S0(_02494_),
    .A0(\i_tinyqv.cpu.instr_data[1][10] ),
    .A1(\i_tinyqv.cpu.instr_data[0][10] ),
    .A2(\i_tinyqv.cpu.instr_data[3][10] ),
    .A3(\i_tinyqv.cpu.instr_data[2][10] ),
    .S1(net2183),
    .X(_02547_));
 sg13g2_mux4_1 _10375_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][9] ),
    .A1(\i_tinyqv.cpu.instr_data[0][9] ),
    .A2(\i_tinyqv.cpu.instr_data[3][9] ),
    .A3(\i_tinyqv.cpu.instr_data[2][9] ),
    .S1(net2182),
    .X(_02548_));
 sg13g2_or2_1 _10376_ (.X(_02549_),
    .B(_02548_),
    .A(net2130));
 sg13g2_mux4_1 _10377_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][8] ),
    .A1(\i_tinyqv.cpu.instr_data[0][8] ),
    .A2(\i_tinyqv.cpu.instr_data[3][8] ),
    .A3(\i_tinyqv.cpu.instr_data[2][8] ),
    .S1(net2182),
    .X(_02550_));
 sg13g2_mux4_1 _10378_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][7] ),
    .A1(\i_tinyqv.cpu.instr_data[0][7] ),
    .A2(\i_tinyqv.cpu.instr_data[3][7] ),
    .A3(\i_tinyqv.cpu.instr_data[2][7] ),
    .S1(net2182),
    .X(_02551_));
 sg13g2_inv_1 _10379_ (.Y(_02552_),
    .A(_02551_));
 sg13g2_mux4_1 _10380_ (.S0(_02494_),
    .A0(\i_tinyqv.cpu.instr_data[1][12] ),
    .A1(\i_tinyqv.cpu.instr_data[0][12] ),
    .A2(\i_tinyqv.cpu.instr_data[3][12] ),
    .A3(\i_tinyqv.cpu.instr_data[2][12] ),
    .S1(net2181),
    .X(_02553_));
 sg13g2_nor4_1 _10381_ (.A(_02549_),
    .B(net2129),
    .C(_02552_),
    .D(net2126),
    .Y(_02554_));
 sg13g2_and2_1 _10382_ (.A(_02545_),
    .B(_02554_),
    .X(_02555_));
 sg13g2_and2_1 _10383_ (.A(_02522_),
    .B(_02555_),
    .X(_02556_));
 sg13g2_nand2_1 _10384_ (.Y(_02557_),
    .A(_02522_),
    .B(_02555_));
 sg13g2_nor2b_2 _10385_ (.A(net2139),
    .B_N(net2142),
    .Y(_02558_));
 sg13g2_nand2_2 _10386_ (.Y(_02559_),
    .A(net2142),
    .B(_02525_));
 sg13g2_nand2_2 _10387_ (.Y(_02560_),
    .A(_02496_),
    .B(_02498_));
 sg13g2_nor2_2 _10388_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 sg13g2_nand3_1 _10389_ (.B(_02498_),
    .C(_02558_),
    .A(_02496_),
    .Y(_02562_));
 sg13g2_nand2_2 _10390_ (.Y(_02563_),
    .A(net2134),
    .B(net2131));
 sg13g2_nor3_2 _10391_ (.A(net2138),
    .B(_02537_),
    .C(_02563_),
    .Y(_02564_));
 sg13g2_nand2_2 _10392_ (.Y(_02565_),
    .A(net2136),
    .B(_02564_));
 sg13g2_o21ai_1 _10393_ (.B1(_02562_),
    .Y(_02566_),
    .A1(net2064),
    .A2(_02565_));
 sg13g2_nand2_1 _10394_ (.Y(_02567_),
    .A(_02522_),
    .B(_02566_));
 sg13g2_nand2_1 _10395_ (.Y(_02568_),
    .A(net1809),
    .B(_02567_));
 sg13g2_nor2_1 _10396_ (.A(net2406),
    .B(net1855),
    .Y(_02569_));
 sg13g2_nor3_1 _10397_ (.A(net4139),
    .B(_02568_),
    .C(_02569_),
    .Y(_02570_));
 sg13g2_nand2_1 _10398_ (.Y(_02571_),
    .A(_01964_),
    .B(_02475_));
 sg13g2_nor2_1 _10399_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_00985_),
    .Y(_02572_));
 sg13g2_nor3_2 _10400_ (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_00985_),
    .C(net2335),
    .Y(_02573_));
 sg13g2_and2_1 _10401_ (.A(net2438),
    .B(_02573_),
    .X(_02574_));
 sg13g2_nand2_1 _10402_ (.Y(_02575_),
    .A(net4156),
    .B(_02574_));
 sg13g2_nand3_1 _10403_ (.B(net4152),
    .C(_02574_),
    .A(net4139),
    .Y(_02576_));
 sg13g2_or2_1 _10404_ (.X(_02577_),
    .B(_02576_),
    .A(_01076_));
 sg13g2_xnor2_1 _10405_ (.Y(_02578_),
    .A(net4158),
    .B(_02577_));
 sg13g2_xnor2_1 _10406_ (.Y(_02579_),
    .A(_02571_),
    .B(_02578_));
 sg13g2_xnor2_1 _10407_ (.Y(_02580_),
    .A(_01076_),
    .B(_02576_));
 sg13g2_xnor2_1 _10408_ (.Y(_02581_),
    .A(_01077_),
    .B(_02575_));
 sg13g2_xor2_1 _10409_ (.B(_02581_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .X(_02582_));
 sg13g2_xnor2_1 _10410_ (.Y(_02583_),
    .A(_00982_),
    .B(_02580_));
 sg13g2_nand3_1 _10411_ (.B(_02582_),
    .C(_02583_),
    .A(_02579_),
    .Y(_02584_));
 sg13g2_nand3_1 _10412_ (.B(net2335),
    .C(_02572_),
    .A(net2438),
    .Y(_02585_));
 sg13g2_or2_1 _10413_ (.X(_02586_),
    .B(_02585_),
    .A(_02584_));
 sg13g2_nand2_1 _10414_ (.Y(_02587_),
    .A(net4057),
    .B(_02586_));
 sg13g2_nor2b_1 _10415_ (.A(_02573_),
    .B_N(_02584_),
    .Y(_02588_));
 sg13g2_o21ai_1 _10416_ (.B1(net2302),
    .Y(_02589_),
    .A1(_01908_),
    .A2(_01914_));
 sg13g2_o21ai_1 _10417_ (.B1(net2438),
    .Y(_02590_),
    .A1(_02588_),
    .A2(_02589_));
 sg13g2_a21oi_1 _10418_ (.A1(_02570_),
    .A2(_02587_),
    .Y(_02591_),
    .B1(_02590_));
 sg13g2_nor2_2 _10419_ (.A(net2435),
    .B(net3423),
    .Y(_02592_));
 sg13g2_nor2_1 _10420_ (.A(net3646),
    .B(_02592_),
    .Y(_02593_));
 sg13g2_a21oi_1 _10421_ (.A1(_01437_),
    .A2(_02593_),
    .Y(_02594_),
    .B1(net4114));
 sg13g2_nor3_2 _10422_ (.A(_01913_),
    .B(_02591_),
    .C(_02594_),
    .Y(_02595_));
 sg13g2_inv_1 _10423_ (.Y(_02596_),
    .A(_02595_));
 sg13g2_a21oi_1 _10424_ (.A1(net2506),
    .A2(_02586_),
    .Y(_02597_),
    .B1(net6));
 sg13g2_o21ai_1 _10425_ (.B1(_02597_),
    .Y(_02598_),
    .A1(net5),
    .A2(_02595_));
 sg13g2_o21ai_1 _10426_ (.B1(net6),
    .Y(_02599_),
    .A1(net2506),
    .A2(debug_data_continue));
 sg13g2_a21oi_1 _10427_ (.A1(net2505),
    .A2(net2234),
    .Y(_02600_),
    .B1(_02599_));
 sg13g2_nor2_1 _10428_ (.A(net7),
    .B(_02600_),
    .Y(_02601_));
 sg13g2_a21oi_1 _10429_ (.A1(net2505),
    .A2(net1809),
    .Y(_02602_),
    .B1(net6));
 sg13g2_o21ai_1 _10430_ (.B1(_02602_),
    .Y(_02603_),
    .A1(net2505),
    .A2(net1892));
 sg13g2_a21oi_1 _10431_ (.A1(_02522_),
    .A2(_02566_),
    .Y(_02604_),
    .B1(net2505));
 sg13g2_a21oi_1 _10432_ (.A1(net2505),
    .A2(net1855),
    .Y(_02605_),
    .B1(_02604_));
 sg13g2_a21oi_1 _10433_ (.A1(net6),
    .A2(_02605_),
    .Y(_02606_),
    .B1(_01151_));
 sg13g2_a21oi_1 _10434_ (.A1(_00923_),
    .A2(net2505),
    .Y(_02607_),
    .B1(net6));
 sg13g2_o21ai_1 _10435_ (.B1(_02607_),
    .Y(_02608_),
    .A1(net2506),
    .A2(_02570_));
 sg13g2_a21oi_1 _10436_ (.A1(net2505),
    .A2(_02476_),
    .Y(_02609_),
    .B1(_01150_));
 sg13g2_o21ai_1 _10437_ (.B1(_02609_),
    .Y(_02610_),
    .A1(net2505),
    .A2(_02574_));
 sg13g2_nand3_1 _10438_ (.B(_02608_),
    .C(_02610_),
    .A(net7),
    .Y(_02611_));
 sg13g2_mux2_1 _10439_ (.A0(_02520_),
    .A1(_01943_),
    .S(net2506),
    .X(_02612_));
 sg13g2_nand2_2 _10440_ (.Y(_02613_),
    .A(net2300),
    .B(_01914_));
 sg13g2_a21oi_1 _10441_ (.A1(net2506),
    .A2(_02613_),
    .Y(_02614_),
    .B1(_01150_));
 sg13g2_o21ai_1 _10442_ (.B1(_02614_),
    .Y(_02615_),
    .A1(net2506),
    .A2(_02429_));
 sg13g2_o21ai_1 _10443_ (.B1(_02615_),
    .Y(_02616_),
    .A1(net6),
    .A2(_02612_));
 sg13g2_a22oi_1 _10444_ (.Y(_02617_),
    .B1(_02603_),
    .B2(_02606_),
    .A2(_02601_),
    .A1(_02598_));
 sg13g2_o21ai_1 _10445_ (.B1(_02611_),
    .Y(_02618_),
    .A1(net7),
    .A2(_02616_));
 sg13g2_a21oi_1 _10446_ (.A1(net8),
    .A2(_02618_),
    .Y(_02619_),
    .B1(\gpio_out_sel[7] ));
 sg13g2_o21ai_1 _10447_ (.B1(_02619_),
    .Y(_02620_),
    .A1(net8),
    .A2(_02617_));
 sg13g2_nor2_1 _10448_ (.A(\i_peripherals.func_sel[47] ),
    .B(\i_peripherals.func_sel[45] ),
    .Y(_02621_));
 sg13g2_nand2_1 _10449_ (.Y(_02622_),
    .A(\i_peripherals.func_sel[43] ),
    .B(_02621_));
 sg13g2_nor4_1 _10450_ (.A(\i_peripherals.func_sel[46] ),
    .B(\i_peripherals.func_sel[44] ),
    .C(\i_peripherals.func_sel[42] ),
    .D(_02622_),
    .Y(_02623_));
 sg13g2_nand2b_1 _10451_ (.Y(_02624_),
    .B(_02623_),
    .A_N(\i_peripherals.i_uart.i_uart_rx.uart_rts ));
 sg13g2_nand3_1 _10452_ (.B(\i_peripherals.func_sel[44] ),
    .C(\i_peripherals.func_sel[42] ),
    .A(\i_peripherals.func_sel[46] ),
    .Y(_02625_));
 sg13g2_o21ai_1 _10453_ (.B1(_02624_),
    .Y(_02626_),
    .A1(_02622_),
    .A2(_02625_));
 sg13g2_o21ai_1 _10454_ (.B1(\gpio_out_sel[7] ),
    .Y(_02627_),
    .A1(\i_peripherals.gpio_out[7] ),
    .A2(_02623_));
 sg13g2_o21ai_1 _10455_ (.B1(_02620_),
    .Y(uo_out[7]),
    .A1(_02626_),
    .A2(_02627_));
 sg13g2_mux2_1 _10456_ (.A0(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .A1(\i_tinyqv.mem.q_ctrl.spi_clk_neg ),
    .S(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ),
    .X(\i_tinyqv.mem.q_ctrl.spi_clk_out ));
 sg13g2_nand2_1 _10457_ (.Y(_02628_),
    .A(\i_tinyqv.cpu.is_load ),
    .B(_02476_));
 sg13g2_nor2_2 _10458_ (.A(net3576),
    .B(net2503),
    .Y(_02629_));
 sg13g2_nor4_1 _10459_ (.A(net3874),
    .B(net2504),
    .C(net2229),
    .D(_01416_),
    .Y(_02630_));
 sg13g2_and2_1 _10460_ (.A(_01403_),
    .B(_02630_),
    .X(_02631_));
 sg13g2_nand2_2 _10461_ (.Y(_02632_),
    .A(_01403_),
    .B(_02630_));
 sg13g2_nand3_1 _10462_ (.B(_02476_),
    .C(net2123),
    .A(\i_tinyqv.cpu.is_load ),
    .Y(_02633_));
 sg13g2_nor4_2 _10463_ (.A(net3576),
    .B(net2504),
    .C(net2229),
    .Y(_02634_),
    .D(_01406_));
 sg13g2_nand4_1 _10464_ (.B(net2232),
    .C(net2303),
    .A(net2357),
    .Y(_02635_),
    .D(_02629_));
 sg13g2_nand2_1 _10465_ (.Y(_02636_),
    .A(_02633_),
    .B(_02635_));
 sg13g2_o21ai_1 _10466_ (.B1(net2490),
    .Y(_02637_),
    .A1(net4002),
    .A2(_02634_));
 sg13g2_a22oi_1 _10467_ (.Y(_00019_),
    .B1(net4003),
    .B2(_02633_),
    .A2(_02636_),
    .A1(_02474_));
 sg13g2_nor2_1 _10468_ (.A(net1862),
    .B(net1812),
    .Y(_02638_));
 sg13g2_nand2_2 _10469_ (.Y(_02639_),
    .A(_02489_),
    .B(net1809));
 sg13g2_nand2_2 _10470_ (.Y(_02640_),
    .A(net2494),
    .B(_02638_));
 sg13g2_nor2b_1 _10471_ (.A(_02640_),
    .B_N(_02579_),
    .Y(_00077_));
 sg13g2_or2_1 _10472_ (.X(_02641_),
    .B(_02640_),
    .A(_02575_));
 sg13g2_nor3_1 _10473_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(_01077_),
    .C(_02641_),
    .Y(_02642_));
 sg13g2_mux2_1 _10474_ (.A0(net3404),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net1754),
    .X(_00078_));
 sg13g2_mux2_1 _10475_ (.A0(net3456),
    .A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .S(net1757),
    .X(_00079_));
 sg13g2_nor2_1 _10476_ (.A(net3207),
    .B(net1755),
    .Y(_02643_));
 sg13g2_a21oi_1 _10477_ (.A1(_01118_),
    .A2(net1755),
    .Y(_00080_),
    .B1(_02643_));
 sg13g2_mux2_1 _10478_ (.A0(net3346),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(net1756),
    .X(_00081_));
 sg13g2_mux2_1 _10479_ (.A0(net3410),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net1754),
    .X(_00082_));
 sg13g2_nor2_1 _10480_ (.A(net3127),
    .B(net1754),
    .Y(_02644_));
 sg13g2_a21oi_1 _10481_ (.A1(_01134_),
    .A2(net1754),
    .Y(_00083_),
    .B1(_02644_));
 sg13g2_mux2_1 _10482_ (.A0(net3527),
    .A1(net2422),
    .S(net1754),
    .X(_00084_));
 sg13g2_nor2_1 _10483_ (.A(net3120),
    .B(net1754),
    .Y(_02645_));
 sg13g2_a21oi_1 _10484_ (.A1(_01124_),
    .A2(net1754),
    .Y(_00085_),
    .B1(_02645_));
 sg13g2_nor2_1 _10485_ (.A(net3373),
    .B(net1755),
    .Y(_02646_));
 sg13g2_a21oi_1 _10486_ (.A1(_01128_),
    .A2(net1755),
    .Y(_00086_),
    .B1(_02646_));
 sg13g2_nor2_1 _10487_ (.A(net3142),
    .B(net1754),
    .Y(_02647_));
 sg13g2_a21oi_1 _10488_ (.A1(_01133_),
    .A2(net1756),
    .Y(_00087_),
    .B1(_02647_));
 sg13g2_mux2_1 _10489_ (.A0(net3623),
    .A1(net2420),
    .S(net1755),
    .X(_00088_));
 sg13g2_nor2_1 _10490_ (.A(net3089),
    .B(net1756),
    .Y(_02648_));
 sg13g2_a21oi_1 _10491_ (.A1(_01125_),
    .A2(net1756),
    .Y(_00089_),
    .B1(_02648_));
 sg13g2_nor2_1 _10492_ (.A(net3056),
    .B(net1757),
    .Y(_02649_));
 sg13g2_a21oi_1 _10493_ (.A1(_01129_),
    .A2(net1757),
    .Y(_00090_),
    .B1(net3057));
 sg13g2_mux2_1 _10494_ (.A0(net3383),
    .A1(net2419),
    .S(net1757),
    .X(_00091_));
 sg13g2_nor3_1 _10495_ (.A(net4067),
    .B(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .C(net2236),
    .Y(_02650_));
 sg13g2_o21ai_1 _10496_ (.B1(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .Y(_02651_),
    .A1(net4067),
    .A2(net2237));
 sg13g2_nand2_1 _10497_ (.Y(_02652_),
    .A(net2486),
    .B(_02651_));
 sg13g2_nor2_1 _10498_ (.A(net4068),
    .B(_02652_),
    .Y(_00092_));
 sg13g2_nor2_1 _10499_ (.A(_01116_),
    .B(_02651_),
    .Y(_02653_));
 sg13g2_a21oi_1 _10500_ (.A1(_01116_),
    .A2(_02651_),
    .Y(_02654_),
    .B1(net2339));
 sg13g2_nor2b_1 _10501_ (.A(_02653_),
    .B_N(net4046),
    .Y(_00093_));
 sg13g2_and2_1 _10502_ (.A(net3729),
    .B(_02653_),
    .X(_02655_));
 sg13g2_o21ai_1 _10503_ (.B1(net2486),
    .Y(_02656_),
    .A1(net3729),
    .A2(_02653_));
 sg13g2_nor2_1 _10504_ (.A(_02655_),
    .B(net3730),
    .Y(_00094_));
 sg13g2_and2_1 _10505_ (.A(net3943),
    .B(_02655_),
    .X(_02657_));
 sg13g2_o21ai_1 _10506_ (.B1(net2486),
    .Y(_02658_),
    .A1(net3943),
    .A2(_02655_));
 sg13g2_nor2_1 _10507_ (.A(_02657_),
    .B(net3944),
    .Y(_00095_));
 sg13g2_mux2_1 _10508_ (.A0(\i_tinyqv.cpu.i_core.i_instrret.add ),
    .A1(\i_tinyqv.cpu.i_core.i_instrret.cy ),
    .S(net2235),
    .X(_02659_));
 sg13g2_and2_1 _10509_ (.A(net3888),
    .B(_02659_),
    .X(_02660_));
 sg13g2_and2_1 _10510_ (.A(net3923),
    .B(_02660_),
    .X(_02661_));
 sg13g2_nand2_1 _10511_ (.Y(_02662_),
    .A(net3899),
    .B(_02661_));
 sg13g2_nor3_1 _10512_ (.A(net2348),
    .B(_01132_),
    .C(_02662_),
    .Y(_00096_));
 sg13g2_nand2_1 _10513_ (.Y(_02663_),
    .A(_01343_),
    .B(_02629_));
 sg13g2_mux2_1 _10514_ (.A0(_01360_),
    .A1(_01367_),
    .S(_01407_),
    .X(_02664_));
 sg13g2_mux2_1 _10515_ (.A0(_02664_),
    .A1(net3575),
    .S(_02663_),
    .X(_00097_));
 sg13g2_and2_1 _10516_ (.A(net2486),
    .B(_02657_),
    .X(_00098_));
 sg13g2_o21ai_1 _10517_ (.B1(net2492),
    .Y(_02665_),
    .A1(net3888),
    .A2(_02659_));
 sg13g2_nor2_1 _10518_ (.A(_02660_),
    .B(net3889),
    .Y(_00099_));
 sg13g2_o21ai_1 _10519_ (.B1(net2492),
    .Y(_02666_),
    .A1(net3923),
    .A2(_02660_));
 sg13g2_nor2_1 _10520_ (.A(_02661_),
    .B(_02666_),
    .Y(_00100_));
 sg13g2_o21ai_1 _10521_ (.B1(net2492),
    .Y(_02667_),
    .A1(net3899),
    .A2(_02661_));
 sg13g2_nor2b_1 _10522_ (.A(net3900),
    .B_N(_02662_),
    .Y(_00101_));
 sg13g2_xnor2_1 _10523_ (.Y(_02668_),
    .A(_01132_),
    .B(_02662_));
 sg13g2_nor2_1 _10524_ (.A(net2348),
    .B(_02668_),
    .Y(_00102_));
 sg13g2_nor3_1 _10525_ (.A(net2234),
    .B(_01957_),
    .C(_02629_),
    .Y(_02669_));
 sg13g2_a21o_1 _10526_ (.A2(net2233),
    .A1(net2968),
    .B1(_02669_),
    .X(_00103_));
 sg13g2_nand2_1 _10527_ (.Y(_02670_),
    .A(net2488),
    .B(_01432_));
 sg13g2_nor2_1 _10528_ (.A(net2228),
    .B(_01716_),
    .Y(_02671_));
 sg13g2_nor2_1 _10529_ (.A(net2504),
    .B(net2232),
    .Y(_02672_));
 sg13g2_nor3_1 _10530_ (.A(_02670_),
    .B(_02671_),
    .C(_02672_),
    .Y(_00104_));
 sg13g2_a21oi_1 _10531_ (.A1(net2504),
    .A2(net2232),
    .Y(_02673_),
    .B1(net3576));
 sg13g2_nor2_1 _10532_ (.A(_02670_),
    .B(net3577),
    .Y(_00105_));
 sg13g2_and2_1 _10533_ (.A(net2236),
    .B(_02483_),
    .X(_02674_));
 sg13g2_nand2_2 _10534_ (.Y(_02675_),
    .A(net2236),
    .B(_02483_));
 sg13g2_a21oi_1 _10535_ (.A1(net2999),
    .A2(_02674_),
    .Y(_02676_),
    .B1(net3038));
 sg13g2_a22oi_1 _10536_ (.Y(_02677_),
    .B1(_02674_),
    .B2(net2999),
    .A2(net2234),
    .A1(net3038));
 sg13g2_inv_1 _10537_ (.Y(_00106_),
    .A(_02677_));
 sg13g2_and2_1 _10538_ (.A(net2231),
    .B(_02657_),
    .X(_02678_));
 sg13g2_and2_1 _10539_ (.A(net3676),
    .B(_02678_),
    .X(_02679_));
 sg13g2_o21ai_1 _10540_ (.B1(net2486),
    .Y(_02680_),
    .A1(net3676),
    .A2(_02678_));
 sg13g2_nor2_1 _10541_ (.A(_02679_),
    .B(net3677),
    .Y(_00107_));
 sg13g2_or2_1 _10542_ (.X(_02681_),
    .B(_02679_),
    .A(net4079));
 sg13g2_nand2_1 _10543_ (.Y(_02682_),
    .A(net4079),
    .B(_02679_));
 sg13g2_and3_1 _10544_ (.X(_00108_),
    .A(net2486),
    .B(_02681_),
    .C(_02682_));
 sg13g2_o21ai_1 _10545_ (.B1(net2486),
    .Y(_02683_),
    .A1(_01066_),
    .A2(_02682_));
 sg13g2_a21oi_1 _10546_ (.A1(_01066_),
    .A2(_02682_),
    .Y(_00109_),
    .B1(_02683_));
 sg13g2_nand3_1 _10547_ (.B(_02363_),
    .C(_02518_),
    .A(\i_tinyqv.cpu.i_core.mie[3] ),
    .Y(_02684_));
 sg13g2_a22oi_1 _10548_ (.Y(_02685_),
    .B1(_02514_),
    .B2(_02684_),
    .A2(net3310),
    .A1(net3409));
 sg13g2_o21ai_1 _10549_ (.B1(net3476),
    .Y(_02686_),
    .A1(_02516_),
    .A2(_02685_));
 sg13g2_nor4_1 _10550_ (.A(net3476),
    .B(_01223_),
    .C(_01282_),
    .D(_01318_),
    .Y(_02687_));
 sg13g2_and2_1 _10551_ (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .B(net2236),
    .X(_02688_));
 sg13g2_nand2_2 _10552_ (.Y(_02689_),
    .A(net3476),
    .B(net2236));
 sg13g2_nand2_2 _10553_ (.Y(_02690_),
    .A(net2236),
    .B(net2146));
 sg13g2_nand2_2 _10554_ (.Y(_02691_),
    .A(_02675_),
    .B(_02689_));
 sg13g2_nor2_1 _10555_ (.A(_02687_),
    .B(_02690_),
    .Y(_02692_));
 sg13g2_o21ai_1 _10556_ (.B1(net2486),
    .Y(_02693_),
    .A1(net3780),
    .A2(_02691_));
 sg13g2_a21oi_1 _10557_ (.A1(_02686_),
    .A2(_02692_),
    .Y(_00110_),
    .B1(_02693_));
 sg13g2_nand2_1 _10558_ (.Y(_02694_),
    .A(_02513_),
    .B(_02518_));
 sg13g2_a221oi_1 _10559_ (.B2(_02694_),
    .C1(_02689_),
    .B1(_02515_),
    .A1(\i_tinyqv.cpu.i_core.mie[16] ),
    .Y(_02695_),
    .A2(\i_tinyqv.cpu.i_core.mip[16] ));
 sg13g2_o21ai_1 _10560_ (.B1(net2487),
    .Y(_02696_),
    .A1(net3468),
    .A2(_02691_));
 sg13g2_nor2_1 _10561_ (.A(_02695_),
    .B(_02696_),
    .Y(_00111_));
 sg13g2_a22oi_1 _10562_ (.Y(_02697_),
    .B1(_02690_),
    .B2(net2937),
    .A2(_02688_),
    .A1(_02516_));
 sg13g2_nor2_1 _10563_ (.A(net2339),
    .B(net2938),
    .Y(_00112_));
 sg13g2_nor2_1 _10564_ (.A(_01367_),
    .B(_02690_),
    .Y(_02698_));
 sg13g2_a22oi_1 _10565_ (.Y(_02699_),
    .B1(_02698_),
    .B2(_02687_),
    .A2(_02690_),
    .A1(net3185));
 sg13g2_nor2_1 _10566_ (.A(net2339),
    .B(net3186),
    .Y(_00113_));
 sg13g2_a22oi_1 _10567_ (.Y(_02700_),
    .B1(_02690_),
    .B2(net3189),
    .A2(_02688_),
    .A1(_02517_));
 sg13g2_nor2_1 _10568_ (.A(net2339),
    .B(net3190),
    .Y(_00114_));
 sg13g2_a21oi_1 _10569_ (.A1(net3060),
    .A2(_02675_),
    .Y(_02701_),
    .B1(_02688_));
 sg13g2_nor2_1 _10570_ (.A(net2339),
    .B(net3061),
    .Y(_00115_));
 sg13g2_a21oi_1 _10571_ (.A1(net2999),
    .A2(net2223),
    .Y(_02702_),
    .B1(_02691_));
 sg13g2_nor2b_1 _10572_ (.A(_02702_),
    .B_N(_02676_),
    .Y(_00116_));
 sg13g2_nand2_1 _10573_ (.Y(_02703_),
    .A(net2837),
    .B(_02002_));
 sg13g2_nand2_2 _10574_ (.Y(_02704_),
    .A(net2485),
    .B(net2295));
 sg13g2_nand2_1 _10575_ (.Y(_02705_),
    .A(net2374),
    .B(_01418_));
 sg13g2_nor2_2 _10576_ (.A(_01410_),
    .B(_01419_),
    .Y(_02706_));
 sg13g2_nor2b_2 _10577_ (.A(_02000_),
    .B_N(_02706_),
    .Y(_02707_));
 sg13g2_nand2b_1 _10578_ (.Y(_02708_),
    .B(_02707_),
    .A_N(_01341_));
 sg13g2_nor2_1 _10579_ (.A(\i_tinyqv.cpu.i_core.mepc[0] ),
    .B(_02707_),
    .Y(_02709_));
 sg13g2_nor2_1 _10580_ (.A(net2145),
    .B(_02709_),
    .Y(_02710_));
 sg13g2_a22oi_1 _10581_ (.Y(_02711_),
    .B1(_02708_),
    .B2(_02710_),
    .A2(net2145),
    .A1(_01348_));
 sg13g2_o21ai_1 _10582_ (.B1(_02703_),
    .Y(_00117_),
    .A1(_02704_),
    .A2(_02711_));
 sg13g2_nand2_1 _10583_ (.Y(_02712_),
    .A(net2861),
    .B(_02002_));
 sg13g2_nand2b_1 _10584_ (.Y(_02713_),
    .B(_02707_),
    .A_N(_01305_));
 sg13g2_nor2_1 _10585_ (.A(\i_tinyqv.cpu.i_core.mepc[1] ),
    .B(_02707_),
    .Y(_02714_));
 sg13g2_nor2_1 _10586_ (.A(net2145),
    .B(_02714_),
    .Y(_02715_));
 sg13g2_a22oi_1 _10587_ (.Y(_02716_),
    .B1(_02713_),
    .B2(_02715_),
    .A2(net2145),
    .A1(_01310_));
 sg13g2_o21ai_1 _10588_ (.B1(_02712_),
    .Y(_00118_),
    .A1(_02704_),
    .A2(_02716_));
 sg13g2_nand2_1 _10589_ (.Y(_02717_),
    .A(net2859),
    .B(_02002_));
 sg13g2_nand2_1 _10590_ (.Y(_02718_),
    .A(_01269_),
    .B(_02707_));
 sg13g2_nor2_1 _10591_ (.A(\i_tinyqv.cpu.i_core.mepc[2] ),
    .B(_02707_),
    .Y(_02719_));
 sg13g2_nor2_1 _10592_ (.A(net2145),
    .B(_02719_),
    .Y(_02720_));
 sg13g2_a22oi_1 _10593_ (.Y(_02721_),
    .B1(_02718_),
    .B2(_02720_),
    .A2(net2145),
    .A1(_01274_));
 sg13g2_o21ai_1 _10594_ (.B1(_02717_),
    .Y(_00119_),
    .A1(_02704_),
    .A2(_02721_));
 sg13g2_nand2_1 _10595_ (.Y(_02722_),
    .A(net2828),
    .B(_02002_));
 sg13g2_nand2_1 _10596_ (.Y(_02723_),
    .A(_01190_),
    .B(_02707_));
 sg13g2_nor2_1 _10597_ (.A(\i_tinyqv.cpu.i_core.mepc[3] ),
    .B(_02707_),
    .Y(_02724_));
 sg13g2_nor2_1 _10598_ (.A(net2146),
    .B(_02724_),
    .Y(_02725_));
 sg13g2_a22oi_1 _10599_ (.Y(_02726_),
    .B1(_02723_),
    .B2(_02725_),
    .A2(net2145),
    .A1(_01210_));
 sg13g2_o21ai_1 _10600_ (.B1(_02722_),
    .Y(_00120_),
    .A1(_02704_),
    .A2(_02726_));
 sg13g2_and2_1 _10601_ (.A(net2487),
    .B(_02676_),
    .X(_02727_));
 sg13g2_nand2_1 _10602_ (.Y(_02728_),
    .A(net2487),
    .B(_02676_));
 sg13g2_nand2_1 _10603_ (.Y(_02729_),
    .A(net2244),
    .B(net1994));
 sg13g2_mux2_1 _10604_ (.A0(\i_peripherals.i_uart.ui_in[0] ),
    .A1(net3129),
    .S(_02729_),
    .X(_00121_));
 sg13g2_mux2_1 _10605_ (.A0(\i_peripherals.i_uart.ui_in[1] ),
    .A1(net3140),
    .S(_02729_),
    .X(_00122_));
 sg13g2_nand2_1 _10606_ (.Y(_02730_),
    .A(_01343_),
    .B(net2223));
 sg13g2_o21ai_1 _10607_ (.B1(_02690_),
    .Y(_02731_),
    .A1(_02248_),
    .A2(_02730_));
 sg13g2_nor2_2 _10608_ (.A(_01189_),
    .B(_02706_),
    .Y(_02732_));
 sg13g2_nor3_1 _10609_ (.A(net2373),
    .B(_01190_),
    .C(_01990_),
    .Y(_02733_));
 sg13g2_nor2_1 _10610_ (.A(_02248_),
    .B(_02733_),
    .Y(_02734_));
 sg13g2_o21ai_1 _10611_ (.B1(_02734_),
    .Y(_02735_),
    .A1(_02705_),
    .A2(_02732_));
 sg13g2_o21ai_1 _10612_ (.B1(_02731_),
    .Y(_02736_),
    .A1(_02730_),
    .A2(_02735_));
 sg13g2_and2_1 _10613_ (.A(_01189_),
    .B(_02706_),
    .X(_02737_));
 sg13g2_o21ai_1 _10614_ (.B1(_02690_),
    .Y(_02738_),
    .A1(_02733_),
    .A2(_02737_));
 sg13g2_nand2b_1 _10615_ (.Y(_02739_),
    .B(_02738_),
    .A_N(_02736_));
 sg13g2_a21oi_1 _10616_ (.A1(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .A2(_02691_),
    .Y(_02740_),
    .B1(_02739_));
 sg13g2_nor2b_1 _10617_ (.A(net3097),
    .B_N(_02736_),
    .Y(_02741_));
 sg13g2_nor3_1 _10618_ (.A(net1993),
    .B(_02740_),
    .C(_02741_),
    .Y(_00123_));
 sg13g2_a221oi_1 _10619_ (.B2(_02250_),
    .C1(_02485_),
    .B1(_02735_),
    .A1(net2236),
    .Y(_02742_),
    .A2(net2146));
 sg13g2_nand3_1 _10620_ (.B(net2186),
    .C(_02690_),
    .A(net3097),
    .Y(_02743_));
 sg13g2_a21oi_1 _10621_ (.A1(_02738_),
    .A2(_02743_),
    .Y(_02744_),
    .B1(_02742_));
 sg13g2_a21oi_1 _10622_ (.A1(net3903),
    .A2(_02742_),
    .Y(_02745_),
    .B1(_02728_));
 sg13g2_nand2b_1 _10623_ (.Y(_00124_),
    .B(_02745_),
    .A_N(_02744_));
 sg13g2_nand2_1 _10624_ (.Y(_02746_),
    .A(net3713),
    .B(_02474_));
 sg13g2_nor3_1 _10625_ (.A(_01432_),
    .B(_02520_),
    .C(_02746_),
    .Y(_02747_));
 sg13g2_nor2b_1 _10626_ (.A(_02747_),
    .B_N(_02511_),
    .Y(_02748_));
 sg13g2_o21ai_1 _10627_ (.B1(_02748_),
    .Y(_02749_),
    .A1(_02477_),
    .A2(net1861));
 sg13g2_nand2_2 _10628_ (.Y(_02750_),
    .A(_02480_),
    .B(_02749_));
 sg13g2_nand2_2 _10629_ (.Y(_02751_),
    .A(net2498),
    .B(_02750_));
 sg13g2_nor2_2 _10630_ (.A(_02528_),
    .B(_02560_),
    .Y(_02752_));
 sg13g2_nor3_1 _10631_ (.A(net2142),
    .B(_02528_),
    .C(_02560_),
    .Y(_02753_));
 sg13g2_nor2_1 _10632_ (.A(_02496_),
    .B(_02528_),
    .Y(_02754_));
 sg13g2_and2_1 _10633_ (.A(net2143),
    .B(_02754_),
    .X(_02755_));
 sg13g2_nand2_1 _10634_ (.Y(_02756_),
    .A(net2143),
    .B(_02754_));
 sg13g2_and2_1 _10635_ (.A(_02526_),
    .B(_02754_),
    .X(_02757_));
 sg13g2_nor2_1 _10636_ (.A(_02527_),
    .B(_02756_),
    .Y(_02758_));
 sg13g2_nor2_2 _10637_ (.A(_02753_),
    .B(_02758_),
    .Y(_02759_));
 sg13g2_and2_1 _10638_ (.A(net2142),
    .B(net2140),
    .X(_02760_));
 sg13g2_inv_1 _10639_ (.Y(_02761_),
    .A(_02760_));
 sg13g2_nand2_2 _10640_ (.Y(_02762_),
    .A(_02752_),
    .B(_02760_));
 sg13g2_inv_1 _10641_ (.Y(_02763_),
    .A(_02762_));
 sg13g2_nor2_2 _10642_ (.A(_02531_),
    .B(_02559_),
    .Y(_02764_));
 sg13g2_nand2_1 _10643_ (.Y(_02765_),
    .A(_02530_),
    .B(_02558_));
 sg13g2_nand2_2 _10644_ (.Y(_02766_),
    .A(net2139),
    .B(_02755_));
 sg13g2_nand4_1 _10645_ (.B(_02762_),
    .C(_02765_),
    .A(_02759_),
    .Y(_02767_),
    .D(_02766_));
 sg13g2_nor2_1 _10646_ (.A(_02533_),
    .B(_02544_),
    .Y(_02768_));
 sg13g2_nor2_1 _10647_ (.A(_02767_),
    .B(_02768_),
    .Y(_02769_));
 sg13g2_nor2b_2 _10648_ (.A(_02560_),
    .B_N(_02528_),
    .Y(_02770_));
 sg13g2_and2_1 _10649_ (.A(_02526_),
    .B(_02770_),
    .X(_02771_));
 sg13g2_nand2_2 _10650_ (.Y(_02772_),
    .A(_02526_),
    .B(_02770_));
 sg13g2_nand3_1 _10651_ (.B(_02769_),
    .C(_02772_),
    .A(net2064),
    .Y(_02773_));
 sg13g2_nor2_2 _10652_ (.A(_02559_),
    .B(_02756_),
    .Y(_02774_));
 sg13g2_nand2_2 _10653_ (.Y(_02775_),
    .A(_02558_),
    .B(_02755_));
 sg13g2_a22oi_1 _10654_ (.Y(_02776_),
    .B1(_02558_),
    .B2(_02752_),
    .A2(net2128),
    .A1(_02545_));
 sg13g2_nand2_2 _10655_ (.Y(_02777_),
    .A(_02759_),
    .B(_02772_));
 sg13g2_and2_1 _10656_ (.A(_02527_),
    .B(_02754_),
    .X(_02778_));
 sg13g2_nand2_1 _10657_ (.Y(_02779_),
    .A(_02527_),
    .B(_02755_));
 sg13g2_nand3_1 _10658_ (.B(_02772_),
    .C(_02779_),
    .A(_02759_),
    .Y(_02780_));
 sg13g2_nor4_2 _10659_ (.A(_02532_),
    .B(_02561_),
    .C(_02767_),
    .Y(_02781_),
    .D(_02780_));
 sg13g2_nor2_1 _10660_ (.A(net2070),
    .B(_02537_),
    .Y(_02782_));
 sg13g2_a22oi_1 _10661_ (.Y(_02783_),
    .B1(_02781_),
    .B2(_02782_),
    .A2(_02773_),
    .A1(_02551_));
 sg13g2_and4_1 _10662_ (.A(_02480_),
    .B(_02775_),
    .C(_02776_),
    .D(_02783_),
    .X(_02784_));
 sg13g2_a21oi_1 _10663_ (.A1(net2502),
    .A2(net1850),
    .Y(_02785_),
    .B1(_02784_));
 sg13g2_mux2_1 _10664_ (.A0(_02785_),
    .A1(net2502),
    .S(_02751_),
    .X(_00125_));
 sg13g2_nor3_1 _10665_ (.A(_02384_),
    .B(_02386_),
    .C(_02480_),
    .Y(_02786_));
 sg13g2_nand2_1 _10666_ (.Y(_02787_),
    .A(net2064),
    .B(net2137));
 sg13g2_inv_1 _10667_ (.Y(_02788_),
    .A(_02787_));
 sg13g2_a221oi_1 _10668_ (.B2(_02788_),
    .C1(net1850),
    .B1(_02781_),
    .A1(net2129),
    .Y(_02789_),
    .A2(_02773_));
 sg13g2_nor3_1 _10669_ (.A(net1806),
    .B(_02786_),
    .C(_02789_),
    .Y(_02790_));
 sg13g2_a21o_1 _10670_ (.A2(net1805),
    .A1(net3917),
    .B1(_02790_),
    .X(_00126_));
 sg13g2_a21oi_1 _10671_ (.A1(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .A2(net4165),
    .Y(_02791_),
    .B1(net2501));
 sg13g2_or2_1 _10672_ (.X(_02792_),
    .B(_02791_),
    .A(_02096_));
 sg13g2_nand2_1 _10673_ (.Y(_02793_),
    .A(net2065),
    .B(net2138));
 sg13g2_inv_1 _10674_ (.Y(_02794_),
    .A(_02793_));
 sg13g2_a221oi_1 _10675_ (.B2(_02794_),
    .C1(net1850),
    .B1(_02781_),
    .A1(_02548_),
    .Y(_02795_),
    .A2(_02773_));
 sg13g2_a21oi_1 _10676_ (.A1(net1850),
    .A2(_02792_),
    .Y(_02796_),
    .B1(_02795_));
 sg13g2_mux2_1 _10677_ (.A0(_02796_),
    .A1(net2501),
    .S(net1805),
    .X(_00127_));
 sg13g2_xnor2_1 _10678_ (.Y(_02797_),
    .A(net2500),
    .B(_02096_));
 sg13g2_or2_1 _10679_ (.X(_02798_),
    .B(_02781_),
    .A(_02771_));
 sg13g2_nand3_1 _10680_ (.B(_02769_),
    .C(_02775_),
    .A(net2064),
    .Y(_02799_));
 sg13g2_a221oi_1 _10681_ (.B2(_02547_),
    .C1(net1850),
    .B1(_02799_),
    .A1(net2064),
    .Y(_02800_),
    .A2(_02798_));
 sg13g2_a21oi_1 _10682_ (.A1(net1850),
    .A2(_02797_),
    .Y(_02801_),
    .B1(_02800_));
 sg13g2_mux2_1 _10683_ (.A0(_02801_),
    .A1(net2500),
    .S(net1806),
    .X(_00128_));
 sg13g2_nand3_1 _10684_ (.B(_01913_),
    .C(_01914_),
    .A(net2302),
    .Y(_02802_));
 sg13g2_nor3_2 _10685_ (.A(\i_tinyqv.mem.qspi_write_done ),
    .B(_01912_),
    .C(_02589_),
    .Y(_02803_));
 sg13g2_nand2b_2 _10686_ (.Y(_02804_),
    .B(_01913_),
    .A_N(_02589_));
 sg13g2_and3_2 _10687_ (.X(_02805_),
    .A(_01913_),
    .B(_02570_),
    .C(_02589_));
 sg13g2_nor2_2 _10688_ (.A(net2438),
    .B(_02805_),
    .Y(_02806_));
 sg13g2_nor2_2 _10689_ (.A(_02803_),
    .B(_02805_),
    .Y(_02807_));
 sg13g2_nor2_1 _10690_ (.A(net2438),
    .B(_02804_),
    .Y(_02808_));
 sg13g2_nand2_1 _10691_ (.Y(_02809_),
    .A(\addr[0] ),
    .B(net2062));
 sg13g2_and2_1 _10692_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .B(_02418_),
    .X(_02810_));
 sg13g2_nand2_1 _10693_ (.Y(_02811_),
    .A(net2781),
    .B(net1752));
 sg13g2_o21ai_1 _10694_ (.B1(_02809_),
    .Y(_00129_),
    .A1(_02810_),
    .A2(_02811_));
 sg13g2_nor2_2 _10695_ (.A(_01907_),
    .B(_01956_),
    .Y(_02812_));
 sg13g2_and2_1 _10696_ (.A(net2387),
    .B(_02812_),
    .X(_02813_));
 sg13g2_o21ai_1 _10697_ (.B1(net2495),
    .Y(_02814_),
    .A1(net3966),
    .A2(_02813_));
 sg13g2_nand2_2 _10698_ (.Y(_02815_),
    .A(_01360_),
    .B(_02043_));
 sg13g2_inv_1 _10699_ (.Y(_02816_),
    .A(_02815_));
 sg13g2_a21oi_1 _10700_ (.A1(_02813_),
    .A2(_02815_),
    .Y(_00130_),
    .B1(_02814_));
 sg13g2_nor2_2 _10701_ (.A(_01328_),
    .B(_02042_),
    .Y(_02817_));
 sg13g2_inv_4 _10702_ (.A(_02817_),
    .Y(_02818_));
 sg13g2_o21ai_1 _10703_ (.B1(net2495),
    .Y(_02819_),
    .A1(net3910),
    .A2(_02813_));
 sg13g2_a21oi_1 _10704_ (.A1(_02813_),
    .A2(_02818_),
    .Y(_00131_),
    .B1(_02819_));
 sg13g2_nand2_2 _10705_ (.Y(_02820_),
    .A(_01292_),
    .B(_02043_));
 sg13g2_inv_1 _10706_ (.Y(_02821_),
    .A(_02820_));
 sg13g2_o21ai_1 _10707_ (.B1(net2495),
    .Y(_02822_),
    .A1(net4106),
    .A2(_02813_));
 sg13g2_a21oi_2 _10708_ (.B1(_02822_),
    .Y(_00132_),
    .A2(_02820_),
    .A1(_02813_));
 sg13g2_nor2_2 _10709_ (.A(_01254_),
    .B(_02042_),
    .Y(_02823_));
 sg13g2_inv_4 _10710_ (.A(_02823_),
    .Y(_02824_));
 sg13g2_o21ai_1 _10711_ (.B1(net2496),
    .Y(_02825_),
    .A1(net4033),
    .A2(_02813_));
 sg13g2_a21oi_1 _10712_ (.A1(_02813_),
    .A2(_02824_),
    .Y(_00133_),
    .B1(_02825_));
 sg13g2_nor2_1 _10713_ (.A(_01107_),
    .B(\time_limit[2] ),
    .Y(_02826_));
 sg13g2_nand2_2 _10714_ (.Y(_02827_),
    .A(net2737),
    .B(net4081));
 sg13g2_nor2_1 _10715_ (.A(\time_count[5] ),
    .B(_01109_),
    .Y(_02828_));
 sg13g2_a22oi_1 _10716_ (.Y(_02829_),
    .B1(\time_count[5] ),
    .B2(_01109_),
    .A2(\time_limit[2] ),
    .A1(_01107_));
 sg13g2_xnor2_1 _10717_ (.Y(_02830_),
    .A(\time_count[6] ),
    .B(\time_limit[6] ));
 sg13g2_xnor2_1 _10718_ (.Y(_02831_),
    .A(\time_count[3] ),
    .B(\time_limit[3] ));
 sg13g2_xnor2_1 _10719_ (.Y(_02832_),
    .A(\time_count[4] ),
    .B(\time_limit[4] ));
 sg13g2_nand4_1 _10720_ (.B(_02830_),
    .C(_02831_),
    .A(_02829_),
    .Y(_02833_),
    .D(_02832_));
 sg13g2_nor4_2 _10721_ (.A(_02826_),
    .B(_02827_),
    .C(_02828_),
    .Y(_02834_),
    .D(_02833_));
 sg13g2_nor2_2 _10722_ (.A(net3912),
    .B(_02834_),
    .Y(_02835_));
 sg13g2_nand2_1 _10723_ (.Y(_02836_),
    .A(\i_tinyqv.cpu.i_timer.i_mtime.cy ),
    .B(net2235));
 sg13g2_o21ai_1 _10724_ (.B1(_02836_),
    .Y(_02837_),
    .A1(net2235),
    .A2(_02835_));
 sg13g2_and2_1 _10725_ (.A(net3948),
    .B(_02837_),
    .X(_02838_));
 sg13g2_nand2_1 _10726_ (.Y(_02839_),
    .A(net3760),
    .B(_02838_));
 sg13g2_nand2b_2 _10727_ (.Y(_02840_),
    .B(_02812_),
    .A_N(\addr[2] ));
 sg13g2_nand4_1 _10728_ (.B(\i_tinyqv.cpu.i_timer.i_mtime.data[2] ),
    .C(\i_tinyqv.cpu.i_timer.i_mtime.data[3] ),
    .A(net2495),
    .Y(_02841_),
    .D(_02840_));
 sg13g2_nor2_1 _10729_ (.A(net3761),
    .B(_02841_),
    .Y(_00134_));
 sg13g2_nand2b_1 _10730_ (.Y(_02842_),
    .B(\i_tinyqv.cpu.i_timer.i_mtime.data[2] ),
    .A_N(\i_tinyqv.cpu.i_timer.mtimecmp[6] ));
 sg13g2_nor2b_1 _10731_ (.A(\i_tinyqv.cpu.i_timer.i_mtime.data[2] ),
    .B_N(\i_tinyqv.cpu.i_timer.mtimecmp[6] ),
    .Y(_02843_));
 sg13g2_xnor2_1 _10732_ (.Y(_02844_),
    .A(\i_tinyqv.cpu.i_timer.i_mtime.data[2] ),
    .B(\i_tinyqv.cpu.i_timer.mtimecmp[6] ));
 sg13g2_o21ai_1 _10733_ (.B1(_01114_),
    .Y(_02845_),
    .A1(\i_tinyqv.cpu.i_timer.mtimecmp[4] ),
    .A2(_01113_));
 sg13g2_a22oi_1 _10734_ (.Y(_02846_),
    .B1(\i_tinyqv.cpu.i_timer.mtimecmp[4] ),
    .B2(_01113_),
    .A2(_01112_),
    .A1(\i_tinyqv.cpu.i_timer.mtimecmp[5] ));
 sg13g2_a22oi_1 _10735_ (.Y(_02847_),
    .B1(_02845_),
    .B2(_02846_),
    .A2(net3760),
    .A1(_01111_));
 sg13g2_o21ai_1 _10736_ (.B1(_02842_),
    .Y(_02848_),
    .A1(_02843_),
    .A2(_02847_));
 sg13g2_o21ai_1 _10737_ (.B1(_02848_),
    .Y(_02849_),
    .A1(net4038),
    .A2(_01115_));
 sg13g2_a21oi_1 _10738_ (.A1(net4038),
    .A2(_01115_),
    .Y(_02850_),
    .B1(_01385_));
 sg13g2_nand2_1 _10739_ (.Y(_00135_),
    .A(_02849_),
    .B(_02850_));
 sg13g2_xnor2_1 _10740_ (.Y(_02851_),
    .A(_02844_),
    .B(_02847_));
 sg13g2_xnor2_1 _10741_ (.Y(_02852_),
    .A(\i_tinyqv.cpu.i_timer.i_mtime.data[3] ),
    .B(\i_tinyqv.cpu.i_timer.mtimecmp[7] ));
 sg13g2_xnor2_1 _10742_ (.Y(_02853_),
    .A(_02843_),
    .B(_02852_));
 sg13g2_nor3_1 _10743_ (.A(net2230),
    .B(_02851_),
    .C(_02853_),
    .Y(_02854_));
 sg13g2_a21o_1 _10744_ (.A2(net2230),
    .A1(net3973),
    .B1(_02854_),
    .X(_00136_));
 sg13g2_nor2_1 _10745_ (.A(net2237),
    .B(net3913),
    .Y(_00137_));
 sg13g2_o21ai_1 _10746_ (.B1(_01699_),
    .Y(_02855_),
    .A1(_01692_),
    .A2(_01700_));
 sg13g2_nand2_1 _10747_ (.Y(_02856_),
    .A(net2454),
    .B(net1999));
 sg13g2_o21ai_1 _10748_ (.B1(_01695_),
    .Y(_02857_),
    .A1(_01694_),
    .A2(_01697_));
 sg13g2_nand2_1 _10749_ (.Y(_02858_),
    .A(net2452),
    .B(net2003));
 sg13g2_nand2_1 _10750_ (.Y(_02859_),
    .A(net2453),
    .B(net2001));
 sg13g2_nand2_1 _10751_ (.Y(_02860_),
    .A(net2452),
    .B(net2001));
 sg13g2_xor2_1 _10752_ (.B(_02859_),
    .A(_02858_),
    .X(_02861_));
 sg13g2_nand2_1 _10753_ (.Y(_02862_),
    .A(_02857_),
    .B(_02861_));
 sg13g2_xnor2_1 _10754_ (.Y(_02863_),
    .A(_02857_),
    .B(_02861_));
 sg13g2_or2_1 _10755_ (.X(_02864_),
    .B(_02863_),
    .A(_02856_));
 sg13g2_xor2_1 _10756_ (.B(_02863_),
    .A(_02856_),
    .X(_02865_));
 sg13g2_nand2_1 _10757_ (.Y(_02866_),
    .A(_02855_),
    .B(_02865_));
 sg13g2_xnor2_1 _10758_ (.Y(_02867_),
    .A(_02855_),
    .B(_02865_));
 sg13g2_a21oi_1 _10759_ (.A1(_01702_),
    .A2(_01704_),
    .Y(_02868_),
    .B1(_02867_));
 sg13g2_nand3_1 _10760_ (.B(_01704_),
    .C(_02867_),
    .A(_01702_),
    .Y(_02869_));
 sg13g2_nand2b_1 _10761_ (.Y(_02870_),
    .B(_02869_),
    .A_N(_02868_));
 sg13g2_a21oi_1 _10762_ (.A1(_01707_),
    .A2(_01709_),
    .Y(_02871_),
    .B1(_02870_));
 sg13g2_nand3_1 _10763_ (.B(_01709_),
    .C(_02870_),
    .A(_01707_),
    .Y(_02872_));
 sg13g2_nor2b_1 _10764_ (.A(_02871_),
    .B_N(_02872_),
    .Y(_00138_));
 sg13g2_nand2b_1 _10765_ (.Y(_02873_),
    .B(_01694_),
    .A_N(_02860_));
 sg13g2_nand2_1 _10766_ (.Y(_02874_),
    .A(net2453),
    .B(net1999));
 sg13g2_xnor2_1 _10767_ (.Y(_02875_),
    .A(_02873_),
    .B(_02874_));
 sg13g2_a21o_2 _10768_ (.A2(_02864_),
    .A1(_02862_),
    .B1(_02875_),
    .X(_02876_));
 sg13g2_nand3_1 _10769_ (.B(_02864_),
    .C(_02875_),
    .A(_02862_),
    .Y(_02877_));
 sg13g2_nand2_1 _10770_ (.Y(_02878_),
    .A(_02876_),
    .B(_02877_));
 sg13g2_nor2_1 _10771_ (.A(_02866_),
    .B(_02878_),
    .Y(_02879_));
 sg13g2_xor2_1 _10772_ (.B(_02878_),
    .A(_02866_),
    .X(_02880_));
 sg13g2_or2_1 _10773_ (.X(_02881_),
    .B(_02871_),
    .A(_02868_));
 sg13g2_xor2_1 _10774_ (.B(_02881_),
    .A(_02880_),
    .X(_00139_));
 sg13g2_nand2_1 _10775_ (.Y(_02882_),
    .A(net2452),
    .B(net1999));
 sg13g2_a21oi_1 _10776_ (.A1(_01694_),
    .A2(_02874_),
    .Y(_02883_),
    .B1(_02860_));
 sg13g2_nand2b_1 _10777_ (.Y(_02884_),
    .B(_02883_),
    .A_N(_02882_));
 sg13g2_xor2_1 _10778_ (.B(_02883_),
    .A(_02882_),
    .X(_02885_));
 sg13g2_xor2_1 _10779_ (.B(_02885_),
    .A(_02876_),
    .X(_02886_));
 sg13g2_a21oi_1 _10780_ (.A1(_02880_),
    .A2(_02881_),
    .Y(_02887_),
    .B1(_02879_));
 sg13g2_nand2b_1 _10781_ (.Y(_02888_),
    .B(_02886_),
    .A_N(_02887_));
 sg13g2_xnor2_1 _10782_ (.Y(_00140_),
    .A(_02886_),
    .B(_02887_));
 sg13g2_o21ai_1 _10783_ (.B1(_02884_),
    .Y(_02889_),
    .A1(_02876_),
    .A2(_02885_));
 sg13g2_nand2b_1 _10784_ (.Y(_00141_),
    .B(_02888_),
    .A_N(_02889_));
 sg13g2_nor2_2 _10785_ (.A(net2443),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[25] ),
    .Y(_02890_));
 sg13g2_or2_1 _10786_ (.X(_02891_),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[25] ),
    .A(net2443));
 sg13g2_nand2_2 _10787_ (.Y(_02892_),
    .A(_01144_),
    .B(_02890_));
 sg13g2_xnor2_1 _10788_ (.Y(_02893_),
    .A(_01144_),
    .B(_02890_));
 sg13g2_xor2_1 _10789_ (.B(_02892_),
    .A(\i_peripherals.i_user_peri39.stage1_math_rec[27] ),
    .X(_02894_));
 sg13g2_or4_1 _10790_ (.A(net3704),
    .B(net3416),
    .C(net3059),
    .D(_02892_),
    .X(_02895_));
 sg13g2_a21oi_2 _10791_ (.B1(net3395),
    .Y(_02896_),
    .A2(_02895_),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[30] ));
 sg13g2_nor2b_2 _10792_ (.A(_02894_),
    .B_N(_02896_),
    .Y(_02897_));
 sg13g2_nor2b_1 _10793_ (.A(_02893_),
    .B_N(_02897_),
    .Y(_02898_));
 sg13g2_nand2_2 _10794_ (.Y(_02899_),
    .A(net2443),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[25] ));
 sg13g2_and2_1 _10795_ (.A(_02891_),
    .B(_02899_),
    .X(_02900_));
 sg13g2_nand2_2 _10796_ (.Y(_02901_),
    .A(_02891_),
    .B(_02899_));
 sg13g2_and2_1 _10797_ (.A(net2450),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[15] ),
    .X(_02902_));
 sg13g2_a21oi_1 _10798_ (.A1(net2329),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[16] ),
    .Y(_02903_),
    .B1(_02902_));
 sg13g2_mux2_1 _10799_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[14] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[13] ),
    .S(net2450),
    .X(_02904_));
 sg13g2_nor2_1 _10800_ (.A(net2441),
    .B(_02904_),
    .Y(_02905_));
 sg13g2_a21oi_1 _10801_ (.A1(net2441),
    .A2(_02903_),
    .Y(_02906_),
    .B1(_02905_));
 sg13g2_mux2_1 _10802_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[12] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[11] ),
    .S(net2449),
    .X(_02907_));
 sg13g2_and2_1 _10803_ (.A(net2449),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[9] ),
    .X(_02908_));
 sg13g2_a21oi_1 _10804_ (.A1(net2329),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[10] ),
    .Y(_02909_),
    .B1(_02908_));
 sg13g2_nand2_1 _10805_ (.Y(_02910_),
    .A(net2442),
    .B(_02907_));
 sg13g2_o21ai_1 _10806_ (.B1(_02910_),
    .Y(_02911_),
    .A1(net2442),
    .A2(_02909_));
 sg13g2_mux2_1 _10807_ (.A0(_02906_),
    .A1(_02911_),
    .S(_02901_),
    .X(_02912_));
 sg13g2_nor3_2 _10808_ (.A(net4168),
    .B(net3702),
    .C(_01055_),
    .Y(_02913_));
 sg13g2_nand3b_1 _10809_ (.B(_01054_),
    .C(net3022),
    .Y(_02914_),
    .A_N(net4171));
 sg13g2_nand2_1 _10810_ (.Y(_02915_),
    .A(\i_peripherals.i_user_peri39.stage1_math_rec[31] ),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[30] ));
 sg13g2_nor2_1 _10811_ (.A(\i_peripherals.i_user_peri39.stage1_math_rec[29] ),
    .B(_02915_),
    .Y(_02916_));
 sg13g2_nor2_1 _10812_ (.A(_02896_),
    .B(_02916_),
    .Y(_02917_));
 sg13g2_and2_1 _10813_ (.A(_02893_),
    .B(_02897_),
    .X(_02918_));
 sg13g2_mux2_1 _10814_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[8] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[7] ),
    .S(net2449),
    .X(_02919_));
 sg13g2_nand2_1 _10815_ (.Y(_02920_),
    .A(net2442),
    .B(_02919_));
 sg13g2_nand2_1 _10816_ (.Y(_02921_),
    .A(net2329),
    .B(_01143_));
 sg13g2_o21ai_1 _10817_ (.B1(_02921_),
    .Y(_02922_),
    .A1(net2329),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[5] ));
 sg13g2_o21ai_1 _10818_ (.B1(_02920_),
    .Y(_02923_),
    .A1(net2442),
    .A2(_02922_));
 sg13g2_nand2_1 _10819_ (.Y(_02924_),
    .A(net2448),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[3] ));
 sg13g2_o21ai_1 _10820_ (.B1(_02924_),
    .Y(_02925_),
    .A1(net2449),
    .A2(_01141_));
 sg13g2_nand2b_1 _10821_ (.Y(_02926_),
    .B(_02925_),
    .A_N(_02899_));
 sg13g2_nand2_1 _10822_ (.Y(_02927_),
    .A(\i_peripherals.i_user_peri39.stage1_math_rec[1] ),
    .B(net2448));
 sg13g2_o21ai_1 _10823_ (.B1(_02927_),
    .Y(_02928_),
    .A1(_01139_),
    .A2(net2448));
 sg13g2_a22oi_1 _10824_ (.Y(_02929_),
    .B1(_02928_),
    .B2(_02890_),
    .A2(_02923_),
    .A1(net2213));
 sg13g2_nand2_1 _10825_ (.Y(_02930_),
    .A(_02926_),
    .B(_02929_));
 sg13g2_and2_1 _10826_ (.A(_02894_),
    .B(_02896_),
    .X(_02931_));
 sg13g2_and2_1 _10827_ (.A(_02893_),
    .B(_02931_),
    .X(_02932_));
 sg13g2_and2_1 _10828_ (.A(net2451),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[19] ),
    .X(_02933_));
 sg13g2_a21oi_1 _10829_ (.A1(net2329),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[20] ),
    .Y(_02934_),
    .B1(_02933_));
 sg13g2_mux2_1 _10830_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[18] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[17] ),
    .S(net2450),
    .X(_02935_));
 sg13g2_nor2_1 _10831_ (.A(net2441),
    .B(_02935_),
    .Y(_02936_));
 sg13g2_a21oi_1 _10832_ (.A1(net2443),
    .A2(_02934_),
    .Y(_02937_),
    .B1(_02936_));
 sg13g2_nor2_1 _10833_ (.A(net2212),
    .B(_02937_),
    .Y(_02938_));
 sg13g2_nand2_1 _10834_ (.Y(_02939_),
    .A(net2451),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[21] ));
 sg13g2_o21ai_1 _10835_ (.B1(_02939_),
    .Y(_02940_),
    .A1(net2451),
    .A2(_01145_));
 sg13g2_nor3_1 _10836_ (.A(\i_peripherals.i_user_peri39.stage1_math_rec[31] ),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[30] ),
    .C(\i_peripherals.i_user_peri39.stage1_math_rec[29] ),
    .Y(_02941_));
 sg13g2_nor3_1 _10837_ (.A(net2329),
    .B(_01142_),
    .C(_02941_),
    .Y(_02942_));
 sg13g2_a21oi_1 _10838_ (.A1(_01142_),
    .A2(_02940_),
    .Y(_02943_),
    .B1(_02942_));
 sg13g2_a21oi_2 _10839_ (.B1(_02938_),
    .Y(_02944_),
    .A2(_02943_),
    .A1(net2212));
 sg13g2_a22oi_1 _10840_ (.Y(_02945_),
    .B1(net1989),
    .B2(_02930_),
    .A2(_02912_),
    .A1(net1990));
 sg13g2_a221oi_1 _10841_ (.B2(_02944_),
    .C1(net2202),
    .B1(_02932_),
    .A1(net3485),
    .Y(_02946_),
    .A2(net2057));
 sg13g2_o21ai_1 _10842_ (.B1(net2284),
    .Y(_02947_),
    .A1(net3749),
    .A2(net2207));
 sg13g2_a21oi_1 _10843_ (.A1(_02945_),
    .A2(_02946_),
    .Y(_00142_),
    .B1(_02947_));
 sg13g2_and2_1 _10844_ (.A(net2450),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[16] ),
    .X(_02948_));
 sg13g2_a21oi_1 _10845_ (.A1(net2329),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[17] ),
    .Y(_02949_),
    .B1(_02948_));
 sg13g2_mux2_1 _10846_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[15] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[14] ),
    .S(net2447),
    .X(_02950_));
 sg13g2_nor2_1 _10847_ (.A(net2440),
    .B(_02950_),
    .Y(_02951_));
 sg13g2_a21oi_1 _10848_ (.A1(net2444),
    .A2(_02949_),
    .Y(_02952_),
    .B1(_02951_));
 sg13g2_mux2_1 _10849_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[13] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[12] ),
    .S(net2450),
    .X(_02953_));
 sg13g2_and2_1 _10850_ (.A(net2450),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[10] ),
    .X(_02954_));
 sg13g2_a21oi_1 _10851_ (.A1(_01140_),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[11] ),
    .Y(_02955_),
    .B1(_02954_));
 sg13g2_nand2_1 _10852_ (.Y(_02956_),
    .A(net2441),
    .B(_02953_));
 sg13g2_o21ai_1 _10853_ (.B1(_02956_),
    .Y(_02957_),
    .A1(net2441),
    .A2(_02955_));
 sg13g2_mux2_1 _10854_ (.A0(_02952_),
    .A1(_02957_),
    .S(net2211),
    .X(_02958_));
 sg13g2_nor2_1 _10855_ (.A(net2448),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[7] ),
    .Y(_02959_));
 sg13g2_a21oi_1 _10856_ (.A1(net2448),
    .A2(_01143_),
    .Y(_02960_),
    .B1(_02959_));
 sg13g2_mux2_1 _10857_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[9] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[8] ),
    .S(net2449),
    .X(_02961_));
 sg13g2_mux2_1 _10858_ (.A0(_02960_),
    .A1(_02961_),
    .S(net2442),
    .X(_02962_));
 sg13g2_o21ai_1 _10859_ (.B1(_02890_),
    .Y(_02963_),
    .A1(net2448),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[3] ));
 sg13g2_a21oi_1 _10860_ (.A1(_01139_),
    .A2(net2448),
    .Y(_02964_),
    .B1(_02963_));
 sg13g2_nor2_1 _10861_ (.A(net2451),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[5] ),
    .Y(_02965_));
 sg13g2_a21oi_1 _10862_ (.A1(net2448),
    .A2(_01141_),
    .Y(_02966_),
    .B1(_02965_));
 sg13g2_nand2b_1 _10863_ (.Y(_02967_),
    .B(_02966_),
    .A_N(_02899_));
 sg13g2_a21oi_1 _10864_ (.A1(net2213),
    .A2(_02962_),
    .Y(_02968_),
    .B1(_02964_));
 sg13g2_nand2_1 _10865_ (.Y(_02969_),
    .A(_02967_),
    .B(_02968_));
 sg13g2_mux2_1 _10866_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[21] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[20] ),
    .S(net2446),
    .X(_02970_));
 sg13g2_mux2_1 _10867_ (.A0(\i_peripherals.i_user_peri39.stage1_math_rec[19] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[18] ),
    .S(net2447),
    .X(_02971_));
 sg13g2_mux2_1 _10868_ (.A0(_02970_),
    .A1(_02971_),
    .S(_01142_),
    .X(_02972_));
 sg13g2_nand2_1 _10869_ (.Y(_02973_),
    .A(net2211),
    .B(_02972_));
 sg13g2_nand2_1 _10870_ (.Y(_02974_),
    .A(_01142_),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[25] ));
 sg13g2_nor2_1 _10871_ (.A(net2446),
    .B(_02941_),
    .Y(_02975_));
 sg13g2_a21oi_2 _10872_ (.B1(_02975_),
    .Y(_02976_),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[22] ),
    .A1(net2446));
 sg13g2_o21ai_1 _10873_ (.B1(_02973_),
    .Y(_02977_),
    .A1(_02974_),
    .A2(_02976_));
 sg13g2_a22oi_1 _10874_ (.Y(_02978_),
    .B1(_02969_),
    .B2(net1988),
    .A2(_02958_),
    .A1(net1991));
 sg13g2_a221oi_1 _10875_ (.B2(_02977_),
    .C1(net2202),
    .B1(_02932_),
    .A1(net3601),
    .Y(_02979_),
    .A2(net2057));
 sg13g2_o21ai_1 _10876_ (.B1(net2284),
    .Y(_02980_),
    .A1(net3830),
    .A2(net2207));
 sg13g2_a21oi_1 _10877_ (.A1(_02978_),
    .A2(_02979_),
    .Y(_00143_),
    .B1(_02980_));
 sg13g2_nor2_1 _10878_ (.A(net2442),
    .B(_02919_),
    .Y(_02981_));
 sg13g2_a21oi_1 _10879_ (.A1(net2442),
    .A2(_02909_),
    .Y(_02982_),
    .B1(_02981_));
 sg13g2_a22oi_1 _10880_ (.Y(_02983_),
    .B1(_02982_),
    .B2(net2213),
    .A2(_02925_),
    .A1(_02890_));
 sg13g2_o21ai_1 _10881_ (.B1(_02983_),
    .Y(_02984_),
    .A1(_02899_),
    .A2(_02922_));
 sg13g2_nand2_1 _10882_ (.Y(_02985_),
    .A(net2441),
    .B(_02935_));
 sg13g2_o21ai_1 _10883_ (.B1(_02985_),
    .Y(_02986_),
    .A1(net2441),
    .A2(_02903_));
 sg13g2_mux4_1 _10884_ (.S0(net2440),
    .A0(\i_peripherals.i_user_peri39.stage1_math_rec[12] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[14] ),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[11] ),
    .A3(\i_peripherals.i_user_peri39.stage1_math_rec[13] ),
    .S1(net2450),
    .X(_02987_));
 sg13g2_mux2_1 _10885_ (.A0(_02986_),
    .A1(_02987_),
    .S(net2211),
    .X(_02988_));
 sg13g2_nor2_1 _10886_ (.A(_01142_),
    .B(_02940_),
    .Y(_02989_));
 sg13g2_a21oi_1 _10887_ (.A1(_01142_),
    .A2(_02934_),
    .Y(_02990_),
    .B1(_02989_));
 sg13g2_nand2_1 _10888_ (.Y(_02991_),
    .A(net2211),
    .B(_02990_));
 sg13g2_nand2b_1 _10889_ (.Y(_02992_),
    .B(net2446),
    .A_N(_02941_));
 sg13g2_o21ai_1 _10890_ (.B1(_02991_),
    .Y(_02993_),
    .A1(_02974_),
    .A2(_02992_));
 sg13g2_a22oi_1 _10891_ (.Y(_02994_),
    .B1(_02993_),
    .B2(_02932_),
    .A2(_02984_),
    .A1(net1987));
 sg13g2_a221oi_1 _10892_ (.B2(net1990),
    .C1(net2202),
    .B1(_02988_),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[2] ),
    .Y(_02995_),
    .A2(net2057));
 sg13g2_o21ai_1 _10893_ (.B1(net2284),
    .Y(_02996_),
    .A1(net3743),
    .A2(net2207));
 sg13g2_a21oi_1 _10894_ (.A1(_02994_),
    .A2(_02995_),
    .Y(_00144_),
    .B1(_02996_));
 sg13g2_nand2_1 _10895_ (.Y(_02997_),
    .A(net2440),
    .B(_02971_));
 sg13g2_o21ai_1 _10896_ (.B1(_02997_),
    .Y(_02998_),
    .A1(net2444),
    .A2(_02949_));
 sg13g2_mux4_1 _10897_ (.S0(net2440),
    .A0(\i_peripherals.i_user_peri39.stage1_math_rec[13] ),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[15] ),
    .A2(\i_peripherals.i_user_peri39.stage1_math_rec[12] ),
    .A3(\i_peripherals.i_user_peri39.stage1_math_rec[14] ),
    .S1(net2450),
    .X(_02999_));
 sg13g2_mux2_1 _10898_ (.A0(_02998_),
    .A1(_02999_),
    .S(net2211),
    .X(_03000_));
 sg13g2_a221oi_1 _10899_ (.B2(net1990),
    .C1(net2202),
    .B1(_03000_),
    .A1(net3649),
    .Y(_03001_),
    .A2(net2057));
 sg13g2_nor2_1 _10900_ (.A(net2440),
    .B(_02970_),
    .Y(_03002_));
 sg13g2_a21oi_1 _10901_ (.A1(net2440),
    .A2(_02976_),
    .Y(_03003_),
    .B1(_03002_));
 sg13g2_and2_1 _10902_ (.A(net2211),
    .B(_03003_),
    .X(_03004_));
 sg13g2_nor2_1 _10903_ (.A(net2442),
    .B(_02961_),
    .Y(_03005_));
 sg13g2_a21oi_1 _10904_ (.A1(net2441),
    .A2(_02955_),
    .Y(_03006_),
    .B1(_03005_));
 sg13g2_nand2_1 _10905_ (.Y(_03007_),
    .A(net2213),
    .B(_03006_));
 sg13g2_nand2b_1 _10906_ (.Y(_03008_),
    .B(_02960_),
    .A_N(_02899_));
 sg13g2_o21ai_1 _10907_ (.B1(_02966_),
    .Y(_03009_),
    .A1(_01144_),
    .A2(_02890_));
 sg13g2_nand3_1 _10908_ (.B(_03008_),
    .C(_03009_),
    .A(_03007_),
    .Y(_03010_));
 sg13g2_a22oi_1 _10909_ (.Y(_03011_),
    .B1(_03010_),
    .B2(net1988),
    .A2(_03004_),
    .A1(_02932_));
 sg13g2_o21ai_1 _10910_ (.B1(net2285),
    .Y(_03012_),
    .A1(net3834),
    .A2(net2207));
 sg13g2_a21oi_1 _10911_ (.A1(_03001_),
    .A2(_03011_),
    .Y(_00145_),
    .B1(_03012_));
 sg13g2_mux2_1 _10912_ (.A0(_02911_),
    .A1(_02923_),
    .S(_02901_),
    .X(_03013_));
 sg13g2_mux2_1 _10913_ (.A0(_02906_),
    .A1(_02937_),
    .S(net2212),
    .X(_03014_));
 sg13g2_nor2_1 _10914_ (.A(net2212),
    .B(_02943_),
    .Y(_03015_));
 sg13g2_a22oi_1 _10915_ (.Y(_03016_),
    .B1(_03014_),
    .B2(net1991),
    .A2(_03013_),
    .A1(net1988));
 sg13g2_a221oi_1 _10916_ (.B2(_03015_),
    .C1(net2202),
    .B1(_02932_),
    .A1(net3871),
    .Y(_03017_),
    .A2(net2057));
 sg13g2_o21ai_1 _10917_ (.B1(net2284),
    .Y(_03018_),
    .A1(net3927),
    .A2(net2208));
 sg13g2_a21oi_1 _10918_ (.A1(_03016_),
    .A2(_03017_),
    .Y(_00146_),
    .B1(_03018_));
 sg13g2_mux2_1 _10919_ (.A0(_02952_),
    .A1(_02972_),
    .S(net2212),
    .X(_03019_));
 sg13g2_nand2_1 _10920_ (.Y(_03020_),
    .A(net2213),
    .B(_02957_));
 sg13g2_nand2_1 _10921_ (.Y(_03021_),
    .A(net2211),
    .B(_02962_));
 sg13g2_nand3_1 _10922_ (.B(_03020_),
    .C(_03021_),
    .A(_02893_),
    .Y(_03022_));
 sg13g2_nor2_1 _10923_ (.A(_02892_),
    .B(_02976_),
    .Y(_03023_));
 sg13g2_nand2_1 _10924_ (.Y(_03024_),
    .A(\i_peripherals.i_user_peri39.stage1_math_rec[27] ),
    .B(_03023_));
 sg13g2_o21ai_1 _10925_ (.B1(_03022_),
    .Y(_03025_),
    .A1(_02893_),
    .A2(_03019_));
 sg13g2_o21ai_1 _10926_ (.B1(_03024_),
    .Y(_03026_),
    .A1(_02894_),
    .A2(_03025_));
 sg13g2_a221oi_1 _10927_ (.B2(net2115),
    .C1(net2203),
    .B1(_03026_),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[5] ),
    .Y(_03027_),
    .A2(net2056));
 sg13g2_o21ai_1 _10928_ (.B1(net2286),
    .Y(_03028_),
    .A1(net3504),
    .A2(net2206));
 sg13g2_nor2_1 _10929_ (.A(_03027_),
    .B(_03028_),
    .Y(_00147_));
 sg13g2_nor2_1 _10930_ (.A(_02891_),
    .B(_02992_),
    .Y(_03029_));
 sg13g2_nor2_1 _10931_ (.A(_02892_),
    .B(_02992_),
    .Y(_03030_));
 sg13g2_a221oi_1 _10932_ (.B2(_03030_),
    .C1(net2203),
    .B1(_02931_),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[6] ),
    .Y(_03031_),
    .A2(net2056));
 sg13g2_mux2_1 _10933_ (.A0(_02986_),
    .A1(_02990_),
    .S(net2212),
    .X(_03032_));
 sg13g2_mux2_1 _10934_ (.A0(_02982_),
    .A1(_02987_),
    .S(net2212),
    .X(_03033_));
 sg13g2_a22oi_1 _10935_ (.Y(_03034_),
    .B1(_03033_),
    .B2(net1987),
    .A2(_03032_),
    .A1(net1991));
 sg13g2_o21ai_1 _10936_ (.B1(net2284),
    .Y(_03035_),
    .A1(net3692),
    .A2(net2207));
 sg13g2_a21oi_1 _10937_ (.A1(_03031_),
    .A2(_03034_),
    .Y(_00148_),
    .B1(_03035_));
 sg13g2_mux2_1 _10938_ (.A0(_02999_),
    .A1(_03006_),
    .S(net2211),
    .X(_03036_));
 sg13g2_mux2_1 _10939_ (.A0(_02998_),
    .A1(_03003_),
    .S(net2212),
    .X(_03037_));
 sg13g2_a22oi_1 _10940_ (.Y(_03038_),
    .B1(net1988),
    .B2(_03036_),
    .A2(net2058),
    .A1(net3811));
 sg13g2_a21oi_1 _10941_ (.A1(net1990),
    .A2(_03037_),
    .Y(_03039_),
    .B1(net2202));
 sg13g2_o21ai_1 _10942_ (.B1(net2285),
    .Y(_03040_),
    .A1(net3959),
    .A2(net2208));
 sg13g2_a21oi_1 _10943_ (.A1(_03038_),
    .A2(_03039_),
    .Y(_00149_),
    .B1(_03040_));
 sg13g2_a22oi_1 _10944_ (.Y(_03041_),
    .B1(net1989),
    .B2(_02912_),
    .A2(net2058),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[8] ));
 sg13g2_a21oi_1 _10945_ (.A1(net1990),
    .A2(_02944_),
    .Y(_03042_),
    .B1(net2203));
 sg13g2_o21ai_1 _10946_ (.B1(net2284),
    .Y(_03043_),
    .A1(net3679),
    .A2(net2207));
 sg13g2_a21oi_1 _10947_ (.A1(_03041_),
    .A2(_03042_),
    .Y(_00150_),
    .B1(_03043_));
 sg13g2_a22oi_1 _10948_ (.Y(_03044_),
    .B1(_02977_),
    .B2(net1991),
    .A2(net2057),
    .A1(net3750));
 sg13g2_a21oi_1 _10949_ (.A1(net1988),
    .A2(_02958_),
    .Y(_03045_),
    .B1(_02914_));
 sg13g2_o21ai_1 _10950_ (.B1(net2285),
    .Y(_03046_),
    .A1(net4000),
    .A2(net2208));
 sg13g2_a21oi_1 _10951_ (.A1(_03044_),
    .A2(_03045_),
    .Y(_00151_),
    .B1(_03046_));
 sg13g2_a22oi_1 _10952_ (.Y(_03047_),
    .B1(net1989),
    .B2(_02988_),
    .A2(net2058),
    .A1(net3810));
 sg13g2_a21oi_1 _10953_ (.A1(net1990),
    .A2(_02993_),
    .Y(_03048_),
    .B1(net2202));
 sg13g2_o21ai_1 _10954_ (.B1(net2284),
    .Y(_03049_),
    .A1(net3846),
    .A2(net2207));
 sg13g2_a21oi_1 _10955_ (.A1(_03047_),
    .A2(_03048_),
    .Y(_00152_),
    .B1(_03049_));
 sg13g2_a22oi_1 _10956_ (.Y(_03050_),
    .B1(_03004_),
    .B2(net1990),
    .A2(net2058),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[11] ));
 sg13g2_a21oi_1 _10957_ (.A1(net1988),
    .A2(_03000_),
    .Y(_03051_),
    .B1(net2203));
 sg13g2_o21ai_1 _10958_ (.B1(net2284),
    .Y(_03052_),
    .A1(net3733),
    .A2(net2208));
 sg13g2_a21oi_1 _10959_ (.A1(_03050_),
    .A2(_03051_),
    .Y(_00153_),
    .B1(_03052_));
 sg13g2_a22oi_1 _10960_ (.Y(_03053_),
    .B1(_03015_),
    .B2(net1990),
    .A2(net2057),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[12] ));
 sg13g2_a21oi_1 _10961_ (.A1(net1987),
    .A2(_03014_),
    .Y(_03054_),
    .B1(net2202));
 sg13g2_o21ai_1 _10962_ (.B1(net2286),
    .Y(_03055_),
    .A1(net3662),
    .A2(net2207));
 sg13g2_a21oi_1 _10963_ (.A1(_03053_),
    .A2(_03054_),
    .Y(_00154_),
    .B1(_03055_));
 sg13g2_nand3_1 _10964_ (.B(_02890_),
    .C(_02897_),
    .A(net3759),
    .Y(_03056_));
 sg13g2_nor2_1 _10965_ (.A(_02976_),
    .B(_03056_),
    .Y(_03057_));
 sg13g2_a221oi_1 _10966_ (.B2(_03019_),
    .C1(_03057_),
    .B1(net1989),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[13] ),
    .Y(_03058_),
    .A2(net2059));
 sg13g2_o21ai_1 _10967_ (.B1(net2282),
    .Y(_03059_),
    .A1(net3875),
    .A2(net2205));
 sg13g2_a21oi_1 _10968_ (.A1(net2205),
    .A2(_03058_),
    .Y(_00155_),
    .B1(_03059_));
 sg13g2_a21oi_1 _10969_ (.A1(\i_peripherals.i_user_peri39.stage1_math_rec[14] ),
    .A2(net2056),
    .Y(_03060_),
    .B1(net2203));
 sg13g2_a22oi_1 _10970_ (.Y(_03061_),
    .B1(_03032_),
    .B2(net1987),
    .A2(_03029_),
    .A1(net1991));
 sg13g2_o21ai_1 _10971_ (.B1(net2286),
    .Y(_03062_),
    .A1(net3850),
    .A2(net2206));
 sg13g2_a21oi_1 _10972_ (.A1(_03060_),
    .A2(_03061_),
    .Y(_00156_),
    .B1(_03062_));
 sg13g2_a22oi_1 _10973_ (.Y(_03063_),
    .B1(net1988),
    .B2(_03037_),
    .A2(net2058),
    .A1(net3774));
 sg13g2_o21ai_1 _10974_ (.B1(net2281),
    .Y(_03064_),
    .A1(net3794),
    .A2(net2205));
 sg13g2_a21oi_1 _10975_ (.A1(net2205),
    .A2(_03063_),
    .Y(_00157_),
    .B1(_03064_));
 sg13g2_a22oi_1 _10976_ (.Y(_03065_),
    .B1(net1987),
    .B2(_02944_),
    .A2(net2056),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[16] ));
 sg13g2_o21ai_1 _10977_ (.B1(net2286),
    .Y(_03066_),
    .A1(net3855),
    .A2(net2206));
 sg13g2_a21oi_1 _10978_ (.A1(net2206),
    .A2(_03065_),
    .Y(_00158_),
    .B1(_03066_));
 sg13g2_a22oi_1 _10979_ (.Y(_03067_),
    .B1(net1988),
    .B2(_02977_),
    .A2(net2057),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[17] ));
 sg13g2_o21ai_1 _10980_ (.B1(net2281),
    .Y(_03068_),
    .A1(net3858),
    .A2(net2204));
 sg13g2_a21oi_1 _10981_ (.A1(net2204),
    .A2(_03067_),
    .Y(_00159_),
    .B1(_03068_));
 sg13g2_a22oi_1 _10982_ (.Y(_03069_),
    .B1(net1987),
    .B2(_02993_),
    .A2(net2056),
    .A1(net3821));
 sg13g2_o21ai_1 _10983_ (.B1(net2286),
    .Y(_03070_),
    .A1(net3886),
    .A2(net2206));
 sg13g2_a21oi_1 _10984_ (.A1(net2206),
    .A2(_03069_),
    .Y(_00160_),
    .B1(_03070_));
 sg13g2_a22oi_1 _10985_ (.Y(_03071_),
    .B1(net1987),
    .B2(_03004_),
    .A2(net2056),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[19] ));
 sg13g2_o21ai_1 _10986_ (.B1(net2281),
    .Y(_03072_),
    .A1(net3768),
    .A2(net2205));
 sg13g2_a21oi_1 _10987_ (.A1(net2205),
    .A2(_03071_),
    .Y(_00161_),
    .B1(_03072_));
 sg13g2_a22oi_1 _10988_ (.Y(_03073_),
    .B1(net1987),
    .B2(_03015_),
    .A2(net2056),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[20] ));
 sg13g2_o21ai_1 _10989_ (.B1(net2282),
    .Y(_03074_),
    .A1(net3790),
    .A2(net2204));
 sg13g2_a21oi_1 _10990_ (.A1(net2204),
    .A2(_03073_),
    .Y(_00162_),
    .B1(_03074_));
 sg13g2_a221oi_1 _10991_ (.B2(_02897_),
    .C1(net2203),
    .B1(_03023_),
    .A1(\i_peripherals.i_user_peri39.stage1_math_rec[21] ),
    .Y(_03075_),
    .A2(net2059));
 sg13g2_o21ai_1 _10992_ (.B1(net2282),
    .Y(_03076_),
    .A1(net3717),
    .A2(net2205));
 sg13g2_nor2_1 _10993_ (.A(_03075_),
    .B(_03076_),
    .Y(_00163_));
 sg13g2_a221oi_1 _10994_ (.B2(_02897_),
    .C1(net2203),
    .B1(_03030_),
    .A1(net3470),
    .Y(_03077_),
    .A2(net2056));
 sg13g2_o21ai_1 _10995_ (.B1(net2281),
    .Y(_03078_),
    .A1(net3661),
    .A2(net2204));
 sg13g2_nor2_1 _10996_ (.A(_03077_),
    .B(_03078_),
    .Y(_00164_));
 sg13g2_and2_1 _10997_ (.A(net2206),
    .B(_02915_),
    .X(_03079_));
 sg13g2_o21ai_1 _10998_ (.B1(_03079_),
    .Y(_03080_),
    .A1(net2445),
    .A2(net2115));
 sg13g2_o21ai_1 _10999_ (.B1(_03080_),
    .Y(_03081_),
    .A1(net3745),
    .A2(net2204));
 sg13g2_nor2_1 _11000_ (.A(net2252),
    .B(_03081_),
    .Y(_00165_));
 sg13g2_xor2_1 _11001_ (.B(net2440),
    .A(net2445),
    .X(_03082_));
 sg13g2_o21ai_1 _11002_ (.B1(_03079_),
    .Y(_03083_),
    .A1(net2115),
    .A2(_03082_));
 sg13g2_o21ai_1 _11003_ (.B1(net2281),
    .Y(_03084_),
    .A1(net3498),
    .A2(net2204));
 sg13g2_nor2b_1 _11004_ (.A(_03084_),
    .B_N(_03083_),
    .Y(_00166_));
 sg13g2_o21ai_1 _11005_ (.B1(net3430),
    .Y(_03085_),
    .A1(net2445),
    .A2(net2440));
 sg13g2_o21ai_1 _11006_ (.B1(_03085_),
    .Y(_03086_),
    .A1(net2446),
    .A2(_02891_));
 sg13g2_nand2b_1 _11007_ (.Y(_03087_),
    .B(_03086_),
    .A_N(net2115));
 sg13g2_o21ai_1 _11008_ (.B1(net2287),
    .Y(_03088_),
    .A1(net3905),
    .A2(net2210));
 sg13g2_a21oi_1 _11009_ (.A1(_03079_),
    .A2(_03087_),
    .Y(_00167_),
    .B1(_03088_));
 sg13g2_o21ai_1 _11010_ (.B1(net3759),
    .Y(_03089_),
    .A1(net2445),
    .A2(_02891_));
 sg13g2_o21ai_1 _11011_ (.B1(_03089_),
    .Y(_03090_),
    .A1(net2445),
    .A2(_02892_));
 sg13g2_nand2b_1 _11012_ (.Y(_03091_),
    .B(_03090_),
    .A_N(net2115));
 sg13g2_o21ai_1 _11013_ (.B1(net2287),
    .Y(_03092_),
    .A1(net3952),
    .A2(net2210));
 sg13g2_a21oi_1 _11014_ (.A1(_03079_),
    .A2(_03091_),
    .Y(_00168_),
    .B1(_03092_));
 sg13g2_nor3_1 _11015_ (.A(net2445),
    .B(\i_peripherals.i_user_peri39.stage1_math_rec[27] ),
    .C(_02892_),
    .Y(_03093_));
 sg13g2_o21ai_1 _11016_ (.B1(\i_peripherals.i_user_peri39.stage1_math_rec[27] ),
    .Y(_03094_),
    .A1(net2445),
    .A2(_02892_));
 sg13g2_nor2b_1 _11017_ (.A(_03093_),
    .B_N(_03094_),
    .Y(_03095_));
 sg13g2_o21ai_1 _11018_ (.B1(_03079_),
    .Y(_03096_),
    .A1(net2115),
    .A2(_03095_));
 sg13g2_o21ai_1 _11019_ (.B1(net2282),
    .Y(_03097_),
    .A1(net3716),
    .A2(net2205));
 sg13g2_nor2b_1 _11020_ (.A(_03097_),
    .B_N(_03096_),
    .Y(_00169_));
 sg13g2_nor2b_1 _11021_ (.A(net3059),
    .B_N(_03093_),
    .Y(_03098_));
 sg13g2_xnor2_1 _11022_ (.Y(_03099_),
    .A(\i_peripherals.i_user_peri39.stage1_math_rec[28] ),
    .B(_03093_));
 sg13g2_o21ai_1 _11023_ (.B1(_03079_),
    .Y(_03100_),
    .A1(net2115),
    .A2(_03099_));
 sg13g2_o21ai_1 _11024_ (.B1(_03100_),
    .Y(_03101_),
    .A1(net3868),
    .A2(net2204));
 sg13g2_nor2_1 _11025_ (.A(net2252),
    .B(_03101_),
    .Y(_00170_));
 sg13g2_xnor2_1 _11026_ (.Y(_03102_),
    .A(net3416),
    .B(_03098_));
 sg13g2_o21ai_1 _11027_ (.B1(_03079_),
    .Y(_03103_),
    .A1(net2115),
    .A2(_03102_));
 sg13g2_o21ai_1 _11028_ (.B1(net2286),
    .Y(_03104_),
    .A1(net3869),
    .A2(net2209));
 sg13g2_nor2b_1 _11029_ (.A(_03104_),
    .B_N(_03103_),
    .Y(_00171_));
 sg13g2_o21ai_1 _11030_ (.B1(net3395),
    .Y(_03105_),
    .A1(net2445),
    .A2(_02895_));
 sg13g2_o21ai_1 _11031_ (.B1(net2287),
    .Y(_03106_),
    .A1(net3714),
    .A2(net2210));
 sg13g2_a21oi_1 _11032_ (.A1(_03079_),
    .A2(_03105_),
    .Y(_00172_),
    .B1(_03106_));
 sg13g2_o21ai_1 _11033_ (.B1(net2288),
    .Y(_03107_),
    .A1(\i_peripherals.i_user_peri39.math_result_reg[31] ),
    .A2(net2209));
 sg13g2_a21oi_1 _11034_ (.A1(_01064_),
    .A2(net2206),
    .Y(_00173_),
    .B1(_03107_));
 sg13g2_nor3_2 _11035_ (.A(net3937),
    .B(_01054_),
    .C(net3022),
    .Y(_03108_));
 sg13g2_nand3b_1 _11036_ (.B(\i_peripherals.i_user_peri39.busy_counter[1] ),
    .C(_01055_),
    .Y(_03109_),
    .A_N(\i_peripherals.i_user_peri39.busy_counter[2] ));
 sg13g2_nand2b_1 _11037_ (.Y(_03110_),
    .B(\i_peripherals.i_user_peri39.instr[18] ),
    .A_N(\i_peripherals.i_user_peri39.instr[19] ));
 sg13g2_nand2b_1 _11038_ (.Y(_03111_),
    .B(_03110_),
    .A_N(\i_peripherals.i_user_peri39.instr[17] ));
 sg13g2_nor2b_1 _11039_ (.A(\i_peripherals.i_user_peri39.instr[18] ),
    .B_N(\i_peripherals.i_user_peri39.instr[19] ),
    .Y(_03112_));
 sg13g2_nand2b_1 _11040_ (.Y(_03113_),
    .B(\i_peripherals.i_user_peri39.instr[19] ),
    .A_N(\i_peripherals.i_user_peri39.instr[18] ));
 sg13g2_nand2_1 _11041_ (.Y(_03114_),
    .A(\i_peripherals.i_user_peri39.instr[17] ),
    .B(_03113_));
 sg13g2_nand3b_1 _11042_ (.B(\i_peripherals.i_user_peri39.instr[17] ),
    .C(\i_peripherals.i_user_peri39.instr[19] ),
    .Y(_03115_),
    .A_N(\i_peripherals.i_user_peri39.instr[18] ));
 sg13g2_o21ai_1 _11043_ (.B1(_03115_),
    .Y(_03116_),
    .A1(\i_peripherals.i_user_peri39.instr[17] ),
    .A2(_03110_));
 sg13g2_xnor2_1 _11044_ (.Y(_03117_),
    .A(\i_peripherals.i_user_peri39.instr[19] ),
    .B(\i_peripherals.i_user_peri39.instr[18] ));
 sg13g2_xor2_1 _11045_ (.B(\i_peripherals.i_user_peri39.instr[18] ),
    .A(\i_peripherals.i_user_peri39.instr[19] ),
    .X(_03118_));
 sg13g2_mux2_1 _11046_ (.A0(_03113_),
    .A1(_03118_),
    .S(\i_peripherals.i_user_peri39.instr[17] ),
    .X(_03119_));
 sg13g2_mux2_1 _11047_ (.A0(_03112_),
    .A1(_03117_),
    .S(\i_peripherals.i_user_peri39.instr[17] ),
    .X(_03120_));
 sg13g2_mux2_1 _11048_ (.A0(_03120_),
    .A1(_03116_),
    .S(\i_peripherals.i_user_peri39.instr[16] ),
    .X(_03121_));
 sg13g2_nand2_1 _11049_ (.Y(_03122_),
    .A(\i_peripherals.i_user_peri39.instr[15] ),
    .B(_03121_));
 sg13g2_a21o_1 _11050_ (.A2(_03119_),
    .A1(\i_peripherals.i_user_peri39.instr[16] ),
    .B1(_03116_),
    .X(_03123_));
 sg13g2_a221oi_1 _11051_ (.B2(\i_peripherals.i_user_peri39.instr[16] ),
    .C1(_01057_),
    .B1(_03119_),
    .A1(_03111_),
    .Y(_03124_),
    .A2(_03114_));
 sg13g2_mux2_1 _11052_ (.A0(_03124_),
    .A1(_01057_),
    .S(_03121_),
    .X(_03125_));
 sg13g2_o21ai_1 _11053_ (.B1(_03122_),
    .Y(_03126_),
    .A1(_03121_),
    .A2(_03124_));
 sg13g2_a21oi_1 _11054_ (.A1(\i_peripherals.i_user_peri39.instr[16] ),
    .A2(_03116_),
    .Y(_03127_),
    .B1(\i_peripherals.i_user_peri39.instr[15] ));
 sg13g2_nand2_1 _11055_ (.Y(_03128_),
    .A(_03123_),
    .B(_03127_));
 sg13g2_a22oi_1 _11056_ (.Y(_03129_),
    .B1(_03123_),
    .B2(_03127_),
    .A2(_03121_),
    .A1(\i_peripherals.i_user_peri39.instr[15] ));
 sg13g2_nand2_1 _11057_ (.Y(_03130_),
    .A(_03122_),
    .B(_03128_));
 sg13g2_mux2_1 _11058_ (.A0(\i_peripherals.i_user_peri39._GEN[127] ),
    .A1(\i_peripherals.i_user_peri39._GEN[63] ),
    .S(net2113),
    .X(_03131_));
 sg13g2_mux2_1 _11059_ (.A0(\i_peripherals.i_user_peri39._GEN[95] ),
    .A1(_03131_),
    .S(net2106),
    .X(_03132_));
 sg13g2_inv_2 _11060_ (.Y(_03133_),
    .A(_03132_));
 sg13g2_nand2b_1 _11061_ (.Y(_03134_),
    .B(\i_peripherals.i_user_peri39.instr[23] ),
    .A_N(\i_peripherals.i_user_peri39.instr[24] ));
 sg13g2_nand2b_1 _11062_ (.Y(_03135_),
    .B(_03134_),
    .A_N(\i_peripherals.i_user_peri39.instr[22] ));
 sg13g2_nor2b_1 _11063_ (.A(\i_peripherals.i_user_peri39.instr[23] ),
    .B_N(\i_peripherals.i_user_peri39.instr[24] ),
    .Y(_03136_));
 sg13g2_nand2b_1 _11064_ (.Y(_03137_),
    .B(\i_peripherals.i_user_peri39.instr[24] ),
    .A_N(\i_peripherals.i_user_peri39.instr[23] ));
 sg13g2_nand2_1 _11065_ (.Y(_03138_),
    .A(\i_peripherals.i_user_peri39.instr[22] ),
    .B(_03137_));
 sg13g2_nand3b_1 _11066_ (.B(\i_peripherals.i_user_peri39.instr[22] ),
    .C(\i_peripherals.i_user_peri39.instr[24] ),
    .Y(_03139_),
    .A_N(\i_peripherals.i_user_peri39.instr[23] ));
 sg13g2_o21ai_1 _11067_ (.B1(_03139_),
    .Y(_03140_),
    .A1(\i_peripherals.i_user_peri39.instr[22] ),
    .A2(_03134_));
 sg13g2_xnor2_1 _11068_ (.Y(_03141_),
    .A(\i_peripherals.i_user_peri39.instr[24] ),
    .B(\i_peripherals.i_user_peri39.instr[23] ));
 sg13g2_xor2_1 _11069_ (.B(\i_peripherals.i_user_peri39.instr[23] ),
    .A(\i_peripherals.i_user_peri39.instr[24] ),
    .X(_03142_));
 sg13g2_mux2_1 _11070_ (.A0(_03137_),
    .A1(_03142_),
    .S(\i_peripherals.i_user_peri39.instr[22] ),
    .X(_03143_));
 sg13g2_mux2_1 _11071_ (.A0(_03136_),
    .A1(_03141_),
    .S(\i_peripherals.i_user_peri39.instr[22] ),
    .X(_03144_));
 sg13g2_mux2_1 _11072_ (.A0(_03144_),
    .A1(_03140_),
    .S(\i_peripherals.i_user_peri39.instr[21] ),
    .X(_03145_));
 sg13g2_and2_1 _11073_ (.A(\i_peripherals.i_user_peri39.instr[20] ),
    .B(_03145_),
    .X(_03146_));
 sg13g2_a21o_1 _11074_ (.A2(_03143_),
    .A1(\i_peripherals.i_user_peri39.instr[21] ),
    .B1(_03140_),
    .X(_03147_));
 sg13g2_a221oi_1 _11075_ (.B2(\i_peripherals.i_user_peri39.instr[21] ),
    .C1(_01056_),
    .B1(_03143_),
    .A1(_03135_),
    .Y(_03148_),
    .A2(_03138_));
 sg13g2_mux2_1 _11076_ (.A0(_03148_),
    .A1(_01056_),
    .S(_03145_),
    .X(_03149_));
 sg13g2_nand2b_1 _11077_ (.Y(_03150_),
    .B(net2103),
    .A_N(\i_peripherals.i_user_peri39._GEN[63] ));
 sg13g2_a21oi_1 _11078_ (.A1(\i_peripherals.i_user_peri39.instr[21] ),
    .A2(_03140_),
    .Y(_03151_),
    .B1(\i_peripherals.i_user_peri39.instr[20] ));
 sg13g2_a22oi_1 _11079_ (.Y(_03152_),
    .B1(_03147_),
    .B2(_03151_),
    .A2(_03145_),
    .A1(\i_peripherals.i_user_peri39.instr[20] ));
 sg13g2_a21o_2 _11080_ (.A2(_03151_),
    .A1(_03147_),
    .B1(_03146_),
    .X(_03153_));
 sg13g2_o21ai_1 _11081_ (.B1(_03150_),
    .Y(_03154_),
    .A1(\i_peripherals.i_user_peri39._GEN[127] ),
    .A2(net2103));
 sg13g2_nand2_1 _11082_ (.Y(_03155_),
    .A(\i_peripherals.i_user_peri39._GEN[95] ),
    .B(net2050));
 sg13g2_o21ai_1 _11083_ (.B1(_03155_),
    .Y(_03156_),
    .A1(net2050),
    .A2(_03154_));
 sg13g2_xnor2_1 _11084_ (.Y(_03157_),
    .A(_03133_),
    .B(_03156_));
 sg13g2_xnor2_1 _11085_ (.Y(_03158_),
    .A(_03132_),
    .B(_03156_));
 sg13g2_mux2_1 _11086_ (.A0(\i_peripherals.i_user_peri39._GEN[124] ),
    .A1(\i_peripherals.i_user_peri39._GEN[60] ),
    .S(net2101),
    .X(_03159_));
 sg13g2_nor2_1 _11087_ (.A(net2050),
    .B(_03159_),
    .Y(_03160_));
 sg13g2_a21oi_2 _11088_ (.B1(_03160_),
    .Y(_03161_),
    .A2(net2050),
    .A1(_01084_));
 sg13g2_mux2_1 _11089_ (.A0(\i_peripherals.i_user_peri39._GEN[125] ),
    .A1(\i_peripherals.i_user_peri39._GEN[61] ),
    .S(net2105),
    .X(_03162_));
 sg13g2_nor2_1 _11090_ (.A(net2051),
    .B(_03162_),
    .Y(_03163_));
 sg13g2_a21oi_2 _11091_ (.B1(_03163_),
    .Y(_03164_),
    .A2(net2051),
    .A1(_01085_));
 sg13g2_mux2_1 _11092_ (.A0(\i_peripherals.i_user_peri39._GEN[119] ),
    .A1(\i_peripherals.i_user_peri39._GEN[55] ),
    .S(net2102),
    .X(_03165_));
 sg13g2_mux2_1 _11093_ (.A0(\i_peripherals.i_user_peri39._GEN[87] ),
    .A1(_03165_),
    .S(net2096),
    .X(_03166_));
 sg13g2_mux2_1 _11094_ (.A0(\i_peripherals.i_user_peri39._GEN[121] ),
    .A1(\i_peripherals.i_user_peri39._GEN[57] ),
    .S(net2102),
    .X(_03167_));
 sg13g2_nor2_1 _11095_ (.A(net2050),
    .B(_03167_),
    .Y(_03168_));
 sg13g2_a21oi_2 _11096_ (.B1(_03168_),
    .Y(_03169_),
    .A2(net2050),
    .A1(_01082_));
 sg13g2_mux2_1 _11097_ (.A0(\i_peripherals.i_user_peri39._GEN[120] ),
    .A1(\i_peripherals.i_user_peri39._GEN[56] ),
    .S(net2102),
    .X(_03170_));
 sg13g2_mux2_1 _11098_ (.A0(\i_peripherals.i_user_peri39._GEN[88] ),
    .A1(_03170_),
    .S(net2100),
    .X(_03171_));
 sg13g2_mux2_1 _11099_ (.A0(\i_peripherals.i_user_peri39._GEN[122] ),
    .A1(\i_peripherals.i_user_peri39._GEN[58] ),
    .S(net2101),
    .X(_03172_));
 sg13g2_mux2_1 _11100_ (.A0(\i_peripherals.i_user_peri39._GEN[90] ),
    .A1(_03172_),
    .S(net2096),
    .X(_03173_));
 sg13g2_mux2_1 _11101_ (.A0(\i_peripherals.i_user_peri39._GEN[123] ),
    .A1(\i_peripherals.i_user_peri39._GEN[59] ),
    .S(net2103),
    .X(_03174_));
 sg13g2_nor2_1 _11102_ (.A(net2051),
    .B(_03174_),
    .Y(_03175_));
 sg13g2_a21oi_1 _11103_ (.A1(_01081_),
    .A2(net2051),
    .Y(_03176_),
    .B1(_03175_));
 sg13g2_mux2_1 _11104_ (.A0(\i_peripherals.i_user_peri39._GEN[126] ),
    .A1(\i_peripherals.i_user_peri39._GEN[62] ),
    .S(net2103),
    .X(_03177_));
 sg13g2_nor2_1 _11105_ (.A(net2051),
    .B(_03177_),
    .Y(_03178_));
 sg13g2_a21oi_2 _11106_ (.B1(_03178_),
    .Y(_03179_),
    .A2(net2051),
    .A1(_01086_));
 sg13g2_nor4_1 _11107_ (.A(_03161_),
    .B(_03171_),
    .C(_03173_),
    .D(_03176_),
    .Y(_03180_));
 sg13g2_nor4_1 _11108_ (.A(_03164_),
    .B(_03166_),
    .C(_03169_),
    .D(_03179_),
    .Y(_03181_));
 sg13g2_nand2_1 _11109_ (.Y(_03182_),
    .A(_03180_),
    .B(_03181_));
 sg13g2_inv_1 _11110_ (.Y(_03183_),
    .A(net1938));
 sg13g2_nor2_1 _11111_ (.A(_03179_),
    .B(net1926),
    .Y(_03184_));
 sg13g2_nand2b_1 _11112_ (.Y(_03185_),
    .B(net1938),
    .A_N(_03161_));
 sg13g2_mux2_1 _11113_ (.A0(\i_peripherals.i_user_peri39._GEN[117] ),
    .A1(\i_peripherals.i_user_peri39._GEN[53] ),
    .S(net2101),
    .X(_03186_));
 sg13g2_mux2_1 _11114_ (.A0(\i_peripherals.i_user_peri39._GEN[85] ),
    .A1(_03186_),
    .S(net2096),
    .X(_03187_));
 sg13g2_inv_1 _11115_ (.Y(_03188_),
    .A(_03187_));
 sg13g2_mux2_1 _11116_ (.A0(\i_peripherals.i_user_peri39._GEN[118] ),
    .A1(\i_peripherals.i_user_peri39._GEN[54] ),
    .S(net2101),
    .X(_03189_));
 sg13g2_mux2_1 _11117_ (.A0(\i_peripherals.i_user_peri39._GEN[86] ),
    .A1(_03189_),
    .S(net2096),
    .X(_03190_));
 sg13g2_inv_1 _11118_ (.Y(_03191_),
    .A(_03190_));
 sg13g2_nor2_1 _11119_ (.A(_03187_),
    .B(_03190_),
    .Y(_03192_));
 sg13g2_inv_2 _11120_ (.Y(_03193_),
    .A(_03192_));
 sg13g2_mux2_1 _11121_ (.A0(\i_peripherals.i_user_peri39._GEN[115] ),
    .A1(\i_peripherals.i_user_peri39._GEN[51] ),
    .S(net2101),
    .X(_03194_));
 sg13g2_mux2_1 _11122_ (.A0(\i_peripherals.i_user_peri39._GEN[83] ),
    .A1(_03194_),
    .S(net2096),
    .X(_03195_));
 sg13g2_inv_1 _11123_ (.Y(_03196_),
    .A(_03195_));
 sg13g2_mux2_1 _11124_ (.A0(\i_peripherals.i_user_peri39._GEN[116] ),
    .A1(\i_peripherals.i_user_peri39._GEN[52] ),
    .S(net2101),
    .X(_03197_));
 sg13g2_mux2_1 _11125_ (.A0(\i_peripherals.i_user_peri39._GEN[84] ),
    .A1(_03197_),
    .S(net2096),
    .X(_03198_));
 sg13g2_inv_1 _11126_ (.Y(_03199_),
    .A(_03198_));
 sg13g2_nor2_1 _11127_ (.A(_03195_),
    .B(_03198_),
    .Y(_03200_));
 sg13g2_inv_1 _11128_ (.Y(_03201_),
    .A(_03200_));
 sg13g2_mux2_1 _11129_ (.A0(\i_peripherals.i_user_peri39._GEN[113] ),
    .A1(\i_peripherals.i_user_peri39._GEN[49] ),
    .S(net2101),
    .X(_03202_));
 sg13g2_mux2_1 _11130_ (.A0(\i_peripherals.i_user_peri39._GEN[81] ),
    .A1(_03202_),
    .S(net2096),
    .X(_03203_));
 sg13g2_inv_2 _11131_ (.Y(_03204_),
    .A(_03203_));
 sg13g2_mux2_1 _11132_ (.A0(\i_peripherals.i_user_peri39._GEN[114] ),
    .A1(\i_peripherals.i_user_peri39._GEN[50] ),
    .S(net2103),
    .X(_03205_));
 sg13g2_mux2_1 _11133_ (.A0(\i_peripherals.i_user_peri39._GEN[82] ),
    .A1(_03205_),
    .S(net2099),
    .X(_03206_));
 sg13g2_inv_2 _11134_ (.Y(_03207_),
    .A(_03206_));
 sg13g2_nor2_2 _11135_ (.A(_03203_),
    .B(_03206_),
    .Y(_03208_));
 sg13g2_mux2_1 _11136_ (.A0(\i_peripherals.i_user_peri39._GEN[111] ),
    .A1(\i_peripherals.i_user_peri39._GEN[47] ),
    .S(net2101),
    .X(_03209_));
 sg13g2_nor2_1 _11137_ (.A(net2050),
    .B(_03209_),
    .Y(_03210_));
 sg13g2_a21oi_2 _11138_ (.B1(_03210_),
    .Y(_03211_),
    .A2(net2050),
    .A1(_01079_));
 sg13g2_mux2_1 _11139_ (.A0(\i_peripherals.i_user_peri39._GEN[112] ),
    .A1(\i_peripherals.i_user_peri39._GEN[48] ),
    .S(net2103),
    .X(_03212_));
 sg13g2_mux2_1 _11140_ (.A0(\i_peripherals.i_user_peri39._GEN[80] ),
    .A1(_03212_),
    .S(net2099),
    .X(_03213_));
 sg13g2_nor2_1 _11141_ (.A(_03211_),
    .B(_03213_),
    .Y(_03214_));
 sg13g2_mux2_1 _11142_ (.A0(\i_peripherals.i_user_peri39._GEN[109] ),
    .A1(\i_peripherals.i_user_peri39._GEN[45] ),
    .S(net2103),
    .X(_03215_));
 sg13g2_mux2_1 _11143_ (.A0(\i_peripherals.i_user_peri39._GEN[77] ),
    .A1(_03215_),
    .S(net2099),
    .X(_03216_));
 sg13g2_inv_2 _11144_ (.Y(_03217_),
    .A(_03216_));
 sg13g2_mux2_1 _11145_ (.A0(\i_peripherals.i_user_peri39._GEN[110] ),
    .A1(\i_peripherals.i_user_peri39._GEN[46] ),
    .S(net2103),
    .X(_03218_));
 sg13g2_mux2_1 _11146_ (.A0(\i_peripherals.i_user_peri39._GEN[78] ),
    .A1(_03218_),
    .S(net2099),
    .X(_03219_));
 sg13g2_inv_2 _11147_ (.Y(_03220_),
    .A(_03219_));
 sg13g2_nand2_1 _11148_ (.Y(_03221_),
    .A(_03217_),
    .B(_03220_));
 sg13g2_mux2_1 _11149_ (.A0(\i_peripherals.i_user_peri39._GEN[108] ),
    .A1(\i_peripherals.i_user_peri39._GEN[44] ),
    .S(net2104),
    .X(_03222_));
 sg13g2_mux2_1 _11150_ (.A0(\i_peripherals.i_user_peri39._GEN[76] ),
    .A1(_03222_),
    .S(net2098),
    .X(_03223_));
 sg13g2_mux2_1 _11151_ (.A0(\i_peripherals.i_user_peri39._GEN[107] ),
    .A1(\i_peripherals.i_user_peri39._GEN[43] ),
    .S(net2105),
    .X(_03224_));
 sg13g2_mux2_1 _11152_ (.A0(\i_peripherals.i_user_peri39._GEN[75] ),
    .A1(_03224_),
    .S(net2097),
    .X(_03225_));
 sg13g2_or2_1 _11153_ (.X(_03226_),
    .B(_03225_),
    .A(_03223_));
 sg13g2_mux2_1 _11154_ (.A0(\i_peripherals.i_user_peri39._GEN[105] ),
    .A1(\i_peripherals.i_user_peri39._GEN[41] ),
    .S(net2102),
    .X(_03227_));
 sg13g2_mux2_1 _11155_ (.A0(\i_peripherals.i_user_peri39._GEN[73] ),
    .A1(_03227_),
    .S(net2100),
    .X(_03228_));
 sg13g2_inv_1 _11156_ (.Y(_03229_),
    .A(_03228_));
 sg13g2_mux2_1 _11157_ (.A0(\i_peripherals.i_user_peri39._GEN[106] ),
    .A1(\i_peripherals.i_user_peri39._GEN[42] ),
    .S(net2104),
    .X(_03230_));
 sg13g2_mux2_1 _11158_ (.A0(\i_peripherals.i_user_peri39._GEN[74] ),
    .A1(_03230_),
    .S(net2098),
    .X(_03231_));
 sg13g2_inv_1 _11159_ (.Y(_03232_),
    .A(_03231_));
 sg13g2_nor2_1 _11160_ (.A(_03228_),
    .B(_03231_),
    .Y(_03233_));
 sg13g2_mux2_1 _11161_ (.A0(\i_peripherals.i_user_peri39._GEN[103] ),
    .A1(\i_peripherals.i_user_peri39._GEN[39] ),
    .S(net2102),
    .X(_03234_));
 sg13g2_mux2_1 _11162_ (.A0(\i_peripherals.i_user_peri39._GEN[71] ),
    .A1(_03234_),
    .S(net2096),
    .X(_03235_));
 sg13g2_mux2_1 _11163_ (.A0(\i_peripherals.i_user_peri39._GEN[104] ),
    .A1(\i_peripherals.i_user_peri39._GEN[40] ),
    .S(net2104),
    .X(_03236_));
 sg13g2_mux2_1 _11164_ (.A0(\i_peripherals.i_user_peri39._GEN[72] ),
    .A1(_03236_),
    .S(net2098),
    .X(_03237_));
 sg13g2_nor2_1 _11165_ (.A(_03235_),
    .B(_03237_),
    .Y(_03238_));
 sg13g2_mux2_1 _11166_ (.A0(\i_peripherals.i_user_peri39._GEN[101] ),
    .A1(\i_peripherals.i_user_peri39._GEN[37] ),
    .S(net2105),
    .X(_03239_));
 sg13g2_mux2_1 _11167_ (.A0(\i_peripherals.i_user_peri39._GEN[69] ),
    .A1(_03239_),
    .S(net2097),
    .X(_03240_));
 sg13g2_inv_2 _11168_ (.Y(_03241_),
    .A(_03240_));
 sg13g2_mux2_1 _11169_ (.A0(\i_peripherals.i_user_peri39._GEN[102] ),
    .A1(\i_peripherals.i_user_peri39._GEN[38] ),
    .S(net2104),
    .X(_03242_));
 sg13g2_mux2_1 _11170_ (.A0(\i_peripherals.i_user_peri39._GEN[70] ),
    .A1(_03242_),
    .S(net2098),
    .X(_03243_));
 sg13g2_inv_1 _11171_ (.Y(_03244_),
    .A(_03243_));
 sg13g2_or2_1 _11172_ (.X(_03245_),
    .B(_03243_),
    .A(_03240_));
 sg13g2_mux2_1 _11173_ (.A0(\i_peripherals.i_user_peri39._GEN[100] ),
    .A1(\i_peripherals.i_user_peri39._GEN[36] ),
    .S(net2102),
    .X(_03246_));
 sg13g2_mux2_1 _11174_ (.A0(\i_peripherals.i_user_peri39._GEN[68] ),
    .A1(_03246_),
    .S(net2100),
    .X(_03247_));
 sg13g2_mux2_1 _11175_ (.A0(\i_peripherals.i_user_peri39._GEN[3] ),
    .A1(\i_peripherals.i_user_peri39._GEN[35] ),
    .S(net2104),
    .X(_03248_));
 sg13g2_or2_1 _11176_ (.X(_03249_),
    .B(_03248_),
    .A(net2051));
 sg13g2_or2_1 _11177_ (.X(_03250_),
    .B(net2097),
    .A(\i_peripherals.i_user_peri39._GEN[67] ));
 sg13g2_mux2_1 _11178_ (.A0(\i_peripherals.i_user_peri39._GEN[67] ),
    .A1(_03248_),
    .S(net2097),
    .X(_03251_));
 sg13g2_nor2b_1 _11179_ (.A(net2097),
    .B_N(\i_peripherals.i_user_peri39._GEN[65] ),
    .Y(_03252_));
 sg13g2_mux2_1 _11180_ (.A0(\i_peripherals.i_user_peri39._GEN[1] ),
    .A1(\i_peripherals.i_user_peri39._GEN[33] ),
    .S(net2104),
    .X(_03253_));
 sg13g2_a21oi_2 _11181_ (.B1(_03252_),
    .Y(_03254_),
    .A2(_03253_),
    .A1(net2097));
 sg13g2_a21o_1 _11182_ (.A2(_03253_),
    .A1(net2097),
    .B1(_03252_),
    .X(_03255_));
 sg13g2_or2_1 _11183_ (.X(_03256_),
    .B(net2099),
    .A(\i_peripherals.i_user_peri39._GEN[66] ));
 sg13g2_mux2_1 _11184_ (.A0(\i_peripherals.i_user_peri39._GEN[2] ),
    .A1(\i_peripherals.i_user_peri39._GEN[34] ),
    .S(net2104),
    .X(_03257_));
 sg13g2_mux2_1 _11185_ (.A0(\i_peripherals.i_user_peri39._GEN[66] ),
    .A1(_03257_),
    .S(net2099),
    .X(_03258_));
 sg13g2_o21ai_1 _11186_ (.B1(_03256_),
    .Y(_03259_),
    .A1(net2051),
    .A2(_03257_));
 sg13g2_nand2_1 _11187_ (.Y(_03260_),
    .A(_03254_),
    .B(_03259_));
 sg13g2_a221oi_1 _11188_ (.B2(_03259_),
    .C1(_03247_),
    .B1(_03254_),
    .A1(_03249_),
    .Y(_03261_),
    .A2(_03250_));
 sg13g2_o21ai_1 _11189_ (.B1(_03238_),
    .Y(_03262_),
    .A1(_03245_),
    .A2(_03261_));
 sg13g2_a21oi_1 _11190_ (.A1(_03233_),
    .A2(_03262_),
    .Y(_03263_),
    .B1(_03226_));
 sg13g2_o21ai_1 _11191_ (.B1(_03214_),
    .Y(_03264_),
    .A1(_03221_),
    .A2(_03263_));
 sg13g2_a21oi_2 _11192_ (.B1(_03201_),
    .Y(_03265_),
    .A2(_03264_),
    .A1(_03208_));
 sg13g2_nor2_2 _11193_ (.A(_03193_),
    .B(_03265_),
    .Y(_03266_));
 sg13g2_nor3_1 _11194_ (.A(net1938),
    .B(_03193_),
    .C(_03265_),
    .Y(_03267_));
 sg13g2_nor2_1 _11195_ (.A(_03171_),
    .B(_03267_),
    .Y(_03268_));
 sg13g2_o21ai_1 _11196_ (.B1(_03166_),
    .Y(_03269_),
    .A1(_03171_),
    .A2(_03267_));
 sg13g2_o21ai_1 _11197_ (.B1(net1926),
    .Y(_03270_),
    .A1(_03193_),
    .A2(_03265_));
 sg13g2_nor2_1 _11198_ (.A(_03193_),
    .B(_03201_),
    .Y(_03271_));
 sg13g2_inv_1 _11199_ (.Y(_03272_),
    .A(_03271_));
 sg13g2_and2_1 _11200_ (.A(_03208_),
    .B(_03214_),
    .X(_03273_));
 sg13g2_nor2_1 _11201_ (.A(_03221_),
    .B(_03226_),
    .Y(_03274_));
 sg13g2_or3_1 _11202_ (.A(_03245_),
    .B(_03247_),
    .C(_03251_),
    .X(_03275_));
 sg13g2_nand3_1 _11203_ (.B(_03238_),
    .C(_03275_),
    .A(_03233_),
    .Y(_03276_));
 sg13g2_nand2_1 _11204_ (.Y(_03277_),
    .A(_03274_),
    .B(_03276_));
 sg13g2_a21oi_2 _11205_ (.B1(_03272_),
    .Y(_03278_),
    .A2(_03277_),
    .A1(_03273_));
 sg13g2_inv_1 _11206_ (.Y(_03279_),
    .A(net1923));
 sg13g2_a21oi_1 _11207_ (.A1(net1926),
    .A2(net1908),
    .Y(_03280_),
    .B1(_03169_));
 sg13g2_a21oi_2 _11208_ (.B1(_03280_),
    .Y(_03281_),
    .A2(_03270_),
    .A1(_03269_));
 sg13g2_nand3_1 _11209_ (.B(_03238_),
    .C(_03274_),
    .A(_03233_),
    .Y(_03282_));
 sg13g2_and2_1 _11210_ (.A(_03271_),
    .B(_03273_),
    .X(_03283_));
 sg13g2_and2_1 _11211_ (.A(_03282_),
    .B(_03283_),
    .X(_03284_));
 sg13g2_nand2_2 _11212_ (.Y(_03285_),
    .A(_03282_),
    .B(_03283_));
 sg13g2_a21oi_1 _11213_ (.A1(net1926),
    .A2(_03285_),
    .Y(_03286_),
    .B1(_03173_));
 sg13g2_nand2b_1 _11214_ (.Y(_03287_),
    .B(_03281_),
    .A_N(_03286_));
 sg13g2_nand2b_2 _11215_ (.Y(_03288_),
    .B(_03283_),
    .A_N(_03282_));
 sg13g2_nand2_1 _11216_ (.Y(_03289_),
    .A(net1927),
    .B(_03288_));
 sg13g2_a21oi_1 _11217_ (.A1(net1926),
    .A2(_03288_),
    .Y(_03290_),
    .B1(_03176_));
 sg13g2_or2_1 _11218_ (.X(_03291_),
    .B(_03290_),
    .A(_03287_));
 sg13g2_nor2b_2 _11219_ (.A(_03291_),
    .B_N(_03185_),
    .Y(_03292_));
 sg13g2_nor2_1 _11220_ (.A(_03164_),
    .B(_03183_),
    .Y(_03293_));
 sg13g2_nand2b_1 _11221_ (.Y(_03294_),
    .B(_03292_),
    .A_N(_03293_));
 sg13g2_nand2_1 _11222_ (.Y(_03295_),
    .A(_03184_),
    .B(_03294_));
 sg13g2_nand2_2 _11223_ (.Y(_03296_),
    .A(net1939),
    .B(_03295_));
 sg13g2_nand2_1 _11224_ (.Y(_03297_),
    .A(\i_peripherals.i_user_peri39._GEN[59] ),
    .B(net2113));
 sg13g2_a21oi_1 _11225_ (.A1(\i_peripherals.i_user_peri39._GEN[123] ),
    .A2(_03126_),
    .Y(_03298_),
    .B1(net2053));
 sg13g2_a22oi_1 _11226_ (.Y(_03299_),
    .B1(_03297_),
    .B2(_03298_),
    .A2(net2053),
    .A1(_01081_));
 sg13g2_mux2_1 _11227_ (.A0(\i_peripherals.i_user_peri39._GEN[119] ),
    .A1(\i_peripherals.i_user_peri39._GEN[55] ),
    .S(net2111),
    .X(_03300_));
 sg13g2_mux2_1 _11228_ (.A0(\i_peripherals.i_user_peri39._GEN[87] ),
    .A1(_03300_),
    .S(net2109),
    .X(_03301_));
 sg13g2_inv_1 _11229_ (.Y(_03302_),
    .A(_03301_));
 sg13g2_nand2_1 _11230_ (.Y(_03303_),
    .A(\i_peripherals.i_user_peri39._GEN[57] ),
    .B(net2111));
 sg13g2_a21oi_1 _11231_ (.A1(\i_peripherals.i_user_peri39._GEN[121] ),
    .A2(net2055),
    .Y(_03304_),
    .B1(net2052));
 sg13g2_a22oi_1 _11232_ (.Y(_03305_),
    .B1(_03303_),
    .B2(_03304_),
    .A2(net2054),
    .A1(_01082_));
 sg13g2_nand2_1 _11233_ (.Y(_03306_),
    .A(\i_peripherals.i_user_peri39._GEN[126] ),
    .B(_03126_));
 sg13g2_a21oi_1 _11234_ (.A1(\i_peripherals.i_user_peri39._GEN[62] ),
    .A2(net2113),
    .Y(_03307_),
    .B1(net2054));
 sg13g2_a22oi_1 _11235_ (.Y(_03308_),
    .B1(_03306_),
    .B2(_03307_),
    .A2(net2053),
    .A1(_01086_));
 sg13g2_nor4_1 _11236_ (.A(_03299_),
    .B(_03301_),
    .C(_03305_),
    .D(_03308_),
    .Y(_03309_));
 sg13g2_nand2_1 _11237_ (.Y(_03310_),
    .A(\i_peripherals.i_user_peri39._GEN[125] ),
    .B(net2055));
 sg13g2_a21oi_1 _11238_ (.A1(\i_peripherals.i_user_peri39._GEN[61] ),
    .A2(net2113),
    .Y(_03311_),
    .B1(net2053));
 sg13g2_a22oi_1 _11239_ (.Y(_03312_),
    .B1(_03310_),
    .B2(_03311_),
    .A2(net2053),
    .A1(_01085_));
 sg13g2_nand2_1 _11240_ (.Y(_03313_),
    .A(\i_peripherals.i_user_peri39._GEN[58] ),
    .B(net2110));
 sg13g2_a21oi_1 _11241_ (.A1(\i_peripherals.i_user_peri39._GEN[122] ),
    .A2(net2055),
    .Y(_03314_),
    .B1(net2052));
 sg13g2_a22oi_1 _11242_ (.Y(_03315_),
    .B1(_03313_),
    .B2(_03314_),
    .A2(net2054),
    .A1(_01083_));
 sg13g2_nand2_1 _11243_ (.Y(_03316_),
    .A(\i_peripherals.i_user_peri39._GEN[124] ),
    .B(net2055));
 sg13g2_a21oi_1 _11244_ (.A1(\i_peripherals.i_user_peri39._GEN[60] ),
    .A2(net2110),
    .Y(_03317_),
    .B1(net2052));
 sg13g2_a22oi_1 _11245_ (.Y(_03318_),
    .B1(_03316_),
    .B2(_03317_),
    .A2(net2054),
    .A1(_01084_));
 sg13g2_mux2_1 _11246_ (.A0(\i_peripherals.i_user_peri39._GEN[120] ),
    .A1(\i_peripherals.i_user_peri39._GEN[56] ),
    .S(net2111),
    .X(_03319_));
 sg13g2_mux2_1 _11247_ (.A0(\i_peripherals.i_user_peri39._GEN[88] ),
    .A1(_03319_),
    .S(net2106),
    .X(_03320_));
 sg13g2_inv_1 _11248_ (.Y(_03321_),
    .A(_03320_));
 sg13g2_nor4_1 _11249_ (.A(_03312_),
    .B(_03315_),
    .C(_03318_),
    .D(_03320_),
    .Y(_03322_));
 sg13g2_nand2_1 _11250_ (.Y(_03323_),
    .A(_03309_),
    .B(_03322_));
 sg13g2_inv_1 _11251_ (.Y(_03324_),
    .A(net1933));
 sg13g2_nor2_1 _11252_ (.A(_03312_),
    .B(net1925),
    .Y(_03325_));
 sg13g2_nor2_1 _11253_ (.A(_03318_),
    .B(net1925),
    .Y(_03326_));
 sg13g2_mux2_1 _11254_ (.A0(\i_peripherals.i_user_peri39._GEN[117] ),
    .A1(\i_peripherals.i_user_peri39._GEN[53] ),
    .S(net2110),
    .X(_03327_));
 sg13g2_mux2_1 _11255_ (.A0(\i_peripherals.i_user_peri39._GEN[85] ),
    .A1(_03327_),
    .S(net2109),
    .X(_03328_));
 sg13g2_inv_1 _11256_ (.Y(_03329_),
    .A(_03328_));
 sg13g2_mux2_1 _11257_ (.A0(\i_peripherals.i_user_peri39._GEN[118] ),
    .A1(\i_peripherals.i_user_peri39._GEN[54] ),
    .S(net2110),
    .X(_03330_));
 sg13g2_mux2_1 _11258_ (.A0(\i_peripherals.i_user_peri39._GEN[86] ),
    .A1(_03330_),
    .S(net2109),
    .X(_03331_));
 sg13g2_nor2_1 _11259_ (.A(_03328_),
    .B(_03331_),
    .Y(_03332_));
 sg13g2_nand2_1 _11260_ (.Y(_03333_),
    .A(\i_peripherals.i_user_peri39._GEN[51] ),
    .B(net2110));
 sg13g2_a21oi_1 _11261_ (.A1(\i_peripherals.i_user_peri39._GEN[115] ),
    .A2(net2055),
    .Y(_03334_),
    .B1(net2052));
 sg13g2_a22oi_1 _11262_ (.Y(_03335_),
    .B1(_03333_),
    .B2(_03334_),
    .A2(net2052),
    .A1(_01080_));
 sg13g2_mux2_1 _11263_ (.A0(\i_peripherals.i_user_peri39._GEN[116] ),
    .A1(\i_peripherals.i_user_peri39._GEN[52] ),
    .S(net2110),
    .X(_03336_));
 sg13g2_mux2_1 _11264_ (.A0(\i_peripherals.i_user_peri39._GEN[84] ),
    .A1(_03336_),
    .S(net2109),
    .X(_03337_));
 sg13g2_nor2_1 _11265_ (.A(_03335_),
    .B(_03337_),
    .Y(_03338_));
 sg13g2_inv_1 _11266_ (.Y(_03339_),
    .A(_03338_));
 sg13g2_nor2_1 _11267_ (.A(\i_peripherals.i_user_peri39._GEN[49] ),
    .B(net2055),
    .Y(_03340_));
 sg13g2_o21ai_1 _11268_ (.B1(net2109),
    .Y(_03341_),
    .A1(\i_peripherals.i_user_peri39._GEN[113] ),
    .A2(net2110));
 sg13g2_nand2_1 _11269_ (.Y(_03342_),
    .A(\i_peripherals.i_user_peri39._GEN[81] ),
    .B(net2052));
 sg13g2_o21ai_1 _11270_ (.B1(_03342_),
    .Y(_03343_),
    .A1(_03340_),
    .A2(_03341_));
 sg13g2_inv_1 _11271_ (.Y(_03344_),
    .A(_03343_));
 sg13g2_mux2_1 _11272_ (.A0(\i_peripherals.i_user_peri39._GEN[114] ),
    .A1(\i_peripherals.i_user_peri39._GEN[50] ),
    .S(net2113),
    .X(_03345_));
 sg13g2_mux2_1 _11273_ (.A0(\i_peripherals.i_user_peri39._GEN[82] ),
    .A1(_03345_),
    .S(net2108),
    .X(_03346_));
 sg13g2_inv_1 _11274_ (.Y(_03347_),
    .A(_03346_));
 sg13g2_nor2_1 _11275_ (.A(_03343_),
    .B(_03346_),
    .Y(_03348_));
 sg13g2_inv_1 _11276_ (.Y(_03349_),
    .A(_03348_));
 sg13g2_nand2_1 _11277_ (.Y(_03350_),
    .A(\i_peripherals.i_user_peri39._GEN[47] ),
    .B(net2110));
 sg13g2_a21oi_1 _11278_ (.A1(\i_peripherals.i_user_peri39._GEN[111] ),
    .A2(net2055),
    .Y(_03351_),
    .B1(net2052));
 sg13g2_a22oi_1 _11279_ (.Y(_03352_),
    .B1(_03350_),
    .B2(_03351_),
    .A2(net2052),
    .A1(_01079_));
 sg13g2_mux2_1 _11280_ (.A0(\i_peripherals.i_user_peri39._GEN[112] ),
    .A1(\i_peripherals.i_user_peri39._GEN[48] ),
    .S(net2113),
    .X(_03353_));
 sg13g2_mux2_1 _11281_ (.A0(\i_peripherals.i_user_peri39._GEN[80] ),
    .A1(_03353_),
    .S(net2108),
    .X(_03354_));
 sg13g2_nor2_1 _11282_ (.A(_03352_),
    .B(_03354_),
    .Y(_03355_));
 sg13g2_mux2_1 _11283_ (.A0(\i_peripherals.i_user_peri39._GEN[109] ),
    .A1(\i_peripherals.i_user_peri39._GEN[45] ),
    .S(net2113),
    .X(_03356_));
 sg13g2_mux2_1 _11284_ (.A0(\i_peripherals.i_user_peri39._GEN[77] ),
    .A1(_03356_),
    .S(net2108),
    .X(_03357_));
 sg13g2_inv_1 _11285_ (.Y(_03358_),
    .A(_03357_));
 sg13g2_mux2_1 _11286_ (.A0(\i_peripherals.i_user_peri39._GEN[110] ),
    .A1(\i_peripherals.i_user_peri39._GEN[46] ),
    .S(net2113),
    .X(_03359_));
 sg13g2_mux2_1 _11287_ (.A0(\i_peripherals.i_user_peri39._GEN[78] ),
    .A1(_03359_),
    .S(net2108),
    .X(_03360_));
 sg13g2_inv_2 _11288_ (.Y(_03361_),
    .A(_03360_));
 sg13g2_nand2_1 _11289_ (.Y(_03362_),
    .A(_03358_),
    .B(_03361_));
 sg13g2_mux2_1 _11290_ (.A0(\i_peripherals.i_user_peri39._GEN[108] ),
    .A1(\i_peripherals.i_user_peri39._GEN[44] ),
    .S(net2112),
    .X(_03363_));
 sg13g2_mux2_1 _11291_ (.A0(\i_peripherals.i_user_peri39._GEN[76] ),
    .A1(_03363_),
    .S(net2106),
    .X(_03364_));
 sg13g2_mux2_1 _11292_ (.A0(\i_peripherals.i_user_peri39._GEN[107] ),
    .A1(\i_peripherals.i_user_peri39._GEN[43] ),
    .S(net2114),
    .X(_03365_));
 sg13g2_mux2_1 _11293_ (.A0(\i_peripherals.i_user_peri39._GEN[75] ),
    .A1(_03365_),
    .S(net2107),
    .X(_03366_));
 sg13g2_nor2_1 _11294_ (.A(_03364_),
    .B(_03366_),
    .Y(_03367_));
 sg13g2_mux2_1 _11295_ (.A0(\i_peripherals.i_user_peri39._GEN[106] ),
    .A1(\i_peripherals.i_user_peri39._GEN[42] ),
    .S(net2114),
    .X(_03368_));
 sg13g2_mux2_1 _11296_ (.A0(\i_peripherals.i_user_peri39._GEN[74] ),
    .A1(_03368_),
    .S(net2106),
    .X(_03369_));
 sg13g2_inv_1 _11297_ (.Y(_03370_),
    .A(_03369_));
 sg13g2_mux2_1 _11298_ (.A0(\i_peripherals.i_user_peri39._GEN[105] ),
    .A1(\i_peripherals.i_user_peri39._GEN[41] ),
    .S(net2111),
    .X(_03371_));
 sg13g2_mux2_1 _11299_ (.A0(\i_peripherals.i_user_peri39._GEN[73] ),
    .A1(_03371_),
    .S(net2109),
    .X(_03372_));
 sg13g2_inv_1 _11300_ (.Y(_03373_),
    .A(_03372_));
 sg13g2_nor2_1 _11301_ (.A(_03369_),
    .B(_03372_),
    .Y(_03374_));
 sg13g2_nor2_1 _11302_ (.A(\i_peripherals.i_user_peri39._GEN[40] ),
    .B(net2055),
    .Y(_03375_));
 sg13g2_o21ai_1 _11303_ (.B1(net2107),
    .Y(_03376_),
    .A1(\i_peripherals.i_user_peri39._GEN[104] ),
    .A2(net2112));
 sg13g2_nand2_1 _11304_ (.Y(_03377_),
    .A(\i_peripherals.i_user_peri39._GEN[72] ),
    .B(net2053));
 sg13g2_o21ai_1 _11305_ (.B1(_03377_),
    .Y(_03378_),
    .A1(_03375_),
    .A2(_03376_));
 sg13g2_mux2_1 _11306_ (.A0(\i_peripherals.i_user_peri39._GEN[103] ),
    .A1(\i_peripherals.i_user_peri39._GEN[39] ),
    .S(net2111),
    .X(_03379_));
 sg13g2_mux2_1 _11307_ (.A0(\i_peripherals.i_user_peri39._GEN[71] ),
    .A1(_03379_),
    .S(net2109),
    .X(_03380_));
 sg13g2_nor2_1 _11308_ (.A(_03378_),
    .B(_03380_),
    .Y(_03381_));
 sg13g2_or2_1 _11309_ (.X(_03382_),
    .B(_03380_),
    .A(_03378_));
 sg13g2_mux2_1 _11310_ (.A0(\i_peripherals.i_user_peri39._GEN[101] ),
    .A1(\i_peripherals.i_user_peri39._GEN[37] ),
    .S(net2114),
    .X(_03383_));
 sg13g2_mux2_1 _11311_ (.A0(\i_peripherals.i_user_peri39._GEN[69] ),
    .A1(_03383_),
    .S(net2107),
    .X(_03384_));
 sg13g2_inv_1 _11312_ (.Y(_03385_),
    .A(_03384_));
 sg13g2_mux2_1 _11313_ (.A0(\i_peripherals.i_user_peri39._GEN[102] ),
    .A1(\i_peripherals.i_user_peri39._GEN[38] ),
    .S(net2112),
    .X(_03386_));
 sg13g2_mux2_1 _11314_ (.A0(\i_peripherals.i_user_peri39._GEN[70] ),
    .A1(_03386_),
    .S(net2106),
    .X(_03387_));
 sg13g2_inv_1 _11315_ (.Y(_03388_),
    .A(_03387_));
 sg13g2_or2_1 _11316_ (.X(_03389_),
    .B(_03387_),
    .A(_03384_));
 sg13g2_mux2_1 _11317_ (.A0(\i_peripherals.i_user_peri39._GEN[100] ),
    .A1(\i_peripherals.i_user_peri39._GEN[36] ),
    .S(net2112),
    .X(_03390_));
 sg13g2_mux2_1 _11318_ (.A0(\i_peripherals.i_user_peri39._GEN[68] ),
    .A1(_03390_),
    .S(net2106),
    .X(_03391_));
 sg13g2_mux2_1 _11319_ (.A0(\i_peripherals.i_user_peri39._GEN[3] ),
    .A1(\i_peripherals.i_user_peri39._GEN[35] ),
    .S(net2112),
    .X(_03392_));
 sg13g2_mux2_1 _11320_ (.A0(\i_peripherals.i_user_peri39._GEN[67] ),
    .A1(_03392_),
    .S(net2106),
    .X(_03393_));
 sg13g2_nor2_1 _11321_ (.A(_03391_),
    .B(_03393_),
    .Y(_03394_));
 sg13g2_mux2_1 _11322_ (.A0(\i_peripherals.i_user_peri39._GEN[1] ),
    .A1(\i_peripherals.i_user_peri39._GEN[33] ),
    .S(net2112),
    .X(_03395_));
 sg13g2_mux2_1 _11323_ (.A0(\i_peripherals.i_user_peri39._GEN[65] ),
    .A1(_03395_),
    .S(net2106),
    .X(_03396_));
 sg13g2_mux2_1 _11324_ (.A0(\i_peripherals.i_user_peri39._GEN[2] ),
    .A1(\i_peripherals.i_user_peri39._GEN[34] ),
    .S(net2112),
    .X(_03397_));
 sg13g2_nor2_1 _11325_ (.A(net2053),
    .B(_03397_),
    .Y(_03398_));
 sg13g2_or2_1 _11326_ (.X(_03399_),
    .B(net2108),
    .A(\i_peripherals.i_user_peri39._GEN[66] ));
 sg13g2_nor2b_1 _11327_ (.A(_03398_),
    .B_N(_03399_),
    .Y(_03400_));
 sg13g2_o21ai_1 _11328_ (.B1(_03399_),
    .Y(_03401_),
    .A1(net2053),
    .A2(_03397_));
 sg13g2_nand2b_1 _11329_ (.Y(_03402_),
    .B(_03401_),
    .A_N(_03396_));
 sg13g2_a21oi_1 _11330_ (.A1(_03394_),
    .A2(_03402_),
    .Y(_03403_),
    .B1(_03389_));
 sg13g2_o21ai_1 _11331_ (.B1(_03374_),
    .Y(_03404_),
    .A1(_03382_),
    .A2(_03403_));
 sg13g2_a21o_1 _11332_ (.A2(_03404_),
    .A1(_03367_),
    .B1(_03362_),
    .X(_03405_));
 sg13g2_a21oi_1 _11333_ (.A1(_03355_),
    .A2(_03405_),
    .Y(_03406_),
    .B1(_03349_));
 sg13g2_o21ai_1 _11334_ (.B1(_03332_),
    .Y(_03407_),
    .A1(_03339_),
    .A2(_03406_));
 sg13g2_inv_2 _11335_ (.Y(_03408_),
    .A(net1902));
 sg13g2_o21ai_1 _11336_ (.B1(_03321_),
    .Y(_03409_),
    .A1(net1933),
    .A2(_03407_));
 sg13g2_a22oi_1 _11337_ (.Y(_03410_),
    .B1(_03409_),
    .B2(_03301_),
    .A2(_03407_),
    .A1(net1925));
 sg13g2_and2_1 _11338_ (.A(_03332_),
    .B(_03338_),
    .X(_03411_));
 sg13g2_inv_1 _11339_ (.Y(_03412_),
    .A(_03411_));
 sg13g2_and2_1 _11340_ (.A(_03348_),
    .B(_03355_),
    .X(_03413_));
 sg13g2_nor2b_1 _11341_ (.A(_03362_),
    .B_N(_03367_),
    .Y(_03414_));
 sg13g2_nand2b_1 _11342_ (.Y(_03415_),
    .B(_03394_),
    .A_N(_03389_));
 sg13g2_nand3_1 _11343_ (.B(_03381_),
    .C(_03415_),
    .A(_03374_),
    .Y(_03416_));
 sg13g2_nand2_1 _11344_ (.Y(_03417_),
    .A(_03414_),
    .B(_03416_));
 sg13g2_a21oi_1 _11345_ (.A1(_03413_),
    .A2(_03417_),
    .Y(_03418_),
    .B1(_03412_));
 sg13g2_nor2_2 _11346_ (.A(net1928),
    .B(net1916),
    .Y(_03419_));
 sg13g2_nor2_1 _11347_ (.A(_03305_),
    .B(_03419_),
    .Y(_03420_));
 sg13g2_nand2_2 _11348_ (.Y(_03421_),
    .A(_03411_),
    .B(_03413_));
 sg13g2_nand3_1 _11349_ (.B(_03381_),
    .C(_03414_),
    .A(_03374_),
    .Y(_03422_));
 sg13g2_nor2b_1 _11350_ (.A(_03421_),
    .B_N(_03422_),
    .Y(_03423_));
 sg13g2_nand2b_2 _11351_ (.Y(_03424_),
    .B(_03422_),
    .A_N(_03421_));
 sg13g2_a21oi_1 _11352_ (.A1(net1925),
    .A2(_03424_),
    .Y(_03425_),
    .B1(_03315_));
 sg13g2_or3_1 _11353_ (.A(_03410_),
    .B(_03420_),
    .C(_03425_),
    .X(_03426_));
 sg13g2_nor2_2 _11354_ (.A(_03421_),
    .B(_03422_),
    .Y(_03427_));
 sg13g2_nor2_2 _11355_ (.A(net1929),
    .B(_03427_),
    .Y(_03428_));
 sg13g2_o21ai_1 _11356_ (.B1(net1924),
    .Y(_03429_),
    .A1(_03421_),
    .A2(_03422_));
 sg13g2_nor2_2 _11357_ (.A(_03299_),
    .B(_03428_),
    .Y(_03430_));
 sg13g2_nor2_1 _11358_ (.A(_03426_),
    .B(_03430_),
    .Y(_03431_));
 sg13g2_nor3_1 _11359_ (.A(_03326_),
    .B(_03426_),
    .C(_03430_),
    .Y(_03432_));
 sg13g2_nor2b_2 _11360_ (.A(_03325_),
    .B_N(_03432_),
    .Y(_03433_));
 sg13g2_nor2_1 _11361_ (.A(_03308_),
    .B(net1925),
    .Y(_03434_));
 sg13g2_o21ai_1 _11362_ (.B1(net1933),
    .Y(_03435_),
    .A1(_03308_),
    .A2(_03433_));
 sg13g2_a21oi_1 _11363_ (.A1(net1939),
    .A2(_03295_),
    .Y(_03436_),
    .B1(_03435_));
 sg13g2_nand2b_2 _11364_ (.Y(_03437_),
    .B(_03296_),
    .A_N(_03435_));
 sg13g2_xor2_1 _11365_ (.B(_03434_),
    .A(_03433_),
    .X(_03438_));
 sg13g2_xor2_1 _11366_ (.B(_03294_),
    .A(_03184_),
    .X(_03439_));
 sg13g2_nand2_1 _11367_ (.Y(_03440_),
    .A(_03438_),
    .B(_03439_));
 sg13g2_mux2_1 _11368_ (.A0(\i_peripherals.i_user_peri39._GEN[0] ),
    .A1(\i_peripherals.i_user_peri39._GEN[32] ),
    .S(net2104),
    .X(_03441_));
 sg13g2_mux2_1 _11369_ (.A0(\i_peripherals.i_user_peri39._GEN[64] ),
    .A1(_03441_),
    .S(net2097),
    .X(_03442_));
 sg13g2_nor4_1 _11370_ (.A(_03260_),
    .B(_03275_),
    .C(_03288_),
    .D(_03442_),
    .Y(_03443_));
 sg13g2_nand4_1 _11371_ (.B(_03179_),
    .C(net1939),
    .A(_03164_),
    .Y(_03444_),
    .D(_03292_));
 sg13g2_nand2_2 _11372_ (.Y(_03445_),
    .A(net1926),
    .B(_03443_));
 sg13g2_xnor2_1 _11373_ (.Y(_03446_),
    .A(_03292_),
    .B(_03293_));
 sg13g2_nand2_1 _11374_ (.Y(_03447_),
    .A(_03445_),
    .B(_03446_));
 sg13g2_o21ai_1 _11375_ (.B1(_03447_),
    .Y(_03448_),
    .A1(_03443_),
    .A2(_03444_));
 sg13g2_mux2_1 _11376_ (.A0(\i_peripherals.i_user_peri39._GEN[0] ),
    .A1(\i_peripherals.i_user_peri39._GEN[32] ),
    .S(net2112),
    .X(_03449_));
 sg13g2_mux2_1 _11377_ (.A0(\i_peripherals.i_user_peri39._GEN[64] ),
    .A1(_03449_),
    .S(net2107),
    .X(_03450_));
 sg13g2_nor3_1 _11378_ (.A(_03402_),
    .B(_03415_),
    .C(_03450_),
    .Y(_03451_));
 sg13g2_and2_1 _11379_ (.A(_03427_),
    .B(_03451_),
    .X(_03452_));
 sg13g2_nand2_2 _11380_ (.Y(_03453_),
    .A(net1925),
    .B(_03452_));
 sg13g2_nand3_1 _11381_ (.B(net1933),
    .C(_03433_),
    .A(_03308_),
    .Y(_03454_));
 sg13g2_nor2_1 _11382_ (.A(_03452_),
    .B(_03454_),
    .Y(_03455_));
 sg13g2_xnor2_1 _11383_ (.Y(_03456_),
    .A(_03325_),
    .B(_03432_));
 sg13g2_o21ai_1 _11384_ (.B1(_03453_),
    .Y(_03457_),
    .A1(_03455_),
    .A2(_03456_));
 sg13g2_nor2_1 _11385_ (.A(_03448_),
    .B(_03457_),
    .Y(_03458_));
 sg13g2_or2_1 _11386_ (.X(_03459_),
    .B(_03457_),
    .A(_03448_));
 sg13g2_xnor2_1 _11387_ (.Y(_03460_),
    .A(_03448_),
    .B(_03457_));
 sg13g2_xnor2_1 _11388_ (.Y(_03461_),
    .A(_03185_),
    .B(_03291_));
 sg13g2_xnor2_1 _11389_ (.Y(_03462_),
    .A(_03326_),
    .B(_03431_));
 sg13g2_nor2b_1 _11390_ (.A(_03461_),
    .B_N(_03462_),
    .Y(_03463_));
 sg13g2_nor2b_2 _11391_ (.A(_03462_),
    .B_N(_03461_),
    .Y(_03464_));
 sg13g2_xor2_1 _11392_ (.B(_03430_),
    .A(_03426_),
    .X(_03465_));
 sg13g2_xor2_1 _11393_ (.B(_03290_),
    .A(_03287_),
    .X(_03466_));
 sg13g2_nor2b_1 _11394_ (.A(_03466_),
    .B_N(_03465_),
    .Y(_03467_));
 sg13g2_xnor2_1 _11395_ (.Y(_03468_),
    .A(_03465_),
    .B(_03466_));
 sg13g2_xor2_1 _11396_ (.B(_03286_),
    .A(_03281_),
    .X(_03469_));
 sg13g2_o21ai_1 _11397_ (.B1(_03425_),
    .Y(_03470_),
    .A1(_03410_),
    .A2(_03420_));
 sg13g2_and2_1 _11398_ (.A(_03426_),
    .B(_03470_),
    .X(_03471_));
 sg13g2_and2_1 _11399_ (.A(_03469_),
    .B(_03471_),
    .X(_03472_));
 sg13g2_or2_1 _11400_ (.X(_03473_),
    .B(_03471_),
    .A(_03469_));
 sg13g2_xor2_1 _11401_ (.B(_03420_),
    .A(_03410_),
    .X(_03474_));
 sg13g2_nand3_1 _11402_ (.B(_03270_),
    .C(_03280_),
    .A(_03269_),
    .Y(_03475_));
 sg13g2_nor2b_2 _11403_ (.A(_03281_),
    .B_N(_03475_),
    .Y(_03476_));
 sg13g2_nand2b_1 _11404_ (.Y(_03477_),
    .B(_03474_),
    .A_N(_03476_));
 sg13g2_nor2b_1 _11405_ (.A(_03474_),
    .B_N(_03476_),
    .Y(_03478_));
 sg13g2_xnor2_1 _11406_ (.Y(_03479_),
    .A(_03474_),
    .B(_03476_));
 sg13g2_xnor2_1 _11407_ (.Y(_03480_),
    .A(_03166_),
    .B(_03268_));
 sg13g2_xnor2_1 _11408_ (.Y(_03481_),
    .A(_03301_),
    .B(_03409_));
 sg13g2_nor2_2 _11409_ (.A(_03480_),
    .B(_03481_),
    .Y(_03482_));
 sg13g2_nand2_1 _11410_ (.Y(_03483_),
    .A(_03480_),
    .B(_03481_));
 sg13g2_nand2_1 _11411_ (.Y(_03484_),
    .A(_03187_),
    .B(_03191_));
 sg13g2_a21oi_1 _11412_ (.A1(_03255_),
    .A2(_03259_),
    .Y(_03485_),
    .B1(_03251_));
 sg13g2_o21ai_1 _11413_ (.B1(_03241_),
    .Y(_03486_),
    .A1(_03247_),
    .A2(_03485_));
 sg13g2_a21oi_1 _11414_ (.A1(_03244_),
    .A2(_03486_),
    .Y(_03487_),
    .B1(_03235_));
 sg13g2_o21ai_1 _11415_ (.B1(_03229_),
    .Y(_03488_),
    .A1(_03237_),
    .A2(_03487_));
 sg13g2_a21oi_1 _11416_ (.A1(_03232_),
    .A2(_03488_),
    .Y(_03489_),
    .B1(_03225_));
 sg13g2_o21ai_1 _11417_ (.B1(_03217_),
    .Y(_03490_),
    .A1(_03223_),
    .A2(_03489_));
 sg13g2_a21oi_1 _11418_ (.A1(_03220_),
    .A2(_03490_),
    .Y(_03491_),
    .B1(_03211_));
 sg13g2_o21ai_1 _11419_ (.B1(_03204_),
    .Y(_03492_),
    .A1(_03213_),
    .A2(_03491_));
 sg13g2_a21oi_1 _11420_ (.A1(_03207_),
    .A2(_03492_),
    .Y(_03493_),
    .B1(_03195_));
 sg13g2_nand2_1 _11421_ (.Y(_03494_),
    .A(_03191_),
    .B(_03199_));
 sg13g2_o21ai_1 _11422_ (.B1(_03484_),
    .Y(_03495_),
    .A1(_03493_),
    .A2(_03494_));
 sg13g2_a21oi_2 _11423_ (.B1(_03166_),
    .Y(_03496_),
    .A2(net1889),
    .A1(net1926));
 sg13g2_nor2_1 _11424_ (.A(_03329_),
    .B(_03331_),
    .Y(_03497_));
 sg13g2_a21oi_1 _11425_ (.A1(_03396_),
    .A2(_03401_),
    .Y(_03498_),
    .B1(_03393_));
 sg13g2_o21ai_1 _11426_ (.B1(_03385_),
    .Y(_03499_),
    .A1(_03391_),
    .A2(_03498_));
 sg13g2_a21oi_1 _11427_ (.A1(_03388_),
    .A2(_03499_),
    .Y(_03500_),
    .B1(_03380_));
 sg13g2_o21ai_1 _11428_ (.B1(_03373_),
    .Y(_03501_),
    .A1(_03378_),
    .A2(_03500_));
 sg13g2_a21oi_1 _11429_ (.A1(_03370_),
    .A2(_03501_),
    .Y(_03502_),
    .B1(_03366_));
 sg13g2_o21ai_1 _11430_ (.B1(_03358_),
    .Y(_03503_),
    .A1(_03364_),
    .A2(_03502_));
 sg13g2_a21oi_1 _11431_ (.A1(_03361_),
    .A2(_03503_),
    .Y(_03504_),
    .B1(_03352_));
 sg13g2_o21ai_1 _11432_ (.B1(_03344_),
    .Y(_03505_),
    .A1(_03354_),
    .A2(_03504_));
 sg13g2_a21o_1 _11433_ (.A2(_03505_),
    .A1(_03347_),
    .B1(_03335_),
    .X(_03506_));
 sg13g2_or2_1 _11434_ (.X(_03507_),
    .B(_03337_),
    .A(_03331_));
 sg13g2_inv_1 _11435_ (.Y(_03508_),
    .A(_03507_));
 sg13g2_a21oi_1 _11436_ (.A1(_03506_),
    .A2(_03508_),
    .Y(_03509_),
    .B1(_03497_));
 sg13g2_o21ai_1 _11437_ (.B1(_03302_),
    .Y(_03510_),
    .A1(net1933),
    .A2(net1884));
 sg13g2_nand2_2 _11438_ (.Y(_03511_),
    .A(_03496_),
    .B(_03510_));
 sg13g2_nor2b_2 _11439_ (.A(_03482_),
    .B_N(_03483_),
    .Y(_03512_));
 sg13g2_inv_1 _11440_ (.Y(_03513_),
    .A(_03512_));
 sg13g2_a21oi_1 _11441_ (.A1(_03496_),
    .A2(_03510_),
    .Y(_03514_),
    .B1(_03513_));
 sg13g2_o21ai_1 _11442_ (.B1(_03479_),
    .Y(_03515_),
    .A1(_03482_),
    .A2(_03514_));
 sg13g2_nand2_1 _11443_ (.Y(_03516_),
    .A(_03477_),
    .B(_03515_));
 sg13g2_nand3b_1 _11444_ (.B(_03477_),
    .C(_03515_),
    .Y(_03517_),
    .A_N(_03472_));
 sg13g2_and3_1 _11445_ (.X(_03518_),
    .A(_03468_),
    .B(_03473_),
    .C(_03517_));
 sg13g2_nor2_1 _11446_ (.A(_03467_),
    .B(_03518_),
    .Y(_03519_));
 sg13g2_nor3_1 _11447_ (.A(_03463_),
    .B(_03467_),
    .C(_03518_),
    .Y(_03520_));
 sg13g2_nor3_1 _11448_ (.A(_03460_),
    .B(_03464_),
    .C(_03520_),
    .Y(_03521_));
 sg13g2_or3_1 _11449_ (.A(_03460_),
    .B(_03464_),
    .C(_03520_),
    .X(_03522_));
 sg13g2_xor2_1 _11450_ (.B(_03439_),
    .A(_03438_),
    .X(_03523_));
 sg13g2_xnor2_1 _11451_ (.Y(_03524_),
    .A(_03438_),
    .B(_03439_));
 sg13g2_a21oi_1 _11452_ (.A1(_03459_),
    .A2(_03522_),
    .Y(_03525_),
    .B1(_03524_));
 sg13g2_o21ai_1 _11453_ (.B1(_03523_),
    .Y(_03526_),
    .A1(_03458_),
    .A2(_03521_));
 sg13g2_xor2_1 _11454_ (.B(_03435_),
    .A(_03296_),
    .X(_03527_));
 sg13g2_a21oi_1 _11455_ (.A1(_03440_),
    .A2(_03526_),
    .Y(_03528_),
    .B1(_03527_));
 sg13g2_a21o_1 _11456_ (.A2(_03526_),
    .A1(_03440_),
    .B1(_03527_),
    .X(_03529_));
 sg13g2_nor2_1 _11457_ (.A(net1871),
    .B(net1849),
    .Y(_03530_));
 sg13g2_nand2_1 _11458_ (.Y(_03531_),
    .A(net1865),
    .B(net1844));
 sg13g2_mux2_1 _11459_ (.A0(_03450_),
    .A1(_03396_),
    .S(net1883),
    .X(_03532_));
 sg13g2_nand2_1 _11460_ (.Y(_03533_),
    .A(net1903),
    .B(_03532_));
 sg13g2_nand2_1 _11461_ (.Y(_03534_),
    .A(net1916),
    .B(_03533_));
 sg13g2_nor2_1 _11462_ (.A(_03391_),
    .B(net1882),
    .Y(_03535_));
 sg13g2_a21oi_1 _11463_ (.A1(_03385_),
    .A2(net1882),
    .Y(_03536_),
    .B1(_03535_));
 sg13g2_nand2_1 _11464_ (.Y(_03537_),
    .A(_03393_),
    .B(net1882));
 sg13g2_o21ai_1 _11465_ (.B1(_03537_),
    .Y(_03538_),
    .A1(_03401_),
    .A2(net1883));
 sg13g2_mux2_1 _11466_ (.A0(_03536_),
    .A1(_03538_),
    .S(net1898),
    .X(_03539_));
 sg13g2_o21ai_1 _11467_ (.B1(_03534_),
    .Y(_03540_),
    .A1(net1916),
    .A2(_03539_));
 sg13g2_nand2_1 _11468_ (.Y(_03541_),
    .A(_03427_),
    .B(_03540_));
 sg13g2_nor2_1 _11469_ (.A(_03378_),
    .B(net1880),
    .Y(_03542_));
 sg13g2_a21oi_1 _11470_ (.A1(_03373_),
    .A2(net1879),
    .Y(_03543_),
    .B1(_03542_));
 sg13g2_nand2_1 _11471_ (.Y(_03544_),
    .A(_03380_),
    .B(net1880));
 sg13g2_o21ai_1 _11472_ (.B1(_03544_),
    .Y(_03545_),
    .A1(_03388_),
    .A2(net1880));
 sg13g2_mux2_1 _11473_ (.A0(_03543_),
    .A1(_03545_),
    .S(net1898),
    .X(_03546_));
 sg13g2_nor2_1 _11474_ (.A(_03364_),
    .B(net1879),
    .Y(_03547_));
 sg13g2_a21oi_1 _11475_ (.A1(_03358_),
    .A2(net1879),
    .Y(_03548_),
    .B1(_03547_));
 sg13g2_nand2_1 _11476_ (.Y(_03549_),
    .A(_03366_),
    .B(net1883));
 sg13g2_o21ai_1 _11477_ (.B1(_03549_),
    .Y(_03550_),
    .A1(_03370_),
    .A2(net1883));
 sg13g2_mux2_1 _11478_ (.A0(_03548_),
    .A1(_03550_),
    .S(net1897),
    .X(_03551_));
 sg13g2_mux2_1 _11479_ (.A0(_03551_),
    .A1(_03546_),
    .S(net1915),
    .X(_03552_));
 sg13g2_o21ai_1 _11480_ (.B1(_03541_),
    .Y(_03553_),
    .A1(_03424_),
    .A2(_03552_));
 sg13g2_nor2_1 _11481_ (.A(net1924),
    .B(_03331_),
    .Y(_03554_));
 sg13g2_nor2_1 _11482_ (.A(_03354_),
    .B(net1878),
    .Y(_03555_));
 sg13g2_a21oi_1 _11483_ (.A1(_03344_),
    .A2(net1878),
    .Y(_03556_),
    .B1(_03555_));
 sg13g2_nand2_1 _11484_ (.Y(_03557_),
    .A(_03352_),
    .B(net1878));
 sg13g2_o21ai_1 _11485_ (.B1(_03557_),
    .Y(_03558_),
    .A1(_03361_),
    .A2(net1878));
 sg13g2_mux2_1 _11486_ (.A0(_03556_),
    .A1(_03558_),
    .S(net1897),
    .X(_03559_));
 sg13g2_nand2_1 _11487_ (.Y(_03560_),
    .A(net1918),
    .B(_03559_));
 sg13g2_nand2_1 _11488_ (.Y(_03561_),
    .A(_03335_),
    .B(net1878));
 sg13g2_o21ai_1 _11489_ (.B1(_03561_),
    .Y(_03562_),
    .A1(_03347_),
    .A2(net1878));
 sg13g2_a21oi_2 _11490_ (.B1(net1930),
    .Y(_03563_),
    .A2(_03413_),
    .A1(_03411_));
 sg13g2_nand2_2 _11491_ (.Y(_03564_),
    .A(net1924),
    .B(_03421_));
 sg13g2_a221oi_1 _11492_ (.B2(net1897),
    .C1(_03564_),
    .B1(_03562_),
    .A1(_03328_),
    .Y(_03565_),
    .A2(_03507_));
 sg13g2_a221oi_1 _11493_ (.B2(_03565_),
    .C1(_03554_),
    .B1(_03560_),
    .A1(net1924),
    .Y(_03566_),
    .A2(_03553_));
 sg13g2_and2_1 _11494_ (.A(net1831),
    .B(_03566_),
    .X(_03567_));
 sg13g2_nand2_1 _11495_ (.Y(_03568_),
    .A(_03237_),
    .B(net1888));
 sg13g2_o21ai_1 _11496_ (.B1(_03568_),
    .Y(_03569_),
    .A1(_03229_),
    .A2(net1890));
 sg13g2_mux2_1 _11497_ (.A0(_03235_),
    .A1(_03243_),
    .S(net1889),
    .X(_03570_));
 sg13g2_mux2_1 _11498_ (.A0(_03569_),
    .A1(_03570_),
    .S(net1912),
    .X(_03571_));
 sg13g2_nand2_1 _11499_ (.Y(_03572_),
    .A(_03223_),
    .B(net1886));
 sg13g2_o21ai_1 _11500_ (.B1(_03572_),
    .Y(_03573_),
    .A1(_03217_),
    .A2(net1887));
 sg13g2_mux2_1 _11501_ (.A0(_03225_),
    .A1(_03231_),
    .S(net1887),
    .X(_03574_));
 sg13g2_mux2_1 _11502_ (.A0(_03573_),
    .A1(_03574_),
    .S(net1910),
    .X(_03575_));
 sg13g2_mux2_1 _11503_ (.A0(_03571_),
    .A1(_03575_),
    .S(net1907),
    .X(_03576_));
 sg13g2_nand2_1 _11504_ (.Y(_03577_),
    .A(net1920),
    .B(_03576_));
 sg13g2_nand2_1 _11505_ (.Y(_03578_),
    .A(_03442_),
    .B(net1889));
 sg13g2_o21ai_1 _11506_ (.B1(_03578_),
    .Y(_03579_),
    .A1(_03254_),
    .A2(net1889));
 sg13g2_nand2b_1 _11507_ (.Y(_03580_),
    .B(_03579_),
    .A_N(net1912));
 sg13g2_nand2_1 _11508_ (.Y(_03581_),
    .A(net1922),
    .B(_03580_));
 sg13g2_nand2_1 _11509_ (.Y(_03582_),
    .A(_03247_),
    .B(net1890));
 sg13g2_o21ai_1 _11510_ (.B1(_03582_),
    .Y(_03583_),
    .A1(_03241_),
    .A2(net1889));
 sg13g2_mux2_1 _11511_ (.A0(_03251_),
    .A1(_03258_),
    .S(net1890),
    .X(_03584_));
 sg13g2_mux2_1 _11512_ (.A0(_03583_),
    .A1(_03584_),
    .S(net1912),
    .X(_03585_));
 sg13g2_o21ai_1 _11513_ (.B1(_03581_),
    .Y(_03586_),
    .A1(net1922),
    .A2(_03585_));
 sg13g2_inv_1 _11514_ (.Y(_03587_),
    .A(_03586_));
 sg13g2_mux2_1 _11515_ (.A0(_03211_),
    .A1(_03219_),
    .S(net1885),
    .X(_03588_));
 sg13g2_nand2_1 _11516_ (.Y(_03589_),
    .A(_03213_),
    .B(net1885));
 sg13g2_o21ai_1 _11517_ (.B1(_03589_),
    .Y(_03590_),
    .A1(_03204_),
    .A2(net1885));
 sg13g2_mux2_1 _11518_ (.A0(_03590_),
    .A1(_03588_),
    .S(net1909),
    .X(_03591_));
 sg13g2_nand2_1 _11519_ (.Y(_03592_),
    .A(_03206_),
    .B(net1885));
 sg13g2_o21ai_1 _11520_ (.B1(_03592_),
    .Y(_03593_),
    .A1(_03196_),
    .A2(net1887));
 sg13g2_a22oi_1 _11521_ (.Y(_03594_),
    .B1(_03593_),
    .B2(net1910),
    .A2(_03494_),
    .A1(_03187_));
 sg13g2_a21oi_1 _11522_ (.A1(net1906),
    .A2(_03594_),
    .Y(_03595_),
    .B1(_03283_));
 sg13g2_o21ai_1 _11523_ (.B1(_03595_),
    .Y(_03596_),
    .A1(net1906),
    .A2(_03591_));
 sg13g2_o21ai_1 _11524_ (.B1(_03596_),
    .Y(_03597_),
    .A1(_03288_),
    .A2(_03586_));
 sg13g2_nor2_1 _11525_ (.A(net1935),
    .B(_03597_),
    .Y(_03598_));
 sg13g2_a22oi_1 _11526_ (.Y(_03599_),
    .B1(_03577_),
    .B2(_03598_),
    .A2(_03191_),
    .A1(net1934));
 sg13g2_a21oi_2 _11527_ (.B1(_03567_),
    .Y(_03600_),
    .A2(_03599_),
    .A1(net1839));
 sg13g2_a21oi_1 _11528_ (.A1(_03473_),
    .A2(_03517_),
    .Y(_03601_),
    .B1(_03468_));
 sg13g2_or2_1 _11529_ (.X(_03602_),
    .B(_03601_),
    .A(_03518_));
 sg13g2_nor2_1 _11530_ (.A(net1840),
    .B(_03602_),
    .Y(_03603_));
 sg13g2_or2_1 _11531_ (.X(_03604_),
    .B(_03510_),
    .A(_03496_));
 sg13g2_inv_1 _11532_ (.Y(_03605_),
    .A(_03604_));
 sg13g2_a21oi_1 _11533_ (.A1(_03483_),
    .A2(_03605_),
    .Y(_03606_),
    .B1(_03482_));
 sg13g2_a21oi_1 _11534_ (.A1(_03479_),
    .A2(_03606_),
    .Y(_03607_),
    .B1(_03478_));
 sg13g2_a21oi_1 _11535_ (.A1(_03473_),
    .A2(_03607_),
    .Y(_03608_),
    .B1(_03472_));
 sg13g2_xor2_1 _11536_ (.B(_03608_),
    .A(_03468_),
    .X(_03609_));
 sg13g2_a21oi_2 _11537_ (.B1(_03603_),
    .Y(_03610_),
    .A2(_03609_),
    .A1(net1841));
 sg13g2_nand3_1 _11538_ (.B(_03526_),
    .C(_03527_),
    .A(_03440_),
    .Y(_03611_));
 sg13g2_nor3_1 _11539_ (.A(_03458_),
    .B(_03521_),
    .C(_03523_),
    .Y(_03612_));
 sg13g2_nor2_1 _11540_ (.A(_03463_),
    .B(_03464_),
    .Y(_03613_));
 sg13g2_xnor2_1 _11541_ (.Y(_03614_),
    .A(_03519_),
    .B(_03613_));
 sg13g2_o21ai_1 _11542_ (.B1(_03460_),
    .Y(_03615_),
    .A1(_03464_),
    .A2(_03520_));
 sg13g2_a21oi_1 _11543_ (.A1(_03522_),
    .A2(_03615_),
    .Y(_03616_),
    .B1(_03614_));
 sg13g2_o21ai_1 _11544_ (.B1(_03616_),
    .Y(_03617_),
    .A1(_03525_),
    .A2(_03612_));
 sg13g2_nor2b_1 _11545_ (.A(_03472_),
    .B_N(_03473_),
    .Y(_03618_));
 sg13g2_xor2_1 _11546_ (.B(_03618_),
    .A(_03516_),
    .X(_03619_));
 sg13g2_or3_1 _11547_ (.A(_03479_),
    .B(_03482_),
    .C(_03514_),
    .X(_03620_));
 sg13g2_and2_1 _11548_ (.A(_03515_),
    .B(_03620_),
    .X(_03621_));
 sg13g2_and2_1 _11549_ (.A(_03511_),
    .B(_03604_),
    .X(_03622_));
 sg13g2_nand2_1 _11550_ (.Y(_03623_),
    .A(_03511_),
    .B(_03604_));
 sg13g2_nor4_1 _11551_ (.A(_03513_),
    .B(_03619_),
    .C(_03621_),
    .D(net1877),
    .Y(_03624_));
 sg13g2_nand2_1 _11552_ (.Y(_03625_),
    .A(_03602_),
    .B(_03624_));
 sg13g2_nand4_1 _11553_ (.B(_03614_),
    .C(_03615_),
    .A(_03522_),
    .Y(_03626_),
    .D(_03625_));
 sg13g2_nor3_1 _11554_ (.A(_03525_),
    .B(_03612_),
    .C(_03626_),
    .Y(_03627_));
 sg13g2_and3_2 _11555_ (.X(_03628_),
    .A(net1846),
    .B(_03611_),
    .C(_03627_));
 sg13g2_a21oi_2 _11556_ (.B1(_03617_),
    .Y(_03629_),
    .A2(_03611_),
    .A1(net1845));
 sg13g2_nor2_2 _11557_ (.A(_03628_),
    .B(_03629_),
    .Y(_03630_));
 sg13g2_xor2_1 _11558_ (.B(_03606_),
    .A(_03479_),
    .X(_03631_));
 sg13g2_mux2_1 _11559_ (.A0(_03621_),
    .A1(_03631_),
    .S(net1840),
    .X(_03632_));
 sg13g2_nor2_2 _11560_ (.A(_03630_),
    .B(_03632_),
    .Y(_03633_));
 sg13g2_or2_1 _11561_ (.X(_03634_),
    .B(_03632_),
    .A(_03630_));
 sg13g2_xnor2_1 _11562_ (.Y(_03635_),
    .A(_03607_),
    .B(_03618_));
 sg13g2_mux2_1 _11563_ (.A0(_03619_),
    .A1(_03635_),
    .S(net1840),
    .X(_03636_));
 sg13g2_nor2_2 _11564_ (.A(_03630_),
    .B(_03636_),
    .Y(_03637_));
 sg13g2_inv_4 _11565_ (.A(net1800),
    .Y(_03638_));
 sg13g2_nor3_2 _11566_ (.A(_03630_),
    .B(_03632_),
    .C(_03636_),
    .Y(_03639_));
 sg13g2_nand2_1 _11567_ (.Y(_03640_),
    .A(net1803),
    .B(net1799));
 sg13g2_o21ai_1 _11568_ (.B1(_03610_),
    .Y(_03641_),
    .A1(_03628_),
    .A2(_03629_));
 sg13g2_inv_4 _11569_ (.A(net1779),
    .Y(_03642_));
 sg13g2_nor2_2 _11570_ (.A(_03636_),
    .B(net1779),
    .Y(_03643_));
 sg13g2_nand2_2 _11571_ (.Y(_03644_),
    .A(_03610_),
    .B(net1799));
 sg13g2_nand2_2 _11572_ (.Y(_03645_),
    .A(_03610_),
    .B(_03639_));
 sg13g2_o21ai_1 _11573_ (.B1(_03511_),
    .Y(_03646_),
    .A1(net1870),
    .A2(net1848));
 sg13g2_nand3_1 _11574_ (.B(net1845),
    .C(_03604_),
    .A(net1866),
    .Y(_03647_));
 sg13g2_a21oi_1 _11575_ (.A1(_03646_),
    .A2(_03647_),
    .Y(_03648_),
    .B1(_03512_));
 sg13g2_and3_1 _11576_ (.X(_03649_),
    .A(_03512_),
    .B(_03646_),
    .C(_03647_));
 sg13g2_or2_1 _11577_ (.X(_03650_),
    .B(_03649_),
    .A(_03648_));
 sg13g2_nor3_1 _11578_ (.A(_03630_),
    .B(_03648_),
    .C(_03649_),
    .Y(_03651_));
 sg13g2_o21ai_1 _11579_ (.B1(_03622_),
    .Y(_03652_),
    .A1(_03628_),
    .A2(_03629_));
 sg13g2_and3_1 _11580_ (.X(_03653_),
    .A(net1866),
    .B(_03453_),
    .C(net1846));
 sg13g2_a21o_2 _11581_ (.A2(net1831),
    .A1(_03445_),
    .B1(_03653_),
    .X(_03654_));
 sg13g2_and3_1 _11582_ (.X(_03655_),
    .A(net1866),
    .B(net1845),
    .C(_03566_));
 sg13g2_a21oi_1 _11583_ (.A1(net1833),
    .A2(_03599_),
    .Y(_03656_),
    .B1(_03655_));
 sg13g2_a21o_1 _11584_ (.A2(_03599_),
    .A1(net1833),
    .B1(_03655_),
    .X(_03657_));
 sg13g2_mux2_1 _11585_ (.A0(_03657_),
    .A1(_03654_),
    .S(net1822),
    .X(_03658_));
 sg13g2_and2_1 _11586_ (.A(net1797),
    .B(_03658_),
    .X(_03659_));
 sg13g2_nand2_1 _11587_ (.Y(_03660_),
    .A(net1797),
    .B(_03658_));
 sg13g2_nand2_1 _11588_ (.Y(_03661_),
    .A(_03639_),
    .B(_03659_));
 sg13g2_nor2_1 _11589_ (.A(_03645_),
    .B(_03660_),
    .Y(_03662_));
 sg13g2_xnor2_1 _11590_ (.Y(_03663_),
    .A(net1947),
    .B(_03662_));
 sg13g2_nand2_1 _11591_ (.Y(_03664_),
    .A(net1932),
    .B(_03378_));
 sg13g2_mux2_1 _11592_ (.A0(_03532_),
    .A1(_03538_),
    .S(net1903),
    .X(_03665_));
 sg13g2_mux2_1 _11593_ (.A0(_03536_),
    .A1(_03545_),
    .S(net1903),
    .X(_03666_));
 sg13g2_mux2_1 _11594_ (.A0(_03666_),
    .A1(_03665_),
    .S(net1916),
    .X(_03667_));
 sg13g2_nand2_1 _11595_ (.Y(_03668_),
    .A(_03563_),
    .B(_03667_));
 sg13g2_and2_1 _11596_ (.A(_03664_),
    .B(_03668_),
    .X(_03669_));
 sg13g2_nor2_1 _11597_ (.A(net1837),
    .B(_03669_),
    .Y(_03670_));
 sg13g2_nor2_2 _11598_ (.A(net1937),
    .B(_03283_),
    .Y(_03671_));
 sg13g2_nand2b_1 _11599_ (.Y(_03672_),
    .B(net1927),
    .A_N(_03283_));
 sg13g2_mux2_1 _11600_ (.A0(_03584_),
    .A1(_03579_),
    .S(net1912),
    .X(_03673_));
 sg13g2_mux2_1 _11601_ (.A0(_03570_),
    .A1(_03583_),
    .S(net1912),
    .X(_03674_));
 sg13g2_mux2_1 _11602_ (.A0(_03673_),
    .A1(_03674_),
    .S(net1907),
    .X(_03675_));
 sg13g2_a22oi_1 _11603_ (.Y(_03676_),
    .B1(_03671_),
    .B2(_03675_),
    .A2(_03237_),
    .A1(net1936));
 sg13g2_inv_2 _11604_ (.Y(_03677_),
    .A(_03676_));
 sg13g2_a21oi_2 _11605_ (.B1(_03670_),
    .Y(_03678_),
    .A2(_03677_),
    .A1(net1837));
 sg13g2_nor2b_2 _11606_ (.A(net1778),
    .B_N(_03636_),
    .Y(_03679_));
 sg13g2_inv_1 _11607_ (.Y(_03680_),
    .A(_03679_));
 sg13g2_nand2_1 _11608_ (.Y(_03681_),
    .A(_03450_),
    .B(net1882));
 sg13g2_nor2_1 _11609_ (.A(net1897),
    .B(_03681_),
    .Y(_03682_));
 sg13g2_mux2_1 _11610_ (.A0(_03393_),
    .A1(_03391_),
    .S(net1882),
    .X(_03683_));
 sg13g2_nor2_1 _11611_ (.A(_03396_),
    .B(net1882),
    .Y(_03684_));
 sg13g2_a21oi_1 _11612_ (.A1(_03401_),
    .A2(net1882),
    .Y(_03685_),
    .B1(_03684_));
 sg13g2_mux2_1 _11613_ (.A0(_03683_),
    .A1(_03685_),
    .S(net1898),
    .X(_03686_));
 sg13g2_mux2_1 _11614_ (.A0(_03686_),
    .A1(_03682_),
    .S(net1916),
    .X(_03687_));
 sg13g2_mux2_1 _11615_ (.A0(_03380_),
    .A1(_03378_),
    .S(net1880),
    .X(_03688_));
 sg13g2_nor2_1 _11616_ (.A(_03384_),
    .B(net1882),
    .Y(_03689_));
 sg13g2_a21oi_1 _11617_ (.A1(_03388_),
    .A2(net1883),
    .Y(_03690_),
    .B1(_03689_));
 sg13g2_mux2_1 _11618_ (.A0(_03688_),
    .A1(_03690_),
    .S(net1898),
    .X(_03691_));
 sg13g2_mux2_1 _11619_ (.A0(_03366_),
    .A1(_03364_),
    .S(net1879),
    .X(_03692_));
 sg13g2_nor2_1 _11620_ (.A(_03372_),
    .B(net1879),
    .Y(_03693_));
 sg13g2_a21oi_1 _11621_ (.A1(_03370_),
    .A2(net1879),
    .Y(_03694_),
    .B1(_03693_));
 sg13g2_mux2_1 _11622_ (.A0(_03692_),
    .A1(_03694_),
    .S(net1898),
    .X(_03695_));
 sg13g2_mux2_1 _11623_ (.A0(_03695_),
    .A1(_03691_),
    .S(net1915),
    .X(_03696_));
 sg13g2_mux2_1 _11624_ (.A0(_03352_),
    .A1(_03354_),
    .S(net1878),
    .X(_03697_));
 sg13g2_nor2_1 _11625_ (.A(_03357_),
    .B(net1879),
    .Y(_03698_));
 sg13g2_a21oi_1 _11626_ (.A1(_03361_),
    .A2(net1879),
    .Y(_03699_),
    .B1(_03698_));
 sg13g2_mux2_1 _11627_ (.A0(_03697_),
    .A1(_03699_),
    .S(net1897),
    .X(_03700_));
 sg13g2_nand2_1 _11628_ (.Y(_03701_),
    .A(net1918),
    .B(_03700_));
 sg13g2_nor2_1 _11629_ (.A(_03343_),
    .B(net1881),
    .Y(_03702_));
 sg13g2_a21oi_1 _11630_ (.A1(_03347_),
    .A2(net1878),
    .Y(_03703_),
    .B1(_03702_));
 sg13g2_mux2_1 _11631_ (.A0(_03335_),
    .A1(_03337_),
    .S(net1884),
    .X(_03704_));
 sg13g2_nand2_1 _11632_ (.Y(_03705_),
    .A(net1902),
    .B(_03704_));
 sg13g2_nand2_1 _11633_ (.Y(_03706_),
    .A(net1897),
    .B(_03703_));
 sg13g2_and4_1 _11634_ (.A(net1924),
    .B(_03701_),
    .C(_03705_),
    .D(_03706_),
    .X(_03707_));
 sg13g2_a22oi_1 _11635_ (.Y(_03708_),
    .B1(_03696_),
    .B2(net1914),
    .A2(_03687_),
    .A1(_03427_));
 sg13g2_a22oi_1 _11636_ (.Y(_03709_),
    .B1(_03707_),
    .B2(_03708_),
    .A2(_03329_),
    .A1(net1928));
 sg13g2_inv_1 _11637_ (.Y(_03710_),
    .A(_03709_));
 sg13g2_nor3_1 _11638_ (.A(net1870),
    .B(net1848),
    .C(_03710_),
    .Y(_03711_));
 sg13g2_mux2_1 _11639_ (.A0(_03223_),
    .A1(_03225_),
    .S(net1886),
    .X(_03712_));
 sg13g2_nand2_1 _11640_ (.Y(_03713_),
    .A(_03228_),
    .B(net1888));
 sg13g2_o21ai_1 _11641_ (.B1(_03713_),
    .Y(_03714_),
    .A1(_03232_),
    .A2(net1888));
 sg13g2_mux2_1 _11642_ (.A0(_03712_),
    .A1(_03714_),
    .S(net1911),
    .X(_03715_));
 sg13g2_and2_1 _11643_ (.A(net1907),
    .B(_03715_),
    .X(_03716_));
 sg13g2_mux2_1 _11644_ (.A0(_03237_),
    .A1(_03235_),
    .S(net1888),
    .X(_03717_));
 sg13g2_nand2_1 _11645_ (.Y(_03718_),
    .A(_03240_),
    .B(net1888));
 sg13g2_o21ai_1 _11646_ (.B1(_03718_),
    .Y(_03719_),
    .A1(_03244_),
    .A2(net1888));
 sg13g2_mux2_1 _11647_ (.A0(_03717_),
    .A1(_03719_),
    .S(net1911),
    .X(_03720_));
 sg13g2_a21oi_1 _11648_ (.A1(net1923),
    .A2(_03720_),
    .Y(_03721_),
    .B1(_03716_));
 sg13g2_nand2b_1 _11649_ (.Y(_03722_),
    .B(_03442_),
    .A_N(net1889));
 sg13g2_nor2_1 _11650_ (.A(net1912),
    .B(_03722_),
    .Y(_03723_));
 sg13g2_mux2_1 _11651_ (.A0(_03247_),
    .A1(_03251_),
    .S(net1889),
    .X(_03724_));
 sg13g2_nand2_1 _11652_ (.Y(_03725_),
    .A(_03255_),
    .B(net1888));
 sg13g2_o21ai_1 _11653_ (.B1(_03725_),
    .Y(_03726_),
    .A1(_03259_),
    .A2(net1889));
 sg13g2_mux2_1 _11654_ (.A0(_03724_),
    .A1(_03726_),
    .S(net1912),
    .X(_03727_));
 sg13g2_mux2_1 _11655_ (.A0(_03723_),
    .A1(_03727_),
    .S(net1908),
    .X(_03728_));
 sg13g2_nand2b_1 _11656_ (.Y(_03729_),
    .B(_03728_),
    .A_N(_03288_));
 sg13g2_nand2_1 _11657_ (.Y(_03730_),
    .A(_03216_),
    .B(net1886));
 sg13g2_o21ai_1 _11658_ (.B1(_03730_),
    .Y(_03731_),
    .A1(_03220_),
    .A2(net1886));
 sg13g2_mux2_1 _11659_ (.A0(_03213_),
    .A1(_03211_),
    .S(net1885),
    .X(_03732_));
 sg13g2_mux2_1 _11660_ (.A0(_03732_),
    .A1(_03731_),
    .S(net1909),
    .X(_03733_));
 sg13g2_nand2_1 _11661_ (.Y(_03734_),
    .A(_03204_),
    .B(net1885));
 sg13g2_o21ai_1 _11662_ (.B1(_03734_),
    .Y(_03735_),
    .A1(_03206_),
    .A2(net1885));
 sg13g2_nand2_1 _11663_ (.Y(_03736_),
    .A(_03195_),
    .B(net1885));
 sg13g2_a21oi_1 _11664_ (.A1(_03198_),
    .A2(_03484_),
    .Y(_03737_),
    .B1(net1909));
 sg13g2_a22oi_1 _11665_ (.Y(_03738_),
    .B1(_03736_),
    .B2(_03737_),
    .A2(_03735_),
    .A1(net1909));
 sg13g2_inv_1 _11666_ (.Y(_03739_),
    .A(_03738_));
 sg13g2_a21oi_1 _11667_ (.A1(net1923),
    .A2(_03733_),
    .Y(_03740_),
    .B1(net1919));
 sg13g2_a22oi_1 _11668_ (.Y(_03741_),
    .B1(_03739_),
    .B2(_03740_),
    .A2(_03721_),
    .A1(net1919));
 sg13g2_nor2_1 _11669_ (.A(net1934),
    .B(_03741_),
    .Y(_03742_));
 sg13g2_a22oi_1 _11670_ (.Y(_03743_),
    .B1(_03729_),
    .B2(_03742_),
    .A2(_03188_),
    .A1(net1934));
 sg13g2_a21oi_1 _11671_ (.A1(net1832),
    .A2(_03743_),
    .Y(_03744_),
    .B1(_03711_));
 sg13g2_a21o_1 _11672_ (.A2(_03743_),
    .A1(net1832),
    .B1(_03711_),
    .X(_03745_));
 sg13g2_and2_1 _11673_ (.A(_03419_),
    .B(_03665_),
    .X(_03746_));
 sg13g2_nor2_1 _11674_ (.A(_03428_),
    .B(_03746_),
    .Y(_03747_));
 sg13g2_mux2_1 _11675_ (.A0(_03543_),
    .A1(_03550_),
    .S(net1902),
    .X(_03748_));
 sg13g2_mux2_1 _11676_ (.A0(_03748_),
    .A1(_03666_),
    .S(net1917),
    .X(_03749_));
 sg13g2_mux2_1 _11677_ (.A0(_03548_),
    .A1(_03558_),
    .S(net1902),
    .X(_03750_));
 sg13g2_inv_1 _11678_ (.Y(_03751_),
    .A(_03750_));
 sg13g2_nand2_1 _11679_ (.Y(_03752_),
    .A(net1897),
    .B(_03556_));
 sg13g2_a21oi_1 _11680_ (.A1(net1902),
    .A2(_03562_),
    .Y(_03753_),
    .B1(net1918));
 sg13g2_nand2_1 _11681_ (.Y(_03754_),
    .A(_03752_),
    .B(_03753_));
 sg13g2_a21oi_1 _11682_ (.A1(net1915),
    .A2(_03751_),
    .Y(_03755_),
    .B1(net1913));
 sg13g2_a221oi_1 _11683_ (.B2(_03755_),
    .C1(_03427_),
    .B1(_03754_),
    .A1(net1913),
    .Y(_03756_),
    .A2(_03749_));
 sg13g2_nor2_1 _11684_ (.A(_03747_),
    .B(_03756_),
    .Y(_03757_));
 sg13g2_a21oi_2 _11685_ (.B1(_03757_),
    .Y(_03758_),
    .A2(_03337_),
    .A1(net1928));
 sg13g2_nor3_1 _11686_ (.A(net1870),
    .B(net1848),
    .C(_03758_),
    .Y(_03759_));
 sg13g2_mux2_1 _11687_ (.A0(_03574_),
    .A1(_03569_),
    .S(net1911),
    .X(_03760_));
 sg13g2_mux2_1 _11688_ (.A0(_03674_),
    .A1(_03760_),
    .S(net1906),
    .X(_03761_));
 sg13g2_nand2_1 _11689_ (.Y(_03762_),
    .A(net1907),
    .B(_03673_));
 sg13g2_inv_1 _11690_ (.Y(_03763_),
    .A(_03762_));
 sg13g2_mux2_1 _11691_ (.A0(_03588_),
    .A1(_03573_),
    .S(net1909),
    .X(_03764_));
 sg13g2_mux2_1 _11692_ (.A0(_03593_),
    .A1(_03590_),
    .S(net1909),
    .X(_03765_));
 sg13g2_o21ai_1 _11693_ (.B1(net1904),
    .Y(_03766_),
    .A1(net1934),
    .A2(_03763_));
 sg13g2_a221oi_1 _11694_ (.B2(net1923),
    .C1(_03765_),
    .B1(_03764_),
    .A1(net1919),
    .Y(_03767_),
    .A2(_03761_));
 sg13g2_a22oi_1 _11695_ (.Y(_03768_),
    .B1(_03766_),
    .B2(_03767_),
    .A2(_03199_),
    .A1(net1934));
 sg13g2_a21oi_1 _11696_ (.A1(net1832),
    .A2(_03768_),
    .Y(_03769_),
    .B1(_03759_));
 sg13g2_a21o_1 _11697_ (.A2(_03768_),
    .A1(net1832),
    .B1(_03759_),
    .X(_03770_));
 sg13g2_mux2_1 _11698_ (.A0(_03770_),
    .A1(_03745_),
    .S(net1821),
    .X(_03771_));
 sg13g2_mux2_1 _11699_ (.A0(_03658_),
    .A1(_03771_),
    .S(net1797),
    .X(_03772_));
 sg13g2_nand2_1 _11700_ (.Y(_03773_),
    .A(net1928),
    .B(_03335_));
 sg13g2_nand2_1 _11701_ (.Y(_03774_),
    .A(net1897),
    .B(_03697_));
 sg13g2_nand2_1 _11702_ (.Y(_03775_),
    .A(net1902),
    .B(_03703_));
 sg13g2_mux2_1 _11703_ (.A0(_03692_),
    .A1(_03699_),
    .S(net1902),
    .X(_03776_));
 sg13g2_a21o_1 _11704_ (.A2(_03775_),
    .A1(_03774_),
    .B1(net1918),
    .X(_03777_));
 sg13g2_nand2_1 _11705_ (.Y(_03778_),
    .A(net1915),
    .B(_03776_));
 sg13g2_nand3_1 _11706_ (.B(_03777_),
    .C(_03778_),
    .A(_03421_),
    .Y(_03779_));
 sg13g2_nor2_1 _11707_ (.A(net1903),
    .B(_03681_),
    .Y(_03780_));
 sg13g2_a21oi_1 _11708_ (.A1(net1903),
    .A2(_03685_),
    .Y(_03781_),
    .B1(_03780_));
 sg13g2_nor2b_1 _11709_ (.A(_03781_),
    .B_N(_03419_),
    .Y(_03782_));
 sg13g2_nor2_1 _11710_ (.A(_03428_),
    .B(_03782_),
    .Y(_03783_));
 sg13g2_mux2_1 _11711_ (.A0(_03688_),
    .A1(_03694_),
    .S(net1902),
    .X(_03784_));
 sg13g2_mux2_1 _11712_ (.A0(_03683_),
    .A1(_03690_),
    .S(net1903),
    .X(_03785_));
 sg13g2_mux2_1 _11713_ (.A0(_03784_),
    .A1(_03785_),
    .S(net1915),
    .X(_03786_));
 sg13g2_o21ai_1 _11714_ (.B1(_03779_),
    .Y(_03787_),
    .A1(_03424_),
    .A2(_03786_));
 sg13g2_o21ai_1 _11715_ (.B1(_03773_),
    .Y(_03788_),
    .A1(_03783_),
    .A2(_03787_));
 sg13g2_and3_1 _11716_ (.X(_03789_),
    .A(net1866),
    .B(net1845),
    .C(_03788_));
 sg13g2_nand2_1 _11717_ (.Y(_03790_),
    .A(net1912),
    .B(_03722_));
 sg13g2_o21ai_1 _11718_ (.B1(_03790_),
    .Y(_03791_),
    .A1(_03266_),
    .A2(_03726_));
 sg13g2_nor2_1 _11719_ (.A(net1922),
    .B(_03791_),
    .Y(_03792_));
 sg13g2_o21ai_1 _11720_ (.B1(net1927),
    .Y(_03793_),
    .A1(net1922),
    .A2(_03791_));
 sg13g2_nand2_1 _11721_ (.Y(_03794_),
    .A(net1904),
    .B(_03793_));
 sg13g2_mux2_1 _11722_ (.A0(_03719_),
    .A1(_03724_),
    .S(net1911),
    .X(_03795_));
 sg13g2_mux2_1 _11723_ (.A0(_03714_),
    .A1(_03717_),
    .S(net1911),
    .X(_03796_));
 sg13g2_mux2_1 _11724_ (.A0(_03795_),
    .A1(_03796_),
    .S(net1907),
    .X(_03797_));
 sg13g2_mux2_1 _11725_ (.A0(_03731_),
    .A1(_03712_),
    .S(net1910),
    .X(_03798_));
 sg13g2_or2_1 _11726_ (.X(_03799_),
    .B(_03798_),
    .A(net1906));
 sg13g2_nand2_1 _11727_ (.Y(_03800_),
    .A(net1909),
    .B(_03732_));
 sg13g2_o21ai_1 _11728_ (.B1(_03800_),
    .Y(_03801_),
    .A1(net1909),
    .A2(_03735_));
 sg13g2_a22oi_1 _11729_ (.Y(_03802_),
    .B1(_03799_),
    .B2(_03801_),
    .A2(_03797_),
    .A1(net1919));
 sg13g2_a22oi_1 _11730_ (.Y(_03803_),
    .B1(_03794_),
    .B2(_03802_),
    .A2(_03196_),
    .A1(net1934));
 sg13g2_a21oi_1 _11731_ (.A1(net1832),
    .A2(_03803_),
    .Y(_03804_),
    .B1(_03789_));
 sg13g2_mux2_1 _11732_ (.A0(_03546_),
    .A1(_03539_),
    .S(net1917),
    .X(_03805_));
 sg13g2_nor2_1 _11733_ (.A(net1917),
    .B(_03533_),
    .Y(_03806_));
 sg13g2_mux2_1 _11734_ (.A0(_03559_),
    .A1(_03551_),
    .S(net1918),
    .X(_03807_));
 sg13g2_a221oi_1 _11735_ (.B2(_03427_),
    .C1(net1928),
    .B1(_03806_),
    .A1(net1913),
    .Y(_03808_),
    .A2(_03805_));
 sg13g2_nand2b_1 _11736_ (.Y(_03809_),
    .B(_03808_),
    .A_N(_03807_));
 sg13g2_o21ai_1 _11737_ (.B1(_03809_),
    .Y(_03810_),
    .A1(net1924),
    .A2(_03346_));
 sg13g2_inv_2 _11738_ (.Y(_03811_),
    .A(_03810_));
 sg13g2_nor3_1 _11739_ (.A(net1870),
    .B(net1848),
    .C(_03810_),
    .Y(_03812_));
 sg13g2_mux2_1 _11740_ (.A0(_03571_),
    .A1(_03585_),
    .S(_03278_),
    .X(_03813_));
 sg13g2_nor2_1 _11741_ (.A(net1922),
    .B(_03580_),
    .Y(_03814_));
 sg13g2_nand2_1 _11742_ (.Y(_03815_),
    .A(net1906),
    .B(_03591_));
 sg13g2_o21ai_1 _11743_ (.B1(net1904),
    .Y(_03816_),
    .A1(net1935),
    .A2(_03814_));
 sg13g2_nand2_1 _11744_ (.Y(_03817_),
    .A(_03815_),
    .B(_03816_));
 sg13g2_a221oi_1 _11745_ (.B2(net1919),
    .C1(_03817_),
    .B1(_03813_),
    .A1(net1922),
    .Y(_03818_),
    .A2(_03575_));
 sg13g2_a21oi_2 _11746_ (.B1(_03818_),
    .Y(_03819_),
    .A2(_03207_),
    .A1(net1934));
 sg13g2_a21oi_1 _11747_ (.A1(net1832),
    .A2(_03819_),
    .Y(_03820_),
    .B1(_03812_));
 sg13g2_mux4_1 _11748_ (.S0(net1832),
    .A0(_03811_),
    .A1(_03819_),
    .A2(_03788_),
    .A3(_03803_),
    .S1(net1821),
    .X(_03821_));
 sg13g2_mux2_1 _11749_ (.A0(_03691_),
    .A1(_03686_),
    .S(net1917),
    .X(_03822_));
 sg13g2_nand2b_2 _11750_ (.Y(_03823_),
    .B(_03682_),
    .A_N(net1916));
 sg13g2_a21oi_1 _11751_ (.A1(net1924),
    .A2(_03823_),
    .Y(_03824_),
    .B1(_03428_));
 sg13g2_mux2_1 _11752_ (.A0(_03700_),
    .A1(_03695_),
    .S(net1915),
    .X(_03825_));
 sg13g2_a21oi_1 _11753_ (.A1(net1914),
    .A2(_03822_),
    .Y(_03826_),
    .B1(_03825_));
 sg13g2_nand2b_1 _11754_ (.Y(_03827_),
    .B(_03826_),
    .A_N(_03824_));
 sg13g2_o21ai_1 _11755_ (.B1(_03827_),
    .Y(_03828_),
    .A1(net1924),
    .A2(_03343_));
 sg13g2_nor3_1 _11756_ (.A(net1869),
    .B(net1847),
    .C(_03828_),
    .Y(_03829_));
 sg13g2_mux2_1 _11757_ (.A0(_03720_),
    .A1(_03727_),
    .S(net1923),
    .X(_03830_));
 sg13g2_and2_1 _11758_ (.A(net1923),
    .B(_03715_),
    .X(_03831_));
 sg13g2_nand2_1 _11759_ (.Y(_03832_),
    .A(net1908),
    .B(_03723_));
 sg13g2_nand2_1 _11760_ (.Y(_03833_),
    .A(net1927),
    .B(_03832_));
 sg13g2_a21oi_1 _11761_ (.A1(net1906),
    .A2(_03733_),
    .Y(_03834_),
    .B1(_03831_));
 sg13g2_a22oi_1 _11762_ (.Y(_03835_),
    .B1(_03833_),
    .B2(net1904),
    .A2(_03830_),
    .A1(net1920));
 sg13g2_a22oi_1 _11763_ (.Y(_03836_),
    .B1(_03834_),
    .B2(_03835_),
    .A2(_03204_),
    .A1(net1935));
 sg13g2_a21oi_1 _11764_ (.A1(net1829),
    .A2(_03836_),
    .Y(_03837_),
    .B1(_03829_));
 sg13g2_a21o_1 _11765_ (.A2(_03836_),
    .A1(net1829),
    .B1(_03829_),
    .X(_03838_));
 sg13g2_nor2_1 _11766_ (.A(net1917),
    .B(_03751_),
    .Y(_03839_));
 sg13g2_a21oi_1 _11767_ (.A1(net1915),
    .A2(_03748_),
    .Y(_03840_),
    .B1(_03839_));
 sg13g2_o21ai_1 _11768_ (.B1(_03428_),
    .Y(_03841_),
    .A1(_03424_),
    .A2(_03667_));
 sg13g2_a21oi_1 _11769_ (.A1(_03424_),
    .A2(_03840_),
    .Y(_03842_),
    .B1(_03841_));
 sg13g2_a21o_2 _11770_ (.A2(_03354_),
    .A1(net1928),
    .B1(_03842_),
    .X(_03843_));
 sg13g2_and3_1 _11771_ (.X(_03844_),
    .A(net1863),
    .B(net1842),
    .C(_03843_));
 sg13g2_nand2_1 _11772_ (.Y(_03845_),
    .A(net1906),
    .B(_03764_));
 sg13g2_a21oi_1 _11773_ (.A1(net1923),
    .A2(_03760_),
    .Y(_03846_),
    .B1(net1919));
 sg13g2_nand2b_1 _11774_ (.Y(_03847_),
    .B(net1920),
    .A_N(_03675_));
 sg13g2_a21oi_1 _11775_ (.A1(_03845_),
    .A2(_03846_),
    .Y(_03848_),
    .B1(net1904));
 sg13g2_a22oi_1 _11776_ (.Y(_03849_),
    .B1(_03847_),
    .B2(_03848_),
    .A2(_03213_),
    .A1(net1934));
 sg13g2_inv_1 _11777_ (.Y(_03850_),
    .A(_03849_));
 sg13g2_a21oi_1 _11778_ (.A1(net1828),
    .A2(_03850_),
    .Y(_03851_),
    .B1(_03844_));
 sg13g2_a21o_1 _11779_ (.A2(_03850_),
    .A1(net1828),
    .B1(_03844_),
    .X(_03852_));
 sg13g2_mux2_1 _11780_ (.A0(_03852_),
    .A1(_03838_),
    .S(net1819),
    .X(_03853_));
 sg13g2_mux4_1 _11781_ (.S0(net1798),
    .A0(_03658_),
    .A1(_03771_),
    .A2(_03821_),
    .A3(_03853_),
    .S1(net1804),
    .X(_03854_));
 sg13g2_mux2_1 _11782_ (.A0(_03776_),
    .A1(_03784_),
    .S(net1915),
    .X(_03855_));
 sg13g2_nand2_1 _11783_ (.Y(_03856_),
    .A(net1916),
    .B(_03781_));
 sg13g2_o21ai_1 _11784_ (.B1(_03856_),
    .Y(_03857_),
    .A1(net1916),
    .A2(_03785_));
 sg13g2_a21oi_1 _11785_ (.A1(net1913),
    .A2(_03857_),
    .Y(_03858_),
    .B1(_03429_));
 sg13g2_a22oi_1 _11786_ (.Y(_03859_),
    .B1(_03855_),
    .B2(_03858_),
    .A2(_03352_),
    .A1(net1928));
 sg13g2_inv_1 _11787_ (.Y(_03860_),
    .A(_03859_));
 sg13g2_nor3_1 _11788_ (.A(net1869),
    .B(net1847),
    .C(_03859_),
    .Y(_03861_));
 sg13g2_nand2_1 _11789_ (.Y(_03862_),
    .A(net1922),
    .B(_03791_));
 sg13g2_o21ai_1 _11790_ (.B1(_03862_),
    .Y(_03863_),
    .A1(net1922),
    .A2(_03795_));
 sg13g2_nand2_1 _11791_ (.Y(_03864_),
    .A(net1923),
    .B(_03796_));
 sg13g2_a21oi_1 _11792_ (.A1(net1906),
    .A2(_03798_),
    .Y(_03865_),
    .B1(net1919));
 sg13g2_a221oi_1 _11793_ (.B2(_03865_),
    .C1(net1904),
    .B1(_03864_),
    .A1(net1919),
    .Y(_03866_),
    .A2(_03863_));
 sg13g2_a21o_2 _11794_ (.A2(_03211_),
    .A1(net1935),
    .B1(_03866_),
    .X(_03867_));
 sg13g2_a21oi_1 _11795_ (.A1(net1828),
    .A2(_03867_),
    .Y(_03868_),
    .B1(_03861_));
 sg13g2_a21o_1 _11796_ (.A2(_03867_),
    .A1(net1828),
    .B1(_03861_),
    .X(_03869_));
 sg13g2_nand2_1 _11797_ (.Y(_03870_),
    .A(net1932),
    .B(_03360_));
 sg13g2_a21oi_1 _11798_ (.A1(net1914),
    .A2(_03540_),
    .Y(_03871_),
    .B1(_03429_));
 sg13g2_o21ai_1 _11799_ (.B1(_03871_),
    .Y(_03872_),
    .A1(net1913),
    .A2(_03552_));
 sg13g2_and2_1 _11800_ (.A(_03870_),
    .B(_03872_),
    .X(_03873_));
 sg13g2_nor3_1 _11801_ (.A(net1869),
    .B(net1847),
    .C(_03873_),
    .Y(_03874_));
 sg13g2_a21oi_1 _11802_ (.A1(net1920),
    .A2(_03586_),
    .Y(_03875_),
    .B1(net1904));
 sg13g2_o21ai_1 _11803_ (.B1(_03875_),
    .Y(_03876_),
    .A1(_03283_),
    .A2(_03576_));
 sg13g2_o21ai_1 _11804_ (.B1(_03876_),
    .Y(_03877_),
    .A1(net1927),
    .A2(_03220_));
 sg13g2_a21oi_1 _11805_ (.A1(net1828),
    .A2(_03877_),
    .Y(_03878_),
    .B1(_03874_));
 sg13g2_a21o_1 _11806_ (.A2(_03877_),
    .A1(net1828),
    .B1(_03874_),
    .X(_03879_));
 sg13g2_mux2_1 _11807_ (.A0(_03878_),
    .A1(_03868_),
    .S(net1819),
    .X(_03880_));
 sg13g2_mux2_1 _11808_ (.A0(_03879_),
    .A1(_03869_),
    .S(net1819),
    .X(_03881_));
 sg13g2_nor2_1 _11809_ (.A(_03424_),
    .B(_03687_),
    .Y(_03882_));
 sg13g2_o21ai_1 _11810_ (.B1(_03428_),
    .Y(_03883_),
    .A1(net1913),
    .A2(_03696_));
 sg13g2_nor2_1 _11811_ (.A(_03882_),
    .B(_03883_),
    .Y(_03884_));
 sg13g2_a21oi_1 _11812_ (.A1(net1929),
    .A2(_03357_),
    .Y(_03885_),
    .B1(_03884_));
 sg13g2_inv_1 _11813_ (.Y(_03886_),
    .A(_03885_));
 sg13g2_nor3_1 _11814_ (.A(net1869),
    .B(net1847),
    .C(_03885_),
    .Y(_03887_));
 sg13g2_a21oi_1 _11815_ (.A1(_03285_),
    .A2(_03721_),
    .Y(_03888_),
    .B1(net1905));
 sg13g2_o21ai_1 _11816_ (.B1(_03888_),
    .Y(_03889_),
    .A1(_03285_),
    .A2(_03728_));
 sg13g2_o21ai_1 _11817_ (.B1(_03889_),
    .Y(_03890_),
    .A1(net1927),
    .A2(_03217_));
 sg13g2_a21oi_1 _11818_ (.A1(net1828),
    .A2(_03890_),
    .Y(_03891_),
    .B1(_03887_));
 sg13g2_nand2_1 _11819_ (.Y(_03892_),
    .A(net1928),
    .B(_03364_));
 sg13g2_nor2_1 _11820_ (.A(net1913),
    .B(_03749_),
    .Y(_03893_));
 sg13g2_a21oi_1 _11821_ (.A1(_03422_),
    .A2(_03746_),
    .Y(_03894_),
    .B1(_03563_));
 sg13g2_o21ai_1 _11822_ (.B1(_03892_),
    .Y(_03895_),
    .A1(_03893_),
    .A2(_03894_));
 sg13g2_inv_1 _11823_ (.Y(_03896_),
    .A(_03895_));
 sg13g2_nor3_1 _11824_ (.A(net1869),
    .B(net1847),
    .C(_03896_),
    .Y(_03897_));
 sg13g2_or2_1 _11825_ (.X(_03898_),
    .B(_03761_),
    .A(net1920));
 sg13g2_a21oi_1 _11826_ (.A1(net1920),
    .A2(_03762_),
    .Y(_03899_),
    .B1(net1904));
 sg13g2_a22oi_1 _11827_ (.Y(_03900_),
    .B1(_03898_),
    .B2(_03899_),
    .A2(_03223_),
    .A1(net1936));
 sg13g2_inv_1 _11828_ (.Y(_03901_),
    .A(_03900_));
 sg13g2_a21oi_1 _11829_ (.A1(net1829),
    .A2(_03901_),
    .Y(_03902_),
    .B1(_03897_));
 sg13g2_mux2_1 _11830_ (.A0(_03902_),
    .A1(_03891_),
    .S(net1819),
    .X(_03903_));
 sg13g2_mux4_1 _11831_ (.S0(net1829),
    .A0(_03895_),
    .A1(_03901_),
    .A2(_03886_),
    .A3(_03890_),
    .S1(net1820),
    .X(_03904_));
 sg13g2_mux2_1 _11832_ (.A0(_03880_),
    .A1(_03903_),
    .S(net1794),
    .X(_03905_));
 sg13g2_nand2b_1 _11833_ (.Y(_03906_),
    .B(net1801),
    .A_N(_03905_));
 sg13g2_nand2b_1 _11834_ (.Y(_03907_),
    .B(_03424_),
    .A_N(_03786_));
 sg13g2_a21o_1 _11835_ (.A2(_03782_),
    .A1(_03422_),
    .B1(_03563_),
    .X(_03908_));
 sg13g2_a22oi_1 _11836_ (.Y(_03909_),
    .B1(_03907_),
    .B2(_03908_),
    .A2(_03366_),
    .A1(net1929));
 sg13g2_nor3_1 _11837_ (.A(net1869),
    .B(net1847),
    .C(_03909_),
    .Y(_03910_));
 sg13g2_nor2_1 _11838_ (.A(net1921),
    .B(_03797_),
    .Y(_03911_));
 sg13g2_nor2_1 _11839_ (.A(_03285_),
    .B(_03792_),
    .Y(_03912_));
 sg13g2_nor3_1 _11840_ (.A(net1905),
    .B(_03911_),
    .C(_03912_),
    .Y(_03913_));
 sg13g2_a21oi_1 _11841_ (.A1(net1936),
    .A2(_03225_),
    .Y(_03914_),
    .B1(_03913_));
 sg13g2_inv_2 _11842_ (.Y(_03915_),
    .A(_03914_));
 sg13g2_a21oi_1 _11843_ (.A1(net1829),
    .A2(_03915_),
    .Y(_03916_),
    .B1(_03910_));
 sg13g2_nor2_1 _11844_ (.A(net1913),
    .B(_03805_),
    .Y(_03917_));
 sg13g2_o21ai_1 _11845_ (.B1(_03428_),
    .Y(_03918_),
    .A1(_03424_),
    .A2(_03806_));
 sg13g2_nor2_1 _11846_ (.A(_03917_),
    .B(_03918_),
    .Y(_03919_));
 sg13g2_a21oi_2 _11847_ (.B1(_03919_),
    .Y(_03920_),
    .A2(_03369_),
    .A1(net1929));
 sg13g2_inv_1 _11848_ (.Y(_03921_),
    .A(_03920_));
 sg13g2_nor3_1 _11849_ (.A(net1869),
    .B(net1847),
    .C(_03920_),
    .Y(_03922_));
 sg13g2_nor2_1 _11850_ (.A(net1920),
    .B(_03813_),
    .Y(_03923_));
 sg13g2_nor2_1 _11851_ (.A(_03285_),
    .B(_03814_),
    .Y(_03924_));
 sg13g2_nor3_1 _11852_ (.A(net1905),
    .B(_03923_),
    .C(_03924_),
    .Y(_03925_));
 sg13g2_a21oi_1 _11853_ (.A1(net1936),
    .A2(_03231_),
    .Y(_03926_),
    .B1(_03925_));
 sg13g2_inv_2 _11854_ (.Y(_03927_),
    .A(_03926_));
 sg13g2_a21oi_1 _11855_ (.A1(net1830),
    .A2(_03927_),
    .Y(_03928_),
    .B1(_03922_));
 sg13g2_mux2_1 _11856_ (.A0(_03928_),
    .A1(_03916_),
    .S(net1820),
    .X(_03929_));
 sg13g2_nand2_1 _11857_ (.Y(_03930_),
    .A(net1932),
    .B(_03372_));
 sg13g2_a21oi_1 _11858_ (.A1(net1914),
    .A2(_03823_),
    .Y(_03931_),
    .B1(_03429_));
 sg13g2_o21ai_1 _11859_ (.B1(_03931_),
    .Y(_03932_),
    .A1(net1914),
    .A2(_03822_));
 sg13g2_and2_1 _11860_ (.A(_03930_),
    .B(_03932_),
    .X(_03933_));
 sg13g2_nor3_2 _11861_ (.A(net1870),
    .B(net1848),
    .C(_03933_),
    .Y(_03934_));
 sg13g2_or2_1 _11862_ (.X(_03935_),
    .B(_03830_),
    .A(net1921));
 sg13g2_a21oi_1 _11863_ (.A1(net1920),
    .A2(_03832_),
    .Y(_03936_),
    .B1(net1905));
 sg13g2_a22oi_1 _11864_ (.Y(_03937_),
    .B1(_03935_),
    .B2(_03936_),
    .A2(_03228_),
    .A1(net1937));
 sg13g2_inv_2 _11865_ (.Y(_03938_),
    .A(_03937_));
 sg13g2_a21oi_2 _11866_ (.B1(_03934_),
    .Y(_03939_),
    .A2(_03938_),
    .A1(net1830));
 sg13g2_nor3_1 _11867_ (.A(net1869),
    .B(net1847),
    .C(_03669_),
    .Y(_03940_));
 sg13g2_a21oi_1 _11868_ (.A1(net1830),
    .A2(_03677_),
    .Y(_03941_),
    .B1(_03940_));
 sg13g2_mux2_1 _11869_ (.A0(_03941_),
    .A1(_03939_),
    .S(net1820),
    .X(_03942_));
 sg13g2_mux2_1 _11870_ (.A0(_03929_),
    .A1(_03942_),
    .S(net1795),
    .X(_03943_));
 sg13g2_o21ai_1 _11871_ (.B1(_03906_),
    .Y(_03944_),
    .A1(net1801),
    .A2(_03943_));
 sg13g2_a22oi_1 _11872_ (.Y(_03945_),
    .B1(_03944_),
    .B2(net1777),
    .A2(_03854_),
    .A1(_03679_));
 sg13g2_xnor2_1 _11873_ (.Y(_03946_),
    .A(net1947),
    .B(_03945_));
 sg13g2_nor2b_1 _11874_ (.A(_03678_),
    .B_N(_03946_),
    .Y(_03947_));
 sg13g2_xnor2_1 _11875_ (.Y(_03948_),
    .A(_03678_),
    .B(_03946_));
 sg13g2_nor2_1 _11876_ (.A(_03564_),
    .B(_03857_),
    .Y(_03949_));
 sg13g2_a21oi_2 _11877_ (.B1(_03949_),
    .Y(_03950_),
    .A2(_03380_),
    .A1(net1930));
 sg13g2_a21oi_1 _11878_ (.A1(net1865),
    .A2(net1843),
    .Y(_03951_),
    .B1(_03950_));
 sg13g2_nand2_1 _11879_ (.Y(_03952_),
    .A(net1936),
    .B(_03235_));
 sg13g2_o21ai_1 _11880_ (.B1(_03952_),
    .Y(_03953_),
    .A1(_03672_),
    .A2(_03863_));
 sg13g2_a21oi_2 _11881_ (.B1(_03951_),
    .Y(_03954_),
    .A2(_03953_),
    .A1(net1837));
 sg13g2_mux2_1 _11882_ (.A0(_03744_),
    .A1(_03656_),
    .S(net1822),
    .X(_03955_));
 sg13g2_mux2_1 _11883_ (.A0(_03804_),
    .A1(_03769_),
    .S(net1821),
    .X(_03956_));
 sg13g2_mux2_1 _11884_ (.A0(_03955_),
    .A1(_03956_),
    .S(net1798),
    .X(_03957_));
 sg13g2_mux2_1 _11885_ (.A0(_03837_),
    .A1(_03820_),
    .S(net1820),
    .X(_03958_));
 sg13g2_mux2_1 _11886_ (.A0(_03868_),
    .A1(_03851_),
    .S(net1819),
    .X(_03959_));
 sg13g2_mux2_1 _11887_ (.A0(_03958_),
    .A1(_03959_),
    .S(net1795),
    .X(_03960_));
 sg13g2_mux2_1 _11888_ (.A0(_03957_),
    .A1(_03960_),
    .S(net1802),
    .X(_03961_));
 sg13g2_mux2_1 _11889_ (.A0(_03891_),
    .A1(_03878_),
    .S(net1819),
    .X(_03962_));
 sg13g2_mux2_1 _11890_ (.A0(_03916_),
    .A1(_03902_),
    .S(net1819),
    .X(_03963_));
 sg13g2_mux2_1 _11891_ (.A0(_03962_),
    .A1(_03963_),
    .S(net1794),
    .X(_03964_));
 sg13g2_mux2_1 _11892_ (.A0(_03939_),
    .A1(_03928_),
    .S(net1819),
    .X(_03965_));
 sg13g2_nor3_1 _11893_ (.A(net1871),
    .B(net1849),
    .C(_03950_),
    .Y(_03966_));
 sg13g2_a21oi_1 _11894_ (.A1(net1830),
    .A2(_03953_),
    .Y(_03967_),
    .B1(_03966_));
 sg13g2_mux2_1 _11895_ (.A0(_03967_),
    .A1(_03941_),
    .S(net1820),
    .X(_03968_));
 sg13g2_mux2_1 _11896_ (.A0(_03965_),
    .A1(_03968_),
    .S(net1794),
    .X(_03969_));
 sg13g2_mux2_1 _11897_ (.A0(_03964_),
    .A1(_03969_),
    .S(net1802),
    .X(_03970_));
 sg13g2_nand2b_1 _11898_ (.Y(_03971_),
    .B(_03654_),
    .A_N(net1821));
 sg13g2_or2_1 _11899_ (.X(_03972_),
    .B(_03971_),
    .A(_03650_));
 sg13g2_inv_1 _11900_ (.Y(_03973_),
    .A(_03972_));
 sg13g2_a21oi_1 _11901_ (.A1(_03639_),
    .A2(_03973_),
    .Y(_03974_),
    .B1(_03642_));
 sg13g2_a221oi_1 _11902_ (.B2(_03643_),
    .C1(_03974_),
    .B1(_03970_),
    .A1(_03679_),
    .Y(_03975_),
    .A2(_03961_));
 sg13g2_xnor2_1 _11903_ (.Y(_03976_),
    .A(net1948),
    .B(_03975_));
 sg13g2_nor2_1 _11904_ (.A(_03954_),
    .B(_03976_),
    .Y(_03977_));
 sg13g2_nand2_1 _11905_ (.Y(_03978_),
    .A(net1930),
    .B(_03387_));
 sg13g2_o21ai_1 _11906_ (.B1(_03978_),
    .Y(_03979_),
    .A1(_03540_),
    .A2(_03564_));
 sg13g2_nand2_1 _11907_ (.Y(_03980_),
    .A(net1937),
    .B(_03243_));
 sg13g2_a22oi_1 _11908_ (.Y(_03981_),
    .B1(_03587_),
    .B2(_03671_),
    .A2(_03243_),
    .A1(net1937));
 sg13g2_o21ai_1 _11909_ (.B1(_03980_),
    .Y(_03982_),
    .A1(_03586_),
    .A2(_03672_));
 sg13g2_nor2_1 _11910_ (.A(net1834),
    .B(_03981_),
    .Y(_03983_));
 sg13g2_a21oi_2 _11911_ (.B1(_03983_),
    .Y(_03984_),
    .A2(_03979_),
    .A1(net1830));
 sg13g2_mux2_1 _11912_ (.A0(_03771_),
    .A1(_03821_),
    .S(net1798),
    .X(_03985_));
 sg13g2_nor2_1 _11913_ (.A(net1795),
    .B(_03853_),
    .Y(_03986_));
 sg13g2_a21oi_1 _11914_ (.A1(net1794),
    .A2(_03880_),
    .Y(_03987_),
    .B1(_03986_));
 sg13g2_mux4_1 _11915_ (.S0(net1797),
    .A0(_03771_),
    .A1(_03821_),
    .A2(_03853_),
    .A3(_03881_),
    .S1(net1804),
    .X(_03988_));
 sg13g2_mux2_1 _11916_ (.A0(_03903_),
    .A1(_03929_),
    .S(net1794),
    .X(_03989_));
 sg13g2_and3_1 _11917_ (.X(_03990_),
    .A(net1865),
    .B(net1844),
    .C(_03979_));
 sg13g2_a21oi_2 _11918_ (.B1(_03990_),
    .Y(_03991_),
    .A2(_03982_),
    .A1(net1830));
 sg13g2_mux2_1 _11919_ (.A0(_03991_),
    .A1(_03967_),
    .S(net1820),
    .X(_03992_));
 sg13g2_mux2_1 _11920_ (.A0(_03942_),
    .A1(_03992_),
    .S(net1794),
    .X(_03993_));
 sg13g2_mux2_1 _11921_ (.A0(_03989_),
    .A1(_03993_),
    .S(net1802),
    .X(_03994_));
 sg13g2_a22oi_1 _11922_ (.Y(_03995_),
    .B1(_03994_),
    .B2(net1777),
    .A2(_03661_),
    .A1(net1778));
 sg13g2_o21ai_1 _11923_ (.B1(_03995_),
    .Y(_03996_),
    .A1(_03680_),
    .A2(_03988_));
 sg13g2_xnor2_1 _11924_ (.Y(_03997_),
    .A(net1941),
    .B(_03996_));
 sg13g2_nor2_1 _11925_ (.A(_03984_),
    .B(_03997_),
    .Y(_03998_));
 sg13g2_and2_1 _11926_ (.A(_03984_),
    .B(_03997_),
    .X(_03999_));
 sg13g2_a22oi_1 _11927_ (.Y(_04000_),
    .B1(_03563_),
    .B2(_03687_),
    .A2(_03384_),
    .A1(net1930));
 sg13g2_inv_1 _11928_ (.Y(_04001_),
    .A(_04000_));
 sg13g2_a21oi_1 _11929_ (.A1(net1865),
    .A2(net1845),
    .Y(_04002_),
    .B1(_04000_));
 sg13g2_nand2_1 _11930_ (.Y(_04003_),
    .A(_03671_),
    .B(_03728_));
 sg13g2_o21ai_1 _11931_ (.B1(_04003_),
    .Y(_04004_),
    .A1(net1927),
    .A2(_03241_));
 sg13g2_a21oi_2 _11932_ (.B1(_04002_),
    .Y(_04005_),
    .A2(_04004_),
    .A1(net1837));
 sg13g2_mux2_1 _11933_ (.A0(_03963_),
    .A1(_03965_),
    .S(net1794),
    .X(_04006_));
 sg13g2_nor3_1 _11934_ (.A(net1871),
    .B(net1849),
    .C(_04000_),
    .Y(_04007_));
 sg13g2_a21oi_2 _11935_ (.B1(_04007_),
    .Y(_04008_),
    .A2(_04004_),
    .A1(net1831));
 sg13g2_mux2_1 _11936_ (.A0(_04008_),
    .A1(_03991_),
    .S(net1820),
    .X(_04009_));
 sg13g2_mux2_1 _11937_ (.A0(_03968_),
    .A1(_04009_),
    .S(net1796),
    .X(_04010_));
 sg13g2_mux2_1 _11938_ (.A0(_04006_),
    .A1(_04010_),
    .S(net1802),
    .X(_04011_));
 sg13g2_mux2_1 _11939_ (.A0(_03971_),
    .A1(_03955_),
    .S(net1797),
    .X(_04012_));
 sg13g2_o21ai_1 _11940_ (.B1(net1778),
    .Y(_04013_),
    .A1(_03640_),
    .A2(_04012_));
 sg13g2_mux2_1 _11941_ (.A0(_03956_),
    .A1(_03958_),
    .S(net1796),
    .X(_04014_));
 sg13g2_mux2_1 _11942_ (.A0(_03959_),
    .A1(_03962_),
    .S(net1794),
    .X(_04015_));
 sg13g2_mux2_1 _11943_ (.A0(_04014_),
    .A1(_04015_),
    .S(net1802),
    .X(_04016_));
 sg13g2_a22oi_1 _11944_ (.Y(_04017_),
    .B1(_04016_),
    .B2(_03679_),
    .A2(_04011_),
    .A1(net1777));
 sg13g2_nand2_1 _11945_ (.Y(_04018_),
    .A(_04013_),
    .B(_04017_));
 sg13g2_xnor2_1 _11946_ (.Y(_04019_),
    .A(net1941),
    .B(_04018_));
 sg13g2_nor2_1 _11947_ (.A(_04005_),
    .B(_04019_),
    .Y(_04020_));
 sg13g2_a22oi_1 _11948_ (.Y(_04021_),
    .B1(_03421_),
    .B2(_03746_),
    .A2(_03391_),
    .A1(net1930));
 sg13g2_a21oi_1 _11949_ (.A1(_03437_),
    .A2(net1845),
    .Y(_04022_),
    .B1(_04021_));
 sg13g2_a22oi_1 _11950_ (.Y(_04023_),
    .B1(_03671_),
    .B2(_03763_),
    .A2(_03247_),
    .A1(net1936));
 sg13g2_inv_2 _11951_ (.Y(_04024_),
    .A(_04023_));
 sg13g2_a21oi_1 _11952_ (.A1(net1839),
    .A2(_04024_),
    .Y(_04025_),
    .B1(_04022_));
 sg13g2_mux4_1 _11953_ (.S0(net1798),
    .A0(_03821_),
    .A1(_03853_),
    .A2(_03881_),
    .A3(_03904_),
    .S1(net1804),
    .X(_04026_));
 sg13g2_nand2_1 _11954_ (.Y(_04027_),
    .A(_03639_),
    .B(_03772_));
 sg13g2_nor3_1 _11955_ (.A(net1871),
    .B(net1849),
    .C(_04021_),
    .Y(_04028_));
 sg13g2_a21oi_2 _11956_ (.B1(_04028_),
    .Y(_04029_),
    .A2(_04024_),
    .A1(net1831));
 sg13g2_mux2_1 _11957_ (.A0(_04029_),
    .A1(_04008_),
    .S(net1821),
    .X(_04030_));
 sg13g2_mux2_1 _11958_ (.A0(_03992_),
    .A1(_04030_),
    .S(net1796),
    .X(_04031_));
 sg13g2_mux2_1 _11959_ (.A0(_03943_),
    .A1(_04031_),
    .S(net1804),
    .X(_04032_));
 sg13g2_a22oi_1 _11960_ (.Y(_04033_),
    .B1(_04032_),
    .B2(net1777),
    .A2(_04027_),
    .A1(net1778));
 sg13g2_o21ai_1 _11961_ (.B1(_04033_),
    .Y(_04034_),
    .A1(_03680_),
    .A2(_04026_));
 sg13g2_xnor2_1 _11962_ (.Y(_04035_),
    .A(net1941),
    .B(_04034_));
 sg13g2_nor2_1 _11963_ (.A(_04025_),
    .B(_04035_),
    .Y(_04036_));
 sg13g2_inv_1 _11964_ (.Y(_04037_),
    .A(_04036_));
 sg13g2_a22oi_1 _11965_ (.Y(_04038_),
    .B1(_03421_),
    .B2(_03782_),
    .A2(_03393_),
    .A1(net1930));
 sg13g2_inv_1 _11966_ (.Y(_04039_),
    .A(_04038_));
 sg13g2_nor2_1 _11967_ (.A(net1838),
    .B(_04038_),
    .Y(_04040_));
 sg13g2_a21o_1 _11968_ (.A2(_03251_),
    .A1(net1937),
    .B1(_03671_),
    .X(_04041_));
 sg13g2_and2_1 _11969_ (.A(_03793_),
    .B(_04041_),
    .X(_04042_));
 sg13g2_a21oi_1 _11970_ (.A1(net1839),
    .A2(_04042_),
    .Y(_04043_),
    .B1(_04040_));
 sg13g2_mux2_1 _11971_ (.A0(_03957_),
    .A1(_03972_),
    .S(net1801),
    .X(_04044_));
 sg13g2_o21ai_1 _11972_ (.B1(net1779),
    .Y(_04045_),
    .A1(_03638_),
    .A2(_04044_));
 sg13g2_mux2_1 _11973_ (.A0(_03960_),
    .A1(_03964_),
    .S(net1802),
    .X(_04046_));
 sg13g2_nor3_1 _11974_ (.A(net1871),
    .B(net1849),
    .C(_04038_),
    .Y(_04047_));
 sg13g2_a21oi_2 _11975_ (.B1(_04047_),
    .Y(_04048_),
    .A2(_04042_),
    .A1(net1831));
 sg13g2_mux2_1 _11976_ (.A0(_04048_),
    .A1(_04029_),
    .S(net1821),
    .X(_04049_));
 sg13g2_mux2_1 _11977_ (.A0(_04009_),
    .A1(_04049_),
    .S(net1797),
    .X(_04050_));
 sg13g2_mux2_1 _11978_ (.A0(_03969_),
    .A1(_04050_),
    .S(net1802),
    .X(_04051_));
 sg13g2_a22oi_1 _11979_ (.Y(_04052_),
    .B1(_04051_),
    .B2(_03643_),
    .A2(_04046_),
    .A1(_03679_));
 sg13g2_nand2_1 _11980_ (.Y(_04053_),
    .A(_04045_),
    .B(_04052_));
 sg13g2_xnor2_1 _11981_ (.Y(_04054_),
    .A(net1942),
    .B(_04053_));
 sg13g2_or2_1 _11982_ (.X(_04055_),
    .B(_04054_),
    .A(_04043_));
 sg13g2_a22oi_1 _11983_ (.Y(_04056_),
    .B1(_03563_),
    .B2(_03806_),
    .A2(_03400_),
    .A1(net1931));
 sg13g2_a21oi_1 _11984_ (.A1(net1866),
    .A2(net1846),
    .Y(_04057_),
    .B1(_04056_));
 sg13g2_a22oi_1 _11985_ (.Y(_04058_),
    .B1(_03671_),
    .B2(_03814_),
    .A2(_03258_),
    .A1(net1936));
 sg13g2_inv_2 _11986_ (.Y(_04059_),
    .A(_04058_));
 sg13g2_a21oi_1 _11987_ (.A1(net1839),
    .A2(_04059_),
    .Y(_04060_),
    .B1(_04057_));
 sg13g2_nand2_1 _11988_ (.Y(_04061_),
    .A(net1803),
    .B(_03985_));
 sg13g2_o21ai_1 _11989_ (.B1(_04061_),
    .Y(_04062_),
    .A1(net1803),
    .A2(_03660_));
 sg13g2_nor2b_1 _11990_ (.A(_03610_),
    .B_N(net1799),
    .Y(_04063_));
 sg13g2_nor2_1 _11991_ (.A(net1801),
    .B(_03989_),
    .Y(_04064_));
 sg13g2_a21oi_1 _11992_ (.A1(net1801),
    .A2(_03987_),
    .Y(_04065_),
    .B1(_04064_));
 sg13g2_nor2_1 _11993_ (.A(net1802),
    .B(_03638_),
    .Y(_04066_));
 sg13g2_nor3_1 _11994_ (.A(net1871),
    .B(net1849),
    .C(_04056_),
    .Y(_04067_));
 sg13g2_a21oi_2 _11995_ (.B1(_04067_),
    .Y(_04068_),
    .A2(_04059_),
    .A1(net1831));
 sg13g2_mux2_1 _11996_ (.A0(_04068_),
    .A1(_04048_),
    .S(net1821),
    .X(_04069_));
 sg13g2_mux2_1 _11997_ (.A0(_04030_),
    .A1(_04069_),
    .S(net1796),
    .X(_04070_));
 sg13g2_and2_1 _11998_ (.A(_03639_),
    .B(_04070_),
    .X(_04071_));
 sg13g2_a221oi_1 _11999_ (.B2(_03993_),
    .C1(_04071_),
    .B1(_04066_),
    .A1(_03638_),
    .Y(_04072_),
    .A2(_04065_));
 sg13g2_a22oi_1 _12000_ (.Y(_04073_),
    .B1(_04072_),
    .B2(_03642_),
    .A2(_04063_),
    .A1(_04062_));
 sg13g2_xnor2_1 _12001_ (.Y(_04074_),
    .A(net1947),
    .B(_04073_));
 sg13g2_nor2b_1 _12002_ (.A(_04060_),
    .B_N(_04074_),
    .Y(_04075_));
 sg13g2_inv_1 _12003_ (.Y(_04076_),
    .A(_04075_));
 sg13g2_xnor2_1 _12004_ (.Y(_04077_),
    .A(_04060_),
    .B(_04074_));
 sg13g2_nand2_1 _12005_ (.Y(_04078_),
    .A(net1930),
    .B(_03396_));
 sg13g2_o21ai_1 _12006_ (.B1(_04078_),
    .Y(_04079_),
    .A1(_03564_),
    .A2(_03823_));
 sg13g2_nand2_1 _12007_ (.Y(_04080_),
    .A(net1831),
    .B(_04079_));
 sg13g2_nor2_1 _12008_ (.A(net1926),
    .B(_03254_),
    .Y(_04081_));
 sg13g2_o21ai_1 _12009_ (.B1(_03833_),
    .Y(_04082_),
    .A1(_03671_),
    .A2(_04081_));
 sg13g2_o21ai_1 _12010_ (.B1(_04080_),
    .Y(_04083_),
    .A1(net1831),
    .A2(_04082_));
 sg13g2_mux2_1 _12011_ (.A0(_04012_),
    .A1(_04014_),
    .S(net1803),
    .X(_04084_));
 sg13g2_nor2b_1 _12012_ (.A(_04084_),
    .B_N(_04063_),
    .Y(_04085_));
 sg13g2_mux2_1 _12013_ (.A0(_04006_),
    .A1(_04015_),
    .S(_03634_),
    .X(_04086_));
 sg13g2_a21oi_1 _12014_ (.A1(net1866),
    .A2(net1845),
    .Y(_04087_),
    .B1(_04082_));
 sg13g2_a21oi_1 _12015_ (.A1(net1838),
    .A2(_04079_),
    .Y(_04088_),
    .B1(_04087_));
 sg13g2_a21o_1 _12016_ (.A2(_04079_),
    .A1(net1838),
    .B1(_04087_),
    .X(_04089_));
 sg13g2_mux2_1 _12017_ (.A0(_04088_),
    .A1(_04068_),
    .S(net1822),
    .X(_04090_));
 sg13g2_mux2_1 _12018_ (.A0(_04049_),
    .A1(_04090_),
    .S(net1797),
    .X(_04091_));
 sg13g2_and2_1 _12019_ (.A(_03639_),
    .B(_04091_),
    .X(_04092_));
 sg13g2_a221oi_1 _12020_ (.B2(_03638_),
    .C1(_04092_),
    .B1(_04086_),
    .A1(_04010_),
    .Y(_04093_),
    .A2(_04066_));
 sg13g2_a21oi_1 _12021_ (.A1(_03642_),
    .A2(_04093_),
    .Y(_04094_),
    .B1(_04085_));
 sg13g2_xnor2_1 _12022_ (.Y(_04095_),
    .A(net1947),
    .B(_04094_));
 sg13g2_and2_1 _12023_ (.A(_04083_),
    .B(_04095_),
    .X(_04096_));
 sg13g2_xnor2_1 _12024_ (.Y(_04097_),
    .A(_04083_),
    .B(_04095_));
 sg13g2_and2_1 _12025_ (.A(net1930),
    .B(_03450_),
    .X(_04098_));
 sg13g2_nand2_1 _12026_ (.Y(_04099_),
    .A(net1834),
    .B(_04098_));
 sg13g2_and2_1 _12027_ (.A(net1939),
    .B(_03442_),
    .X(_04100_));
 sg13g2_nand2_1 _12028_ (.Y(_04101_),
    .A(net1939),
    .B(_03442_));
 sg13g2_o21ai_1 _12029_ (.B1(_04099_),
    .Y(_04102_),
    .A1(net1834),
    .A2(_04101_));
 sg13g2_nand2_1 _12030_ (.Y(_04103_),
    .A(_03854_),
    .B(_04063_));
 sg13g2_and2_1 _12031_ (.A(net1840),
    .B(_04098_),
    .X(_04104_));
 sg13g2_nand3_1 _12032_ (.B(net1845),
    .C(_04098_),
    .A(net1866),
    .Y(_04105_));
 sg13g2_a21oi_1 _12033_ (.A1(net1834),
    .A2(_04100_),
    .Y(_04106_),
    .B1(_04104_));
 sg13g2_o21ai_1 _12034_ (.B1(_04105_),
    .Y(_04107_),
    .A1(net1840),
    .A2(_04101_));
 sg13g2_nor2_1 _12035_ (.A(net1821),
    .B(_04107_),
    .Y(_04108_));
 sg13g2_a21oi_1 _12036_ (.A1(net1822),
    .A2(_04088_),
    .Y(_04109_),
    .B1(_04108_));
 sg13g2_mux4_1 _12037_ (.S0(net1798),
    .A0(_04068_),
    .A1(_04106_),
    .A2(_04048_),
    .A3(_04088_),
    .S1(net1822),
    .X(_04110_));
 sg13g2_mux4_1 _12038_ (.S0(net1804),
    .A0(_03905_),
    .A1(_03943_),
    .A2(_04031_),
    .A3(_04110_),
    .S1(net1799),
    .X(_04111_));
 sg13g2_o21ai_1 _12039_ (.B1(_04103_),
    .Y(_04112_),
    .A1(net1779),
    .A2(_04111_));
 sg13g2_xnor2_1 _12040_ (.Y(_04113_),
    .A(net1941),
    .B(_04112_));
 sg13g2_nand2_1 _12041_ (.Y(_04114_),
    .A(_04102_),
    .B(_04113_));
 sg13g2_xor2_1 _12042_ (.B(_04113_),
    .A(_04102_),
    .X(_04115_));
 sg13g2_xnor2_1 _12043_ (.Y(_04116_),
    .A(_04102_),
    .B(_04113_));
 sg13g2_nand2_1 _12044_ (.Y(_04117_),
    .A(_03638_),
    .B(_03970_));
 sg13g2_nand2_1 _12045_ (.Y(_04118_),
    .A(net1822),
    .B(_04107_));
 sg13g2_mux2_1 _12046_ (.A0(_04090_),
    .A1(_04118_),
    .S(net1797),
    .X(_04119_));
 sg13g2_a22oi_1 _12047_ (.Y(_04120_),
    .B1(_04119_),
    .B2(_03639_),
    .A2(_04066_),
    .A1(_04050_));
 sg13g2_nand2_1 _12048_ (.Y(_04121_),
    .A(_04117_),
    .B(_04120_));
 sg13g2_nor2_2 _12049_ (.A(net1801),
    .B(net1800),
    .Y(_04122_));
 sg13g2_nand2b_1 _12050_ (.Y(_04123_),
    .B(_04122_),
    .A_N(_03972_));
 sg13g2_o21ai_1 _12051_ (.B1(_04123_),
    .Y(_04124_),
    .A1(_03638_),
    .A2(_03961_));
 sg13g2_nor2_1 _12052_ (.A(_03642_),
    .B(_04124_),
    .Y(_04125_));
 sg13g2_a21oi_1 _12053_ (.A1(_03642_),
    .A2(_04121_),
    .Y(_04126_),
    .B1(_04125_));
 sg13g2_a21o_1 _12054_ (.A2(_04121_),
    .A1(_03642_),
    .B1(_04125_),
    .X(_04127_));
 sg13g2_and4_1 _12055_ (.A(_03638_),
    .B(_04011_),
    .C(_04032_),
    .D(_04051_),
    .X(_04128_));
 sg13g2_nand3_1 _12056_ (.B(_04110_),
    .C(_04119_),
    .A(_04091_),
    .Y(_04129_));
 sg13g2_nand2_1 _12057_ (.Y(_04130_),
    .A(net1804),
    .B(_03650_));
 sg13g2_o21ai_1 _12058_ (.B1(net1799),
    .Y(_04131_),
    .A1(_04118_),
    .A2(_04130_));
 sg13g2_a21oi_1 _12059_ (.A1(_03634_),
    .A2(_04129_),
    .Y(_04132_),
    .B1(_04131_));
 sg13g2_o21ai_1 _12060_ (.B1(_03642_),
    .Y(_04133_),
    .A1(_04128_),
    .A2(_04132_));
 sg13g2_mux2_1 _12061_ (.A0(_04044_),
    .A1(_04046_),
    .S(net1799),
    .X(_04134_));
 sg13g2_nand4_1 _12062_ (.B(_03769_),
    .C(_03804_),
    .A(_03744_),
    .Y(_04135_),
    .D(_03820_));
 sg13g2_a21oi_1 _12063_ (.A1(net1801),
    .A2(_03654_),
    .Y(_04136_),
    .B1(_04135_));
 sg13g2_o21ai_1 _12064_ (.B1(net1779),
    .Y(_04137_),
    .A1(net1799),
    .A2(_04136_));
 sg13g2_nand2b_1 _12065_ (.Y(_04138_),
    .B(net1800),
    .A_N(_04016_));
 sg13g2_nand2b_1 _12066_ (.Y(_04139_),
    .B(_04122_),
    .A_N(_04012_));
 sg13g2_a22oi_1 _12067_ (.Y(_04140_),
    .B1(_04122_),
    .B2(_03772_),
    .A2(_04026_),
    .A1(net1800));
 sg13g2_nor2b_1 _12068_ (.A(_04137_),
    .B_N(_04140_),
    .Y(_04141_));
 sg13g2_nand4_1 _12069_ (.B(_04138_),
    .C(_04139_),
    .A(_04134_),
    .Y(_04142_),
    .D(_04141_));
 sg13g2_nor3_1 _12070_ (.A(_03838_),
    .B(_03852_),
    .C(_03869_),
    .Y(_04143_));
 sg13g2_a21oi_1 _12071_ (.A1(_03878_),
    .A2(_04143_),
    .Y(_04144_),
    .B1(_03639_));
 sg13g2_nand4_1 _12072_ (.B(_03902_),
    .C(_03916_),
    .A(_03891_),
    .Y(_04145_),
    .D(_03928_));
 sg13g2_o21ai_1 _12073_ (.B1(_03641_),
    .Y(_04146_),
    .A1(_04144_),
    .A2(_04145_));
 sg13g2_o21ai_1 _12074_ (.B1(_03645_),
    .Y(_04147_),
    .A1(_04089_),
    .A2(_04107_));
 sg13g2_nand4_1 _12075_ (.B(_04029_),
    .C(_04048_),
    .A(_04008_),
    .Y(_04148_),
    .D(_04068_));
 sg13g2_nand4_1 _12076_ (.B(_03941_),
    .C(_03967_),
    .A(_03939_),
    .Y(_04149_),
    .D(_03991_));
 sg13g2_o21ai_1 _12077_ (.B1(_03610_),
    .Y(_04150_),
    .A1(net1804),
    .A2(net1799));
 sg13g2_a22oi_1 _12078_ (.Y(_04151_),
    .B1(_04149_),
    .B2(_04150_),
    .A2(_04148_),
    .A1(_03644_));
 sg13g2_nand3_1 _12079_ (.B(_04147_),
    .C(_04151_),
    .A(_04146_),
    .Y(_04152_));
 sg13g2_a21o_2 _12080_ (.A2(_04142_),
    .A1(_04133_),
    .B1(_04152_),
    .X(_04153_));
 sg13g2_a22oi_1 _12081_ (.Y(_04154_),
    .B1(_04122_),
    .B2(_03659_),
    .A2(_03988_),
    .A1(net1800));
 sg13g2_nand2b_1 _12082_ (.Y(_04155_),
    .B(net1801),
    .A_N(_04070_));
 sg13g2_nand3_1 _12083_ (.B(_03650_),
    .C(_04109_),
    .A(net1804),
    .Y(_04156_));
 sg13g2_nand3_1 _12084_ (.B(_04155_),
    .C(_04156_),
    .A(net1777),
    .Y(_04157_));
 sg13g2_a22oi_1 _12085_ (.Y(_04158_),
    .B1(_04154_),
    .B2(net1778),
    .A2(_03994_),
    .A1(_03679_));
 sg13g2_nand2_1 _12086_ (.Y(_04159_),
    .A(_04157_),
    .B(_04158_));
 sg13g2_nand2_1 _12087_ (.Y(_04160_),
    .A(net1947),
    .B(_04159_));
 sg13g2_nor2_1 _12088_ (.A(_04153_),
    .B(_04160_),
    .Y(_04161_));
 sg13g2_nand2_1 _12089_ (.Y(_04162_),
    .A(_04127_),
    .B(_04161_));
 sg13g2_or4_1 _12090_ (.A(_04116_),
    .B(_04126_),
    .C(_04153_),
    .D(_04160_),
    .X(_04163_));
 sg13g2_a21oi_1 _12091_ (.A1(_04114_),
    .A2(_04163_),
    .Y(_04164_),
    .B1(_04097_));
 sg13g2_o21ai_1 _12092_ (.B1(_04077_),
    .Y(_04165_),
    .A1(_04096_),
    .A2(_04164_));
 sg13g2_xor2_1 _12093_ (.B(_04054_),
    .A(_04043_),
    .X(_04166_));
 sg13g2_inv_1 _12094_ (.Y(_04167_),
    .A(_04166_));
 sg13g2_a21o_1 _12095_ (.A2(_04165_),
    .A1(_04076_),
    .B1(_04167_),
    .X(_04168_));
 sg13g2_xor2_1 _12096_ (.B(_04035_),
    .A(_04025_),
    .X(_04169_));
 sg13g2_inv_1 _12097_ (.Y(_04170_),
    .A(_04169_));
 sg13g2_a21o_1 _12098_ (.A2(_04168_),
    .A1(_04055_),
    .B1(_04170_),
    .X(_04171_));
 sg13g2_xor2_1 _12099_ (.B(_04019_),
    .A(_04005_),
    .X(_04172_));
 sg13g2_inv_1 _12100_ (.Y(_04173_),
    .A(_04172_));
 sg13g2_a21oi_1 _12101_ (.A1(_04037_),
    .A2(_04171_),
    .Y(_04174_),
    .B1(_04173_));
 sg13g2_nor2_1 _12102_ (.A(_04020_),
    .B(_04174_),
    .Y(_04175_));
 sg13g2_nor3_1 _12103_ (.A(_03998_),
    .B(_04020_),
    .C(_04174_),
    .Y(_04176_));
 sg13g2_or2_1 _12104_ (.X(_04177_),
    .B(_04176_),
    .A(_03999_));
 sg13g2_xnor2_1 _12105_ (.Y(_04178_),
    .A(_03954_),
    .B(_03976_));
 sg13g2_inv_1 _12106_ (.Y(_04179_),
    .A(_04178_));
 sg13g2_nor2_1 _12107_ (.A(_04177_),
    .B(_04178_),
    .Y(_04180_));
 sg13g2_nor2_1 _12108_ (.A(_03977_),
    .B(_04180_),
    .Y(_04181_));
 sg13g2_nand2_1 _12109_ (.Y(_04182_),
    .A(_03948_),
    .B(_04179_));
 sg13g2_nor3_1 _12110_ (.A(_03999_),
    .B(_04176_),
    .C(_04182_),
    .Y(_04183_));
 sg13g2_a21o_1 _12111_ (.A2(_03977_),
    .A1(_03948_),
    .B1(_03947_),
    .X(_04184_));
 sg13g2_or2_1 _12112_ (.X(_04185_),
    .B(_04184_),
    .A(_04183_));
 sg13g2_a21oi_1 _12113_ (.A1(net1864),
    .A2(net1842),
    .Y(_04186_),
    .B1(_03933_));
 sg13g2_a21oi_2 _12114_ (.B1(_04186_),
    .Y(_04187_),
    .A2(_03938_),
    .A1(net1835));
 sg13g2_nand2b_1 _12115_ (.Y(_04188_),
    .B(_03643_),
    .A_N(_04086_));
 sg13g2_o21ai_1 _12116_ (.B1(_04188_),
    .Y(_04189_),
    .A1(_03680_),
    .A2(_04084_));
 sg13g2_xnor2_1 _12117_ (.Y(_04190_),
    .A(net1941),
    .B(_04189_));
 sg13g2_nand2b_1 _12118_ (.Y(_04191_),
    .B(_04190_),
    .A_N(_04187_));
 sg13g2_xor2_1 _12119_ (.B(_04190_),
    .A(_04187_),
    .X(_04192_));
 sg13g2_nor2_1 _12120_ (.A(net1836),
    .B(_03920_),
    .Y(_04193_));
 sg13g2_a21oi_2 _12121_ (.B1(_04193_),
    .Y(_04194_),
    .A2(_03927_),
    .A1(net1835));
 sg13g2_nand2_1 _12122_ (.Y(_04195_),
    .A(_03679_),
    .B(_04062_));
 sg13g2_o21ai_1 _12123_ (.B1(_04195_),
    .Y(_04196_),
    .A1(_03644_),
    .A2(_04065_));
 sg13g2_xnor2_1 _12124_ (.Y(_04197_),
    .A(net1942),
    .B(_04196_));
 sg13g2_nor2b_1 _12125_ (.A(_04194_),
    .B_N(_04197_),
    .Y(_04198_));
 sg13g2_inv_1 _12126_ (.Y(_04199_),
    .A(_04198_));
 sg13g2_xor2_1 _12127_ (.B(_04197_),
    .A(_04194_),
    .X(_04200_));
 sg13g2_nor2_1 _12128_ (.A(_04192_),
    .B(_04200_),
    .Y(_04201_));
 sg13g2_o21ai_1 _12129_ (.B1(_04201_),
    .Y(_04202_),
    .A1(_04183_),
    .A2(_04184_));
 sg13g2_a21oi_2 _12130_ (.B1(_03896_),
    .Y(_04203_),
    .A2(net1843),
    .A1(net1864));
 sg13g2_nor2_2 _12131_ (.A(net1829),
    .B(_03900_),
    .Y(_04204_));
 sg13g2_nor2_1 _12132_ (.A(net1778),
    .B(_04140_),
    .Y(_04205_));
 sg13g2_xnor2_1 _12133_ (.Y(_04206_),
    .A(net1941),
    .B(_04205_));
 sg13g2_nor3_1 _12134_ (.A(_04203_),
    .B(_04204_),
    .C(_04206_),
    .Y(_04207_));
 sg13g2_a21oi_2 _12135_ (.B1(_03909_),
    .Y(_04208_),
    .A2(net1842),
    .A1(net1863));
 sg13g2_a21oi_2 _12136_ (.B1(_04208_),
    .Y(_04209_),
    .A2(_03915_),
    .A1(net1835));
 sg13g2_nor2_1 _12137_ (.A(net1778),
    .B(_04134_),
    .Y(_04210_));
 sg13g2_xnor2_1 _12138_ (.Y(_04211_),
    .A(net1943),
    .B(_04210_));
 sg13g2_nand2b_1 _12139_ (.Y(_04212_),
    .B(_04211_),
    .A_N(_04209_));
 sg13g2_inv_1 _12140_ (.Y(_04213_),
    .A(_04212_));
 sg13g2_o21ai_1 _12141_ (.B1(_04206_),
    .Y(_04214_),
    .A1(_04203_),
    .A2(_04204_));
 sg13g2_nor2_1 _12142_ (.A(_04191_),
    .B(_04200_),
    .Y(_04215_));
 sg13g2_a21oi_1 _12143_ (.A1(_04212_),
    .A2(_04214_),
    .Y(_04216_),
    .B1(_04207_));
 sg13g2_nor3_1 _12144_ (.A(_04198_),
    .B(_04215_),
    .C(_04216_),
    .Y(_04217_));
 sg13g2_nand2b_1 _12145_ (.Y(_04218_),
    .B(_04209_),
    .A_N(_04211_));
 sg13g2_nand2b_1 _12146_ (.Y(_04219_),
    .B(_04218_),
    .A_N(_04207_));
 sg13g2_a22oi_1 _12147_ (.Y(_04220_),
    .B1(_04219_),
    .B2(_04214_),
    .A2(_04217_),
    .A1(_04202_));
 sg13g2_nor2_1 _12148_ (.A(net1835),
    .B(_03859_),
    .Y(_04221_));
 sg13g2_a21oi_2 _12149_ (.B1(_04221_),
    .Y(_04222_),
    .A2(_03867_),
    .A1(net1835));
 sg13g2_nand2_1 _12150_ (.Y(_04223_),
    .A(_03642_),
    .B(_04124_));
 sg13g2_xnor2_1 _12151_ (.Y(_04224_),
    .A(net1943),
    .B(_04223_));
 sg13g2_nor2_1 _12152_ (.A(_04222_),
    .B(_04224_),
    .Y(_04225_));
 sg13g2_inv_1 _12153_ (.Y(_04226_),
    .A(_04225_));
 sg13g2_xnor2_1 _12154_ (.Y(_04227_),
    .A(_04222_),
    .B(_04224_));
 sg13g2_nand2_1 _12155_ (.Y(_04228_),
    .A(net1777),
    .B(_03854_));
 sg13g2_xnor2_1 _12156_ (.Y(_04229_),
    .A(net1943),
    .B(_04228_));
 sg13g2_nor2_1 _12157_ (.A(net1828),
    .B(_03849_),
    .Y(_04230_));
 sg13g2_a21oi_2 _12158_ (.B1(_04230_),
    .Y(_04231_),
    .A2(_03843_),
    .A1(net1829));
 sg13g2_nand2_1 _12159_ (.Y(_04232_),
    .A(_04229_),
    .B(_04231_));
 sg13g2_nor2_1 _12160_ (.A(_04229_),
    .B(_04231_),
    .Y(_04233_));
 sg13g2_xnor2_1 _12161_ (.Y(_04234_),
    .A(_04229_),
    .B(_04231_));
 sg13g2_nor2_1 _12162_ (.A(_04227_),
    .B(_04234_),
    .Y(_04235_));
 sg13g2_inv_1 _12163_ (.Y(_04236_),
    .A(_04235_));
 sg13g2_nor2_1 _12164_ (.A(net1835),
    .B(_03885_),
    .Y(_04237_));
 sg13g2_a21oi_2 _12165_ (.B1(_04237_),
    .Y(_04238_),
    .A2(_03890_),
    .A1(net1836));
 sg13g2_a21oi_1 _12166_ (.A1(_04138_),
    .A2(_04139_),
    .Y(_04239_),
    .B1(net1778));
 sg13g2_xnor2_1 _12167_ (.Y(_04240_),
    .A(net1947),
    .B(_04239_));
 sg13g2_nor2_1 _12168_ (.A(_04238_),
    .B(_04240_),
    .Y(_04241_));
 sg13g2_xor2_1 _12169_ (.B(_04240_),
    .A(_04238_),
    .X(_04242_));
 sg13g2_a21oi_1 _12170_ (.A1(net1863),
    .A2(net1842),
    .Y(_04243_),
    .B1(_03873_));
 sg13g2_a21oi_2 _12171_ (.B1(_04243_),
    .Y(_04244_),
    .A2(_03877_),
    .A1(net1835));
 sg13g2_nor2_1 _12172_ (.A(net1779),
    .B(_04154_),
    .Y(_04245_));
 sg13g2_xnor2_1 _12173_ (.Y(_04246_),
    .A(net1947),
    .B(_04245_));
 sg13g2_nand2_1 _12174_ (.Y(_04247_),
    .A(_04244_),
    .B(_04246_));
 sg13g2_nor2_1 _12175_ (.A(_04244_),
    .B(_04246_),
    .Y(_04248_));
 sg13g2_xnor2_1 _12176_ (.Y(_04249_),
    .A(_04244_),
    .B(_04246_));
 sg13g2_nor2_1 _12177_ (.A(_04236_),
    .B(_04249_),
    .Y(_04250_));
 sg13g2_nand2_1 _12178_ (.Y(_04251_),
    .A(_04242_),
    .B(_04250_));
 sg13g2_a221oi_1 _12179_ (.B2(_04214_),
    .C1(_04251_),
    .B1(_04219_),
    .A1(_04202_),
    .Y(_04252_),
    .A2(_04217_));
 sg13g2_o21ai_1 _12180_ (.B1(_04247_),
    .Y(_04253_),
    .A1(_04241_),
    .A2(_04248_));
 sg13g2_o21ai_1 _12181_ (.B1(_04232_),
    .Y(_04254_),
    .A1(_04225_),
    .A2(_04233_));
 sg13g2_o21ai_1 _12182_ (.B1(_04254_),
    .Y(_04255_),
    .A1(_04236_),
    .A2(_04253_));
 sg13g2_nor2_1 _12183_ (.A(_04252_),
    .B(_04255_),
    .Y(_04256_));
 sg13g2_mux2_1 _12184_ (.A0(_03788_),
    .A1(_03803_),
    .S(net1838),
    .X(_04257_));
 sg13g2_nor2_1 _12185_ (.A(_03644_),
    .B(_04044_),
    .Y(_04258_));
 sg13g2_xnor2_1 _12186_ (.Y(_04259_),
    .A(net1948),
    .B(_04258_));
 sg13g2_inv_1 _12187_ (.Y(_04260_),
    .A(_04259_));
 sg13g2_nand2_1 _12188_ (.Y(_04261_),
    .A(_04257_),
    .B(_04260_));
 sg13g2_xnor2_1 _12189_ (.Y(_04262_),
    .A(_04257_),
    .B(_04259_));
 sg13g2_nand3_1 _12190_ (.B(net1777),
    .C(_03772_),
    .A(net1803),
    .Y(_04263_));
 sg13g2_xnor2_1 _12191_ (.Y(_04264_),
    .A(net1948),
    .B(_04263_));
 sg13g2_nor2_1 _12192_ (.A(net1838),
    .B(_03758_),
    .Y(_04265_));
 sg13g2_a21o_1 _12193_ (.A2(_03768_),
    .A1(net1838),
    .B1(_04265_),
    .X(_04266_));
 sg13g2_nor2_1 _12194_ (.A(_04264_),
    .B(_04266_),
    .Y(_04267_));
 sg13g2_nand2_1 _12195_ (.Y(_04268_),
    .A(_04264_),
    .B(_04266_));
 sg13g2_nor2b_1 _12196_ (.A(_04267_),
    .B_N(_04268_),
    .Y(_04269_));
 sg13g2_nand2_1 _12197_ (.Y(_04270_),
    .A(_04262_),
    .B(_04269_));
 sg13g2_inv_1 _12198_ (.Y(_04271_),
    .A(_04270_));
 sg13g2_nor2_2 _12199_ (.A(net1836),
    .B(_03828_),
    .Y(_04272_));
 sg13g2_a21oi_2 _12200_ (.B1(_04272_),
    .Y(_04273_),
    .A2(_03836_),
    .A1(net1836));
 sg13g2_nor2_1 _12201_ (.A(_03644_),
    .B(_04084_),
    .Y(_04274_));
 sg13g2_xnor2_1 _12202_ (.Y(_04275_),
    .A(net1948),
    .B(_04274_));
 sg13g2_nor2_1 _12203_ (.A(_04273_),
    .B(_04275_),
    .Y(_04276_));
 sg13g2_inv_1 _12204_ (.Y(_04277_),
    .A(_04276_));
 sg13g2_xnor2_1 _12205_ (.Y(_04278_),
    .A(_04273_),
    .B(_04275_));
 sg13g2_nor2_1 _12206_ (.A(net1838),
    .B(_03810_),
    .Y(_04279_));
 sg13g2_a21oi_2 _12207_ (.B1(_04279_),
    .Y(_04280_),
    .A2(_03819_),
    .A1(net1838));
 sg13g2_nand2_1 _12208_ (.Y(_04281_),
    .A(net1777),
    .B(_04062_));
 sg13g2_xnor2_1 _12209_ (.Y(_04282_),
    .A(net1943),
    .B(_04281_));
 sg13g2_xor2_1 _12210_ (.B(_04282_),
    .A(_04280_),
    .X(_04283_));
 sg13g2_nand2b_1 _12211_ (.Y(_04284_),
    .B(_04283_),
    .A_N(_04278_));
 sg13g2_nor2_1 _12212_ (.A(_04270_),
    .B(_04284_),
    .Y(_04285_));
 sg13g2_o21ai_1 _12213_ (.B1(_04285_),
    .Y(_04286_),
    .A1(_04252_),
    .A2(_04255_));
 sg13g2_a21o_1 _12214_ (.A2(_04282_),
    .A1(_04280_),
    .B1(_04277_),
    .X(_04287_));
 sg13g2_o21ai_1 _12215_ (.B1(_04287_),
    .Y(_04288_),
    .A1(_04280_),
    .A2(_04282_));
 sg13g2_inv_1 _12216_ (.Y(_04289_),
    .A(_04288_));
 sg13g2_a21oi_1 _12217_ (.A1(_04261_),
    .A2(_04268_),
    .Y(_04290_),
    .B1(_04267_));
 sg13g2_a21oi_1 _12218_ (.A1(_04271_),
    .A2(_04288_),
    .Y(_04291_),
    .B1(_04290_));
 sg13g2_nor2_1 _12219_ (.A(_03645_),
    .B(_04012_),
    .Y(_04292_));
 sg13g2_xnor2_1 _12220_ (.Y(_04293_),
    .A(net1947),
    .B(_04292_));
 sg13g2_nand2_1 _12221_ (.Y(_04294_),
    .A(net1839),
    .B(_03743_));
 sg13g2_o21ai_1 _12222_ (.B1(_04294_),
    .Y(_04295_),
    .A1(net1839),
    .A2(_03710_));
 sg13g2_nand2b_1 _12223_ (.Y(_04296_),
    .B(_04295_),
    .A_N(_04293_));
 sg13g2_xor2_1 _12224_ (.B(_04295_),
    .A(_04293_),
    .X(_04297_));
 sg13g2_a21o_1 _12225_ (.A2(_04291_),
    .A1(_04286_),
    .B1(_04297_),
    .X(_04298_));
 sg13g2_or2_1 _12226_ (.X(_04299_),
    .B(_03663_),
    .A(_03600_));
 sg13g2_and2_1 _12227_ (.A(_04296_),
    .B(_04299_),
    .X(_04300_));
 sg13g2_a22oi_1 _12228_ (.Y(_04301_),
    .B1(_04298_),
    .B2(_04300_),
    .A2(_03663_),
    .A1(_03600_));
 sg13g2_or2_1 _12229_ (.X(_04302_),
    .B(_03453_),
    .A(_03445_));
 sg13g2_nor2_2 _12230_ (.A(_03645_),
    .B(_03972_),
    .Y(_04303_));
 sg13g2_nor2_1 _12231_ (.A(net1949),
    .B(_04303_),
    .Y(_04304_));
 sg13g2_xnor2_1 _12232_ (.Y(_04305_),
    .A(net1950),
    .B(_04303_));
 sg13g2_xnor2_1 _12233_ (.Y(_04306_),
    .A(_04302_),
    .B(_04305_));
 sg13g2_nand2_1 _12234_ (.Y(_04307_),
    .A(_04301_),
    .B(_04306_));
 sg13g2_xnor2_1 _12235_ (.Y(_04308_),
    .A(_04301_),
    .B(_04306_));
 sg13g2_nand2_1 _12236_ (.Y(_04309_),
    .A(net1949),
    .B(_04308_));
 sg13g2_nor3_2 _12237_ (.A(net1946),
    .B(_03645_),
    .C(_03650_),
    .Y(_04310_));
 sg13g2_or3_1 _12238_ (.A(net1946),
    .B(_03645_),
    .C(_03650_),
    .X(_04311_));
 sg13g2_a21oi_1 _12239_ (.A1(_04304_),
    .A2(_04307_),
    .Y(_04312_),
    .B1(net1774));
 sg13g2_a21oi_2 _12240_ (.B1(_03622_),
    .Y(_04313_),
    .A2(net1843),
    .A1(net1864));
 sg13g2_a21oi_1 _12241_ (.A1(net1865),
    .A2(net1844),
    .Y(_04314_),
    .B1(net1877));
 sg13g2_a221oi_1 _12242_ (.B2(net1825),
    .C1(_03940_),
    .B1(_03979_),
    .A1(_03622_),
    .Y(_04315_),
    .A2(_03951_));
 sg13g2_nor2_1 _12243_ (.A(_03953_),
    .B(_04315_),
    .Y(_04316_));
 sg13g2_nand2_1 _12244_ (.Y(_04317_),
    .A(_03953_),
    .B(_04315_));
 sg13g2_xor2_1 _12245_ (.B(_04315_),
    .A(_03953_),
    .X(_04318_));
 sg13g2_a221oi_1 _12246_ (.B2(_03979_),
    .C1(_03966_),
    .B1(net1824),
    .A1(net1877),
    .Y(_04319_),
    .A2(_04002_));
 sg13g2_nor2_1 _12247_ (.A(_03982_),
    .B(_04319_),
    .Y(_04320_));
 sg13g2_xnor2_1 _12248_ (.Y(_04321_),
    .A(_03981_),
    .B(_04319_));
 sg13g2_and2_1 _12249_ (.A(_04318_),
    .B(_04321_),
    .X(_04322_));
 sg13g2_nand2_1 _12250_ (.Y(_04323_),
    .A(_04318_),
    .B(_04321_));
 sg13g2_a221oi_1 _12251_ (.B2(_04039_),
    .C1(_04028_),
    .B1(net1823),
    .A1(net1877),
    .Y(_04324_),
    .A2(_04057_));
 sg13g2_nor2_1 _12252_ (.A(_04042_),
    .B(_04324_),
    .Y(_04325_));
 sg13g2_nand2_1 _12253_ (.Y(_04326_),
    .A(_04042_),
    .B(_04324_));
 sg13g2_a221oi_1 _12254_ (.B2(net1825),
    .C1(_04047_),
    .B1(_04079_),
    .A1(_03622_),
    .Y(_04327_),
    .A2(_04057_));
 sg13g2_nor2_1 _12255_ (.A(_04059_),
    .B(_04327_),
    .Y(_04328_));
 sg13g2_a221oi_1 _12256_ (.B2(_04079_),
    .C1(_04067_),
    .B1(net1823),
    .A1(_04098_),
    .Y(_04329_),
    .A2(net1825));
 sg13g2_nand2b_1 _12257_ (.Y(_04330_),
    .B(_04082_),
    .A_N(_04329_));
 sg13g2_a22oi_1 _12258_ (.Y(_04331_),
    .B1(_04098_),
    .B2(net1823),
    .A2(_04079_),
    .A1(net1840));
 sg13g2_and2_1 _12259_ (.A(_04100_),
    .B(_04331_),
    .X(_04332_));
 sg13g2_nor2b_1 _12260_ (.A(_04082_),
    .B_N(_04329_),
    .Y(_04333_));
 sg13g2_xnor2_1 _12261_ (.Y(_04334_),
    .A(_04082_),
    .B(_04329_));
 sg13g2_o21ai_1 _12262_ (.B1(_04330_),
    .Y(_04335_),
    .A1(_04332_),
    .A2(_04333_));
 sg13g2_xnor2_1 _12263_ (.Y(_04336_),
    .A(_04058_),
    .B(_04327_));
 sg13g2_a21oi_1 _12264_ (.A1(_04335_),
    .A2(_04336_),
    .Y(_04337_),
    .B1(_04328_));
 sg13g2_xor2_1 _12265_ (.B(_04324_),
    .A(_04042_),
    .X(_04338_));
 sg13g2_and2_1 _12266_ (.A(_04336_),
    .B(_04338_),
    .X(_04339_));
 sg13g2_a221oi_1 _12267_ (.B2(_04339_),
    .C1(_04325_),
    .B1(_04335_),
    .A1(_04326_),
    .Y(_04340_),
    .A2(_04328_));
 sg13g2_a221oi_1 _12268_ (.B2(_04001_),
    .C1(_03990_),
    .B1(net1823),
    .A1(net1877),
    .Y(_04341_),
    .A2(_04022_));
 sg13g2_nor2_1 _12269_ (.A(_04004_),
    .B(_04341_),
    .Y(_04342_));
 sg13g2_nand2_1 _12270_ (.Y(_04343_),
    .A(_04004_),
    .B(_04341_));
 sg13g2_xnor2_1 _12271_ (.Y(_04344_),
    .A(_04004_),
    .B(_04341_));
 sg13g2_a221oi_1 _12272_ (.B2(net1826),
    .C1(_04007_),
    .B1(_04039_),
    .A1(_03622_),
    .Y(_04345_),
    .A2(_04022_));
 sg13g2_nor2_1 _12273_ (.A(_04024_),
    .B(_04345_),
    .Y(_04346_));
 sg13g2_inv_1 _12274_ (.Y(_04347_),
    .A(_04346_));
 sg13g2_xnor2_1 _12275_ (.Y(_04348_),
    .A(_04023_),
    .B(_04345_));
 sg13g2_inv_1 _12276_ (.Y(_04349_),
    .A(_04348_));
 sg13g2_nand2b_1 _12277_ (.Y(_04350_),
    .B(_04348_),
    .A_N(_04344_));
 sg13g2_a21o_1 _12278_ (.A2(_04346_),
    .A1(_04343_),
    .B1(_04342_),
    .X(_04351_));
 sg13g2_a21oi_1 _12279_ (.A1(_04343_),
    .A2(_04346_),
    .Y(_04352_),
    .B1(_04342_));
 sg13g2_or2_1 _12280_ (.X(_04353_),
    .B(_04350_),
    .A(_04323_));
 sg13g2_a221oi_1 _12281_ (.B2(_04351_),
    .C1(_04316_),
    .B1(_04322_),
    .A1(_04317_),
    .Y(_04354_),
    .A2(_04320_));
 sg13g2_o21ai_1 _12282_ (.B1(_04354_),
    .Y(_04355_),
    .A1(_04340_),
    .A2(_04353_));
 sg13g2_a221oi_1 _12283_ (.B2(_03511_),
    .C1(_03920_),
    .B1(_03604_),
    .A1(net1863),
    .Y(_04356_),
    .A2(net1842));
 sg13g2_a221oi_1 _12284_ (.B2(_03622_),
    .C1(_04356_),
    .B1(_04208_),
    .A1(net1836),
    .Y(_04357_),
    .A2(_03895_));
 sg13g2_nand2b_1 _12285_ (.Y(_04358_),
    .B(_03914_),
    .A_N(_04357_));
 sg13g2_and2_1 _12286_ (.A(_03915_),
    .B(_04357_),
    .X(_04359_));
 sg13g2_xnor2_1 _12287_ (.Y(_04360_),
    .A(_03915_),
    .B(_04357_));
 sg13g2_a221oi_1 _12288_ (.B2(_03921_),
    .C1(_03910_),
    .B1(net1824),
    .A1(net1876),
    .Y(_04361_),
    .A2(_04186_));
 sg13g2_nand2b_1 _12289_ (.Y(_04362_),
    .B(_03926_),
    .A_N(_04361_));
 sg13g2_xnor2_1 _12290_ (.Y(_04363_),
    .A(_03927_),
    .B(_04361_));
 sg13g2_a221oi_1 _12291_ (.B2(_03511_),
    .C1(_03669_),
    .B1(_03604_),
    .A1(net1863),
    .Y(_04364_),
    .A2(net1843));
 sg13g2_a221oi_1 _12292_ (.B2(_03932_),
    .C1(net1876),
    .B1(_03930_),
    .A1(net1863),
    .Y(_04365_),
    .A2(net1842));
 sg13g2_or3_1 _12293_ (.A(_03922_),
    .B(_04364_),
    .C(_04365_),
    .X(_04366_));
 sg13g2_nor2_1 _12294_ (.A(_03937_),
    .B(_04366_),
    .Y(_04367_));
 sg13g2_xnor2_1 _12295_ (.Y(_04368_),
    .A(_03938_),
    .B(_04366_));
 sg13g2_a221oi_1 _12296_ (.B2(_03511_),
    .C1(_03950_),
    .B1(_03604_),
    .A1(net1865),
    .Y(_04369_),
    .A2(net1843));
 sg13g2_a221oi_1 _12297_ (.B2(_03668_),
    .C1(net1876),
    .B1(_03664_),
    .A1(net1863),
    .Y(_04370_),
    .A2(net1842));
 sg13g2_nor3_1 _12298_ (.A(_03934_),
    .B(_04369_),
    .C(_04370_),
    .Y(_04371_));
 sg13g2_or3_1 _12299_ (.A(_03934_),
    .B(_04369_),
    .C(_04370_),
    .X(_04372_));
 sg13g2_nor2_1 _12300_ (.A(_03677_),
    .B(_04371_),
    .Y(_04373_));
 sg13g2_xnor2_1 _12301_ (.Y(_04374_),
    .A(_03676_),
    .B(_04371_));
 sg13g2_nand2_1 _12302_ (.Y(_04375_),
    .A(_04368_),
    .B(_04374_));
 sg13g2_inv_1 _12303_ (.Y(_04376_),
    .A(_04375_));
 sg13g2_nor3_1 _12304_ (.A(_04360_),
    .B(_04363_),
    .C(_04375_),
    .Y(_04377_));
 sg13g2_a221oi_1 _12305_ (.B2(_03872_),
    .C1(net1876),
    .B1(_03870_),
    .A1(net1863),
    .Y(_04378_),
    .A2(net1842));
 sg13g2_a221oi_1 _12306_ (.B2(net1825),
    .C1(_04378_),
    .B1(_03886_),
    .A1(net1835),
    .Y(_04379_),
    .A2(_03860_));
 sg13g2_nor2_1 _12307_ (.A(_03877_),
    .B(_04379_),
    .Y(_04380_));
 sg13g2_xor2_1 _12308_ (.B(_04379_),
    .A(_03877_),
    .X(_04381_));
 sg13g2_xnor2_1 _12309_ (.Y(_04382_),
    .A(_03877_),
    .B(_04379_));
 sg13g2_a221oi_1 _12310_ (.B2(_03860_),
    .C1(_03844_),
    .B1(net1824),
    .A1(net1876),
    .Y(_04383_),
    .A2(_04243_));
 sg13g2_nor2_1 _12311_ (.A(_03867_),
    .B(_04383_),
    .Y(_04384_));
 sg13g2_nand2_1 _12312_ (.Y(_04385_),
    .A(_03867_),
    .B(_04383_));
 sg13g2_xor2_1 _12313_ (.B(_04383_),
    .A(_03867_),
    .X(_04386_));
 sg13g2_and2_1 _12314_ (.A(_04381_),
    .B(_04386_),
    .X(_04387_));
 sg13g2_a221oi_1 _12315_ (.B2(_03895_),
    .C1(_03887_),
    .B1(net1824),
    .A1(net1876),
    .Y(_04388_),
    .A2(_04208_));
 sg13g2_nand2b_1 _12316_ (.Y(_04389_),
    .B(_03900_),
    .A_N(_04388_));
 sg13g2_xnor2_1 _12317_ (.Y(_04390_),
    .A(_03900_),
    .B(_04388_));
 sg13g2_a221oi_1 _12318_ (.B2(_03886_),
    .C1(_03874_),
    .B1(net1824),
    .A1(net1876),
    .Y(_04391_),
    .A2(_04203_));
 sg13g2_and2_1 _12319_ (.A(_03890_),
    .B(_04391_),
    .X(_04392_));
 sg13g2_or2_1 _12320_ (.X(_04393_),
    .B(_04391_),
    .A(_03890_));
 sg13g2_xor2_1 _12321_ (.B(_04391_),
    .A(_03890_),
    .X(_04394_));
 sg13g2_and4_1 _12322_ (.A(_04381_),
    .B(_04386_),
    .C(_04390_),
    .D(_04394_),
    .X(_04395_));
 sg13g2_and2_1 _12323_ (.A(_04377_),
    .B(_04395_),
    .X(_04396_));
 sg13g2_a22oi_1 _12324_ (.Y(_04397_),
    .B1(_04372_),
    .B2(_03676_),
    .A2(_04366_),
    .A1(_03937_));
 sg13g2_nor2_1 _12325_ (.A(_04367_),
    .B(_04397_),
    .Y(_04398_));
 sg13g2_nor4_1 _12326_ (.A(_04360_),
    .B(_04363_),
    .C(_04367_),
    .D(_04397_),
    .Y(_04399_));
 sg13g2_o21ai_1 _12327_ (.B1(_04358_),
    .Y(_04400_),
    .A1(_04359_),
    .A2(_04362_));
 sg13g2_or2_1 _12328_ (.X(_04401_),
    .B(_04400_),
    .A(_04399_));
 sg13g2_o21ai_1 _12329_ (.B1(_04395_),
    .Y(_04402_),
    .A1(_04399_),
    .A2(_04400_));
 sg13g2_and2_1 _12330_ (.A(_04389_),
    .B(_04393_),
    .X(_04403_));
 sg13g2_a21oi_1 _12331_ (.A1(_04389_),
    .A2(_04393_),
    .Y(_04404_),
    .B1(_04392_));
 sg13g2_a221oi_1 _12332_ (.B2(_04404_),
    .C1(_04384_),
    .B1(_04387_),
    .A1(_04380_),
    .Y(_04405_),
    .A2(_04385_));
 sg13g2_nand2_1 _12333_ (.Y(_04406_),
    .A(_04402_),
    .B(_04405_));
 sg13g2_a21oi_1 _12334_ (.A1(_04355_),
    .A2(_04396_),
    .Y(_04407_),
    .B1(_04406_));
 sg13g2_a21o_1 _12335_ (.A2(_04396_),
    .A1(_04355_),
    .B1(_04406_),
    .X(_04408_));
 sg13g2_a221oi_1 _12336_ (.B2(_03843_),
    .C1(_03829_),
    .B1(net1824),
    .A1(_03860_),
    .Y(_04409_),
    .A2(net1825));
 sg13g2_nand2b_1 _12337_ (.Y(_04410_),
    .B(_03849_),
    .A_N(_04409_));
 sg13g2_inv_1 _12338_ (.Y(_04411_),
    .A(_04410_));
 sg13g2_xnor2_1 _12339_ (.Y(_04412_),
    .A(_03849_),
    .B(_04409_));
 sg13g2_nand2_1 _12340_ (.Y(_04413_),
    .A(_03843_),
    .B(net1825));
 sg13g2_a22oi_1 _12341_ (.Y(_04414_),
    .B1(_04272_),
    .B2(_03622_),
    .A2(_03811_),
    .A1(net1836));
 sg13g2_and3_1 _12342_ (.X(_04415_),
    .A(_03836_),
    .B(_04413_),
    .C(_04414_));
 sg13g2_nand3_1 _12343_ (.B(_04413_),
    .C(_04414_),
    .A(_03836_),
    .Y(_04416_));
 sg13g2_a21oi_1 _12344_ (.A1(_04413_),
    .A2(_04414_),
    .Y(_04417_),
    .B1(_03836_));
 sg13g2_nor2_1 _12345_ (.A(_04415_),
    .B(_04417_),
    .Y(_04418_));
 sg13g2_nand2_1 _12346_ (.Y(_04419_),
    .A(_04412_),
    .B(_04418_));
 sg13g2_inv_1 _12347_ (.Y(_04420_),
    .A(_04419_));
 sg13g2_o21ai_1 _12348_ (.B1(_04416_),
    .Y(_04421_),
    .A1(_04411_),
    .A2(_04417_));
 sg13g2_nand2_1 _12349_ (.Y(_04422_),
    .A(_03811_),
    .B(net1825));
 sg13g2_a21oi_1 _12350_ (.A1(_03788_),
    .A2(net1823),
    .Y(_04423_),
    .B1(_03759_));
 sg13g2_and3_1 _12351_ (.X(_04424_),
    .A(_03803_),
    .B(_04422_),
    .C(_04423_));
 sg13g2_nand2_1 _12352_ (.Y(_04425_),
    .A(net1876),
    .B(_04272_));
 sg13g2_a21oi_1 _12353_ (.A1(_03811_),
    .A2(net1823),
    .Y(_04426_),
    .B1(_03789_));
 sg13g2_a21oi_1 _12354_ (.A1(_04425_),
    .A2(_04426_),
    .Y(_04427_),
    .B1(_03819_));
 sg13g2_a21oi_1 _12355_ (.A1(_04422_),
    .A2(_04423_),
    .Y(_04428_),
    .B1(_03803_));
 sg13g2_nor2_1 _12356_ (.A(_04427_),
    .B(_04428_),
    .Y(_04429_));
 sg13g2_o21ai_1 _12357_ (.B1(_04421_),
    .Y(_04430_),
    .A1(_04424_),
    .A2(_04429_));
 sg13g2_a21oi_1 _12358_ (.A1(_04408_),
    .A2(_04420_),
    .Y(_04431_),
    .B1(_04430_));
 sg13g2_and3_1 _12359_ (.X(_04432_),
    .A(_03819_),
    .B(_04425_),
    .C(_04426_));
 sg13g2_nand2b_1 _12360_ (.Y(_04433_),
    .B(_04432_),
    .A_N(_04428_));
 sg13g2_nand2b_1 _12361_ (.Y(_04434_),
    .B(_04433_),
    .A_N(_04424_));
 sg13g2_nor2_1 _12362_ (.A(_04431_),
    .B(_04434_),
    .Y(_04435_));
 sg13g2_a221oi_1 _12363_ (.B2(_03566_),
    .C1(_03653_),
    .B1(net1823),
    .A1(_03709_),
    .Y(_04436_),
    .A2(net1826));
 sg13g2_or2_1 _12364_ (.X(_04437_),
    .B(_04436_),
    .A(_03599_));
 sg13g2_xnor2_1 _12365_ (.Y(_04438_),
    .A(_03599_),
    .B(_04436_));
 sg13g2_a22oi_1 _12366_ (.Y(_04439_),
    .B1(net1823),
    .B2(_03453_),
    .A2(net1826),
    .A1(_03566_));
 sg13g2_nor2_1 _12367_ (.A(_03445_),
    .B(_04439_),
    .Y(_04440_));
 sg13g2_xor2_1 _12368_ (.B(_04439_),
    .A(_03445_),
    .X(_04441_));
 sg13g2_nor2b_1 _12369_ (.A(_04438_),
    .B_N(_04441_),
    .Y(_04442_));
 sg13g2_a221oi_1 _12370_ (.B2(_03788_),
    .C1(_03711_),
    .B1(net1825),
    .A1(_03622_),
    .Y(_04443_),
    .A2(_04265_));
 sg13g2_nor2_1 _12371_ (.A(_03768_),
    .B(_04443_),
    .Y(_04444_));
 sg13g2_xnor2_1 _12372_ (.Y(_04445_),
    .A(_03768_),
    .B(_04443_));
 sg13g2_inv_1 _12373_ (.Y(_04446_),
    .A(_04445_));
 sg13g2_nand2b_1 _12374_ (.Y(_04447_),
    .B(net1826),
    .A_N(_03758_));
 sg13g2_a21oi_1 _12375_ (.A1(_03709_),
    .A2(net1824),
    .Y(_04448_),
    .B1(_03655_));
 sg13g2_a21oi_1 _12376_ (.A1(_04447_),
    .A2(_04448_),
    .Y(_04449_),
    .B1(_03743_));
 sg13g2_nand3_1 _12377_ (.B(_04447_),
    .C(_04448_),
    .A(_03743_),
    .Y(_04450_));
 sg13g2_nand2b_1 _12378_ (.Y(_04451_),
    .B(_04450_),
    .A_N(_04449_));
 sg13g2_nor2_1 _12379_ (.A(_04445_),
    .B(_04451_),
    .Y(_04452_));
 sg13g2_nand2_1 _12380_ (.Y(_04453_),
    .A(_04442_),
    .B(_04452_));
 sg13g2_nor3_2 _12381_ (.A(_04431_),
    .B(_04434_),
    .C(_04453_),
    .Y(_04454_));
 sg13g2_a21oi_1 _12382_ (.A1(_04444_),
    .A2(_04450_),
    .Y(_04455_),
    .B1(_04449_));
 sg13g2_inv_1 _12383_ (.Y(_04456_),
    .A(_04455_));
 sg13g2_a21oi_1 _12384_ (.A1(_03445_),
    .A2(_04439_),
    .Y(_04457_),
    .B1(_04437_));
 sg13g2_a21oi_1 _12385_ (.A1(_04442_),
    .A2(_04456_),
    .Y(_04458_),
    .B1(_04440_));
 sg13g2_nand2b_2 _12386_ (.Y(_04459_),
    .B(_04458_),
    .A_N(_04457_));
 sg13g2_o21ai_1 _12387_ (.B1(net1827),
    .Y(_04460_),
    .A1(_04454_),
    .A2(_04459_));
 sg13g2_inv_1 _12388_ (.Y(_04461_),
    .A(_04460_));
 sg13g2_nor3_1 _12389_ (.A(net1827),
    .B(_04454_),
    .C(_04459_),
    .Y(_04462_));
 sg13g2_or3_1 _12390_ (.A(net1827),
    .B(_04454_),
    .C(_04459_),
    .X(_04463_));
 sg13g2_a21o_1 _12391_ (.A2(_04452_),
    .A1(_04435_),
    .B1(_04456_),
    .X(_04464_));
 sg13g2_nand2b_1 _12392_ (.Y(_04465_),
    .B(_04464_),
    .A_N(_04438_));
 sg13g2_xor2_1 _12393_ (.B(_04464_),
    .A(_04438_),
    .X(_04466_));
 sg13g2_or2_1 _12394_ (.X(_04467_),
    .B(_04466_),
    .A(_04463_));
 sg13g2_a21oi_1 _12395_ (.A1(_04435_),
    .A2(_04446_),
    .Y(_04468_),
    .B1(_04444_));
 sg13g2_xnor2_1 _12396_ (.Y(_04469_),
    .A(_04451_),
    .B(_04468_));
 sg13g2_inv_1 _12397_ (.Y(_04470_),
    .A(_04469_));
 sg13g2_xnor2_1 _12398_ (.Y(_04471_),
    .A(_04407_),
    .B(_04412_));
 sg13g2_a21oi_1 _12399_ (.A1(_04355_),
    .A2(_04377_),
    .Y(_04472_),
    .B1(_04401_));
 sg13g2_nand2b_1 _12400_ (.Y(_04473_),
    .B(_04390_),
    .A_N(_04472_));
 sg13g2_a21oi_1 _12401_ (.A1(_04403_),
    .A2(_04473_),
    .Y(_04474_),
    .B1(_04392_));
 sg13g2_a221oi_1 _12402_ (.B2(_04473_),
    .C1(_04382_),
    .B1(_04403_),
    .A1(_03890_),
    .Y(_04475_),
    .A2(_04391_));
 sg13g2_or3_1 _12403_ (.A(_04380_),
    .B(_04386_),
    .C(_04475_),
    .X(_04476_));
 sg13g2_o21ai_1 _12404_ (.B1(_04386_),
    .Y(_04477_),
    .A1(_04380_),
    .A2(_04475_));
 sg13g2_nand2_1 _12405_ (.Y(_04478_),
    .A(_04476_),
    .B(_04477_));
 sg13g2_a21oi_2 _12406_ (.B1(_04471_),
    .Y(_04479_),
    .A2(_04477_),
    .A1(_04476_));
 sg13g2_xnor2_1 _12407_ (.Y(_04480_),
    .A(_04382_),
    .B(_04474_));
 sg13g2_nand2_1 _12408_ (.Y(_04481_),
    .A(_04389_),
    .B(_04473_));
 sg13g2_xor2_1 _12409_ (.B(_04481_),
    .A(_04394_),
    .X(_04482_));
 sg13g2_xor2_1 _12410_ (.B(_04374_),
    .A(_04355_),
    .X(_04483_));
 sg13g2_o21ai_1 _12411_ (.B1(_04352_),
    .Y(_04484_),
    .A1(_04340_),
    .A2(_04350_));
 sg13g2_xnor2_1 _12412_ (.Y(_04485_),
    .A(_04321_),
    .B(_04484_));
 sg13g2_xnor2_1 _12413_ (.Y(_04486_),
    .A(_04100_),
    .B(_04331_));
 sg13g2_nor2_1 _12414_ (.A(_04104_),
    .B(_04486_),
    .Y(_04487_));
 sg13g2_xnor2_1 _12415_ (.Y(_04488_),
    .A(_04332_),
    .B(_04334_));
 sg13g2_inv_1 _12416_ (.Y(_04489_),
    .A(_04488_));
 sg13g2_nand2b_1 _12417_ (.Y(_04490_),
    .B(_04487_),
    .A_N(_04488_));
 sg13g2_xnor2_1 _12418_ (.Y(_04491_),
    .A(_04335_),
    .B(_04336_));
 sg13g2_nand2b_2 _12419_ (.Y(_04492_),
    .B(_04491_),
    .A_N(_04490_));
 sg13g2_xnor2_1 _12420_ (.Y(_04493_),
    .A(_04337_),
    .B(_04338_));
 sg13g2_inv_1 _12421_ (.Y(_04494_),
    .A(_04493_));
 sg13g2_xnor2_1 _12422_ (.Y(_04495_),
    .A(_04340_),
    .B(_04348_));
 sg13g2_nor3_1 _12423_ (.A(_04492_),
    .B(_04493_),
    .C(_04495_),
    .Y(_04496_));
 sg13g2_inv_1 _12424_ (.Y(_04497_),
    .A(_04496_));
 sg13g2_o21ai_1 _12425_ (.B1(_04347_),
    .Y(_04498_),
    .A1(_04340_),
    .A2(_04349_));
 sg13g2_xor2_1 _12426_ (.B(_04498_),
    .A(_04344_),
    .X(_04499_));
 sg13g2_and2_1 _12427_ (.A(_04496_),
    .B(_04499_),
    .X(_04500_));
 sg13g2_nand3_1 _12428_ (.B(_04496_),
    .C(_04499_),
    .A(_04485_),
    .Y(_04501_));
 sg13g2_inv_1 _12429_ (.Y(_04502_),
    .A(_04501_));
 sg13g2_a21oi_1 _12430_ (.A1(_04321_),
    .A2(_04484_),
    .Y(_04503_),
    .B1(_04320_));
 sg13g2_xnor2_1 _12431_ (.Y(_04504_),
    .A(_04318_),
    .B(_04503_));
 sg13g2_nor2_1 _12432_ (.A(_04501_),
    .B(_04504_),
    .Y(_04505_));
 sg13g2_nor3_1 _12433_ (.A(_04483_),
    .B(_04501_),
    .C(_04504_),
    .Y(_04506_));
 sg13g2_a21oi_1 _12434_ (.A1(_04355_),
    .A2(_04374_),
    .Y(_04507_),
    .B1(_04373_));
 sg13g2_xnor2_1 _12435_ (.Y(_04508_),
    .A(_04368_),
    .B(_04507_));
 sg13g2_nor4_2 _12436_ (.A(_04483_),
    .B(_04501_),
    .C(_04504_),
    .Y(_04509_),
    .D(_04508_));
 sg13g2_a21oi_1 _12437_ (.A1(_04355_),
    .A2(_04376_),
    .Y(_04510_),
    .B1(_04398_));
 sg13g2_xnor2_1 _12438_ (.Y(_04511_),
    .A(_04363_),
    .B(_04510_));
 sg13g2_nand2_1 _12439_ (.Y(_04512_),
    .A(_04509_),
    .B(_04511_));
 sg13g2_o21ai_1 _12440_ (.B1(_04362_),
    .Y(_04513_),
    .A1(_04363_),
    .A2(_04510_));
 sg13g2_xor2_1 _12441_ (.B(_04513_),
    .A(_04360_),
    .X(_04514_));
 sg13g2_nand3_1 _12442_ (.B(_04511_),
    .C(_04514_),
    .A(_04509_),
    .Y(_04515_));
 sg13g2_nand2_1 _12443_ (.Y(_04516_),
    .A(net1728),
    .B(_04515_));
 sg13g2_xnor2_1 _12444_ (.Y(_04517_),
    .A(_04390_),
    .B(_04472_));
 sg13g2_inv_1 _12445_ (.Y(_04518_),
    .A(_04517_));
 sg13g2_nand4_1 _12446_ (.B(_04511_),
    .C(_04514_),
    .A(_04509_),
    .Y(_04519_),
    .D(_04518_));
 sg13g2_nand2_1 _12447_ (.Y(_04520_),
    .A(net1728),
    .B(_04519_));
 sg13g2_nor3_2 _12448_ (.A(_04480_),
    .B(_04482_),
    .C(_04519_),
    .Y(_04521_));
 sg13g2_a21oi_1 _12449_ (.A1(_04479_),
    .A2(_04521_),
    .Y(_04522_),
    .B1(_04463_));
 sg13g2_or2_1 _12450_ (.X(_04523_),
    .B(_04432_),
    .A(_04427_));
 sg13g2_inv_1 _12451_ (.Y(_04524_),
    .A(_04523_));
 sg13g2_o21ai_1 _12452_ (.B1(_04421_),
    .Y(_04525_),
    .A1(_04407_),
    .A2(_04419_));
 sg13g2_xnor2_1 _12453_ (.Y(_04526_),
    .A(_04524_),
    .B(_04525_));
 sg13g2_a21oi_1 _12454_ (.A1(_04408_),
    .A2(_04412_),
    .Y(_04527_),
    .B1(_04411_));
 sg13g2_xor2_1 _12455_ (.B(_04527_),
    .A(_04418_),
    .X(_04528_));
 sg13g2_and2_1 _12456_ (.A(_04526_),
    .B(_04528_),
    .X(_04529_));
 sg13g2_nand3_1 _12457_ (.B(_04521_),
    .C(_04529_),
    .A(_04479_),
    .Y(_04530_));
 sg13g2_nand2_1 _12458_ (.Y(_04531_),
    .A(net1728),
    .B(_04530_));
 sg13g2_xnor2_1 _12459_ (.Y(_04532_),
    .A(_04435_),
    .B(_04445_));
 sg13g2_nor2_1 _12460_ (.A(_04424_),
    .B(_04428_),
    .Y(_04533_));
 sg13g2_a21oi_1 _12461_ (.A1(_04524_),
    .A2(_04525_),
    .Y(_04534_),
    .B1(_04427_));
 sg13g2_xor2_1 _12462_ (.B(_04534_),
    .A(_04533_),
    .X(_04535_));
 sg13g2_inv_1 _12463_ (.Y(_04536_),
    .A(_04535_));
 sg13g2_nor2b_1 _12464_ (.A(_04532_),
    .B_N(_04535_),
    .Y(_04537_));
 sg13g2_nand4_1 _12465_ (.B(_04521_),
    .C(_04529_),
    .A(_04479_),
    .Y(_04538_),
    .D(_04537_));
 sg13g2_nand2_1 _12466_ (.Y(_04539_),
    .A(net1728),
    .B(_04538_));
 sg13g2_o21ai_1 _12467_ (.B1(net1728),
    .Y(_04540_),
    .A1(_04470_),
    .A2(_04538_));
 sg13g2_and2_1 _12468_ (.A(_04437_),
    .B(_04465_),
    .X(_04541_));
 sg13g2_xor2_1 _12469_ (.B(_04541_),
    .A(_04441_),
    .X(_04542_));
 sg13g2_a21o_2 _12470_ (.A2(_04540_),
    .A1(_04467_),
    .B1(_04542_),
    .X(_04543_));
 sg13g2_nand3_1 _12471_ (.B(_04540_),
    .C(_04542_),
    .A(_04467_),
    .Y(_04544_));
 sg13g2_a21oi_1 _12472_ (.A1(_04543_),
    .A2(_04544_),
    .Y(_04545_),
    .B1(_04461_));
 sg13g2_xnor2_1 _12473_ (.Y(_04546_),
    .A(_04470_),
    .B(_04539_));
 sg13g2_xnor2_1 _12474_ (.Y(_04547_),
    .A(_04466_),
    .B(_04540_));
 sg13g2_nor2b_1 _12475_ (.A(_04546_),
    .B_N(_04547_),
    .Y(_04548_));
 sg13g2_and2_1 _12476_ (.A(_04545_),
    .B(_04548_),
    .X(_04549_));
 sg13g2_o21ai_1 _12477_ (.B1(net1728),
    .Y(_04550_),
    .A1(_04530_),
    .A2(_04536_));
 sg13g2_xor2_1 _12478_ (.B(_04550_),
    .A(_04532_),
    .X(_04551_));
 sg13g2_xnor2_1 _12479_ (.Y(_04552_),
    .A(_04532_),
    .B(_04550_));
 sg13g2_xnor2_1 _12480_ (.Y(_04553_),
    .A(_04531_),
    .B(_04535_));
 sg13g2_xnor2_1 _12481_ (.Y(_04554_),
    .A(_04531_),
    .B(_04536_));
 sg13g2_nor2_1 _12482_ (.A(_04552_),
    .B(_04554_),
    .Y(_04555_));
 sg13g2_nand3_1 _12483_ (.B(_04521_),
    .C(_04528_),
    .A(_04479_),
    .Y(_04556_));
 sg13g2_nand2_1 _12484_ (.Y(_04557_),
    .A(net1729),
    .B(_04556_));
 sg13g2_xor2_1 _12485_ (.B(_04557_),
    .A(_04526_),
    .X(_04558_));
 sg13g2_xnor2_1 _12486_ (.Y(_04559_),
    .A(_04526_),
    .B(_04557_));
 sg13g2_xnor2_1 _12487_ (.Y(_04560_),
    .A(_04522_),
    .B(_04528_));
 sg13g2_nand2b_1 _12488_ (.Y(_04561_),
    .B(_04559_),
    .A_N(_04560_));
 sg13g2_nor4_2 _12489_ (.A(_04552_),
    .B(_04554_),
    .C(_04558_),
    .Y(_04562_),
    .D(_04560_));
 sg13g2_xnor2_1 _12490_ (.Y(_04563_),
    .A(_04516_),
    .B(_04518_));
 sg13g2_nand2_1 _12491_ (.Y(_04564_),
    .A(net1728),
    .B(_04512_));
 sg13g2_xnor2_1 _12492_ (.Y(_04565_),
    .A(_04514_),
    .B(_04564_));
 sg13g2_nand2_1 _12493_ (.Y(_04566_),
    .A(_04563_),
    .B(_04565_));
 sg13g2_nor4_1 _12494_ (.A(net1827),
    .B(_04454_),
    .C(_04459_),
    .D(_04509_),
    .Y(_04567_));
 sg13g2_xnor2_1 _12495_ (.Y(_04568_),
    .A(_04511_),
    .B(_04567_));
 sg13g2_nor4_1 _12496_ (.A(net1827),
    .B(_04454_),
    .C(_04459_),
    .D(_04506_),
    .Y(_04569_));
 sg13g2_xor2_1 _12497_ (.B(_04569_),
    .A(_04508_),
    .X(_04570_));
 sg13g2_nor2_1 _12498_ (.A(_04568_),
    .B(_04570_),
    .Y(_04571_));
 sg13g2_nand3_1 _12499_ (.B(_04565_),
    .C(_04571_),
    .A(_04563_),
    .Y(_04572_));
 sg13g2_nor2_1 _12500_ (.A(_04463_),
    .B(_04521_),
    .Y(_04573_));
 sg13g2_a21oi_1 _12501_ (.A1(_04478_),
    .A2(_04521_),
    .Y(_04574_),
    .B1(_04463_));
 sg13g2_xor2_1 _12502_ (.B(_04574_),
    .A(_04471_),
    .X(_04575_));
 sg13g2_xnor2_1 _12503_ (.Y(_04576_),
    .A(_04471_),
    .B(_04574_));
 sg13g2_xnor2_1 _12504_ (.Y(_04577_),
    .A(_04478_),
    .B(_04573_));
 sg13g2_nand2b_1 _12505_ (.Y(_04578_),
    .B(_04576_),
    .A_N(_04577_));
 sg13g2_xor2_1 _12506_ (.B(_04520_),
    .A(_04482_),
    .X(_04579_));
 sg13g2_o21ai_1 _12507_ (.B1(net1728),
    .Y(_04580_),
    .A1(_04482_),
    .A2(_04519_));
 sg13g2_xor2_1 _12508_ (.B(_04580_),
    .A(_04480_),
    .X(_04581_));
 sg13g2_nand2_1 _12509_ (.Y(_04582_),
    .A(_04579_),
    .B(_04581_));
 sg13g2_inv_1 _12510_ (.Y(_04583_),
    .A(_04582_));
 sg13g2_nor4_1 _12511_ (.A(_04572_),
    .B(_04575_),
    .C(_04577_),
    .D(_04582_),
    .Y(_04584_));
 sg13g2_nand3_1 _12512_ (.B(_04562_),
    .C(_04584_),
    .A(_04549_),
    .Y(_04585_));
 sg13g2_xnor2_1 _12513_ (.Y(_04586_),
    .A(_04492_),
    .B(_04493_));
 sg13g2_nand2b_1 _12514_ (.Y(_04587_),
    .B(_04494_),
    .A_N(net1727));
 sg13g2_nand2_1 _12515_ (.Y(_04588_),
    .A(net1727),
    .B(_04586_));
 sg13g2_mux2_1 _12516_ (.A0(_04494_),
    .A1(_04586_),
    .S(net1727),
    .X(_04589_));
 sg13g2_inv_1 _12517_ (.Y(_04590_),
    .A(_04589_));
 sg13g2_o21ai_1 _12518_ (.B1(_04495_),
    .Y(_04591_),
    .A1(_04492_),
    .A2(_04493_));
 sg13g2_nor2b_1 _12519_ (.A(_04496_),
    .B_N(_04591_),
    .Y(_04592_));
 sg13g2_mux2_1 _12520_ (.A0(_04495_),
    .A1(_04592_),
    .S(net1727),
    .X(_04593_));
 sg13g2_xor2_1 _12521_ (.B(_04488_),
    .A(_04487_),
    .X(_04594_));
 sg13g2_mux2_1 _12522_ (.A0(_04489_),
    .A1(_04594_),
    .S(net1727),
    .X(_04595_));
 sg13g2_inv_1 _12523_ (.Y(_04596_),
    .A(_04595_));
 sg13g2_xor2_1 _12524_ (.B(_04491_),
    .A(_04490_),
    .X(_04597_));
 sg13g2_mux2_1 _12525_ (.A0(_04491_),
    .A1(_04597_),
    .S(net1727),
    .X(_04598_));
 sg13g2_nand2_1 _12526_ (.Y(_04599_),
    .A(_04595_),
    .B(_04598_));
 sg13g2_or3_1 _12527_ (.A(_04590_),
    .B(_04593_),
    .C(_04599_),
    .X(_04600_));
 sg13g2_nor4_1 _12528_ (.A(net1827),
    .B(_04454_),
    .C(_04459_),
    .D(_04505_),
    .Y(_04601_));
 sg13g2_xnor2_1 _12529_ (.Y(_04602_),
    .A(_04483_),
    .B(_04601_));
 sg13g2_nor4_1 _12530_ (.A(_04313_),
    .B(_04454_),
    .C(_04459_),
    .D(_04502_),
    .Y(_04603_));
 sg13g2_xor2_1 _12531_ (.B(_04603_),
    .A(_04504_),
    .X(_04604_));
 sg13g2_xnor2_1 _12532_ (.Y(_04605_),
    .A(_04504_),
    .B(_04603_));
 sg13g2_and2_1 _12533_ (.A(_04602_),
    .B(_04605_),
    .X(_04606_));
 sg13g2_nand2_1 _12534_ (.Y(_04607_),
    .A(_04602_),
    .B(_04605_));
 sg13g2_a21o_1 _12535_ (.A2(_04497_),
    .A1(net1727),
    .B1(_04499_),
    .X(_04608_));
 sg13g2_nand3_1 _12536_ (.B(_04497_),
    .C(_04499_),
    .A(net1727),
    .Y(_04609_));
 sg13g2_nand2_1 _12537_ (.Y(_04610_),
    .A(_04608_),
    .B(_04609_));
 sg13g2_nor4_1 _12538_ (.A(_04313_),
    .B(_04454_),
    .C(_04459_),
    .D(_04500_),
    .Y(_04611_));
 sg13g2_xor2_1 _12539_ (.B(_04611_),
    .A(_04485_),
    .X(_04612_));
 sg13g2_nand3_1 _12540_ (.B(_04609_),
    .C(_04612_),
    .A(_04608_),
    .Y(_04613_));
 sg13g2_nor2_1 _12541_ (.A(_04607_),
    .B(_04613_),
    .Y(_04614_));
 sg13g2_nand2b_1 _12542_ (.Y(_04615_),
    .B(_04614_),
    .A_N(_04600_));
 sg13g2_nand2_1 _12543_ (.Y(_04616_),
    .A(_04584_),
    .B(_04615_));
 sg13g2_and3_1 _12544_ (.X(_04617_),
    .A(_04549_),
    .B(_04562_),
    .C(_04616_));
 sg13g2_nand4_1 _12545_ (.B(_04548_),
    .C(_04562_),
    .A(_04545_),
    .Y(_04618_),
    .D(_04616_));
 sg13g2_a21oi_1 _12546_ (.A1(_04600_),
    .A2(_04614_),
    .Y(_04619_),
    .B1(_04572_));
 sg13g2_nor3_1 _12547_ (.A(_04578_),
    .B(_04582_),
    .C(_04619_),
    .Y(_04620_));
 sg13g2_nand2b_2 _12548_ (.Y(_04621_),
    .B(_04562_),
    .A_N(_04620_));
 sg13g2_and2_1 _12549_ (.A(_04549_),
    .B(_04621_),
    .X(_04622_));
 sg13g2_nand2_1 _12550_ (.Y(_04623_),
    .A(_04549_),
    .B(_04621_));
 sg13g2_a221oi_1 _12551_ (.B2(_04598_),
    .C1(_04593_),
    .B1(_04595_),
    .A1(_04587_),
    .Y(_04624_),
    .A2(_04588_));
 sg13g2_o21ai_1 _12552_ (.B1(_04606_),
    .Y(_04625_),
    .A1(_04613_),
    .A2(_04624_));
 sg13g2_a21o_1 _12553_ (.A2(_04625_),
    .A1(_04571_),
    .B1(_04566_),
    .X(_04626_));
 sg13g2_a21oi_1 _12554_ (.A1(_04583_),
    .A2(_04626_),
    .Y(_04627_),
    .B1(_04578_));
 sg13g2_o21ai_1 _12555_ (.B1(_04555_),
    .Y(_04628_),
    .A1(_04561_),
    .A2(_04627_));
 sg13g2_a221oi_1 _12556_ (.B2(_04628_),
    .C1(_04461_),
    .B1(_04548_),
    .A1(_04543_),
    .Y(_04629_),
    .A2(_04544_));
 sg13g2_nand2_1 _12557_ (.Y(_04630_),
    .A(_04598_),
    .B(net1707));
 sg13g2_o21ai_1 _12558_ (.B1(_04630_),
    .Y(_04631_),
    .A1(_04593_),
    .A2(net1707));
 sg13g2_and2_1 _12559_ (.A(net1720),
    .B(_04631_),
    .X(_04632_));
 sg13g2_mux2_1 _12560_ (.A0(_04602_),
    .A1(_04612_),
    .S(net1710),
    .X(_04633_));
 sg13g2_a21oi_1 _12561_ (.A1(net1719),
    .A2(_04633_),
    .Y(_04634_),
    .B1(_04632_));
 sg13g2_xnor2_1 _12562_ (.Y(_04635_),
    .A(_04105_),
    .B(_04486_));
 sg13g2_nor2b_1 _12563_ (.A(net1708),
    .B_N(_04635_),
    .Y(_04636_));
 sg13g2_nand2_2 _12564_ (.Y(_04637_),
    .A(net1716),
    .B(_04636_));
 sg13g2_inv_1 _12565_ (.Y(_04638_),
    .A(_04637_));
 sg13g2_nor2_1 _12566_ (.A(net1721),
    .B(_04634_),
    .Y(_04639_));
 sg13g2_a21oi_1 _12567_ (.A1(net1721),
    .A2(_04637_),
    .Y(_04640_),
    .B1(_04639_));
 sg13g2_nor2_1 _12568_ (.A(_04563_),
    .B(net1711),
    .Y(_04641_));
 sg13g2_a21oi_1 _12569_ (.A1(_04568_),
    .A2(net1710),
    .Y(_04642_),
    .B1(_04641_));
 sg13g2_nand2_1 _12570_ (.Y(_04643_),
    .A(_04581_),
    .B(net1714));
 sg13g2_o21ai_1 _12571_ (.B1(_04643_),
    .Y(_04644_),
    .A1(_04575_),
    .A2(net1714));
 sg13g2_mux2_1 _12572_ (.A0(_04642_),
    .A1(_04644_),
    .S(net1718),
    .X(_04645_));
 sg13g2_inv_1 _12573_ (.Y(_04646_),
    .A(_04645_));
 sg13g2_mux2_1 _12574_ (.A0(_04551_),
    .A1(_04559_),
    .S(net1712),
    .X(_04647_));
 sg13g2_nor2_1 _12575_ (.A(net1718),
    .B(_04647_),
    .Y(_04648_));
 sg13g2_a21oi_1 _12576_ (.A1(_04543_),
    .A2(_04544_),
    .Y(_04649_),
    .B1(_04547_));
 sg13g2_nor3_1 _12577_ (.A(_04461_),
    .B(_04648_),
    .C(_04649_),
    .Y(_04650_));
 sg13g2_inv_1 _12578_ (.Y(_04651_),
    .A(_04650_));
 sg13g2_mux4_1 _12579_ (.S0(net1723),
    .A0(_04634_),
    .A1(_04638_),
    .A2(_04651_),
    .A3(_04646_),
    .S1(_04585_),
    .X(_04652_));
 sg13g2_and2_1 _12580_ (.A(net1775),
    .B(_04652_),
    .X(_04653_));
 sg13g2_a21oi_1 _12581_ (.A1(_04309_),
    .A2(_04312_),
    .Y(_04654_),
    .B1(_04653_));
 sg13g2_a21o_1 _12582_ (.A2(_04312_),
    .A1(_04309_),
    .B1(_04653_),
    .X(_04655_));
 sg13g2_nor2_1 _12583_ (.A(net1941),
    .B(_04159_),
    .Y(_04656_));
 sg13g2_a221oi_1 _12584_ (.B2(_04656_),
    .C1(_04161_),
    .B1(_04153_),
    .A1(net1942),
    .Y(_04657_),
    .A2(_04127_));
 sg13g2_and2_1 _12585_ (.A(net1774),
    .B(_04585_),
    .X(_04658_));
 sg13g2_nand2_2 _12586_ (.Y(_04659_),
    .A(net1774),
    .B(_04585_));
 sg13g2_nor2_1 _12587_ (.A(_04105_),
    .B(net1707),
    .Y(_04660_));
 sg13g2_nand2_1 _12588_ (.Y(_04661_),
    .A(net1715),
    .B(_04660_));
 sg13g2_nor2_1 _12589_ (.A(net1724),
    .B(_04661_),
    .Y(_04662_));
 sg13g2_nor2_1 _12590_ (.A(net1773),
    .B(net1725),
    .Y(_04663_));
 sg13g2_a21o_2 _12591_ (.A2(_04662_),
    .A1(_04658_),
    .B1(_04657_),
    .X(_04664_));
 sg13g2_nand3_1 _12592_ (.B(_04157_),
    .C(_04158_),
    .A(net1941),
    .Y(_04665_));
 sg13g2_nand2b_2 _12593_ (.Y(_04666_),
    .B(_04665_),
    .A_N(_04153_));
 sg13g2_o21ai_1 _12594_ (.B1(_03296_),
    .Y(_04667_),
    .A1(_03435_),
    .A2(net1776));
 sg13g2_inv_1 _12595_ (.Y(_04668_),
    .A(_04667_));
 sg13g2_nor2_1 _12596_ (.A(net1773),
    .B(_04585_),
    .Y(_04669_));
 sg13g2_or2_1 _12597_ (.X(_04670_),
    .B(_04585_),
    .A(net1773));
 sg13g2_nor2_1 _12598_ (.A(net1840),
    .B(net1776),
    .Y(_04671_));
 sg13g2_mux2_1 _12599_ (.A0(_03466_),
    .A1(_03465_),
    .S(net1764),
    .X(_04672_));
 sg13g2_and2_1 _12600_ (.A(net1704),
    .B(_04672_),
    .X(_04673_));
 sg13g2_nor2_1 _12601_ (.A(_03480_),
    .B(net1765),
    .Y(_04674_));
 sg13g2_a221oi_1 _12602_ (.B2(_03481_),
    .C1(_04674_),
    .B1(net1765),
    .A1(net1776),
    .Y(_04675_),
    .A2(net1709));
 sg13g2_nor2_1 _12603_ (.A(net1944),
    .B(net1775),
    .Y(_04676_));
 sg13g2_nand2_2 _12604_ (.Y(_04677_),
    .A(net1950),
    .B(net1773));
 sg13g2_nor2_1 _12605_ (.A(_03496_),
    .B(net1764),
    .Y(_04678_));
 sg13g2_a21oi_2 _12606_ (.B1(_04678_),
    .Y(_04679_),
    .A2(net1764),
    .A1(_03510_));
 sg13g2_nand2b_2 _12607_ (.Y(_04680_),
    .B(net1761),
    .A_N(_04679_));
 sg13g2_nand3_1 _12608_ (.B(net1709),
    .C(_04674_),
    .A(net1776),
    .Y(_04681_));
 sg13g2_nand2b_1 _12609_ (.Y(_04682_),
    .B(_04681_),
    .A_N(_04675_));
 sg13g2_a21oi_2 _12610_ (.B1(_04675_),
    .Y(_04683_),
    .A2(_04681_),
    .A1(_04680_));
 sg13g2_nand3_1 _12611_ (.B(_04549_),
    .C(_04621_),
    .A(net1775),
    .Y(_04684_));
 sg13g2_mux2_1 _12612_ (.A0(_03476_),
    .A1(_03474_),
    .S(net1764),
    .X(_04685_));
 sg13g2_and2_1 _12613_ (.A(_04684_),
    .B(_04685_),
    .X(_04686_));
 sg13g2_nand2_1 _12614_ (.Y(_04687_),
    .A(_04684_),
    .B(_04685_));
 sg13g2_xnor2_1 _12615_ (.Y(_04688_),
    .A(_04684_),
    .B(_04685_));
 sg13g2_nand2_1 _12616_ (.Y(_04689_),
    .A(_03471_),
    .B(net1764));
 sg13g2_o21ai_1 _12617_ (.B1(_04689_),
    .Y(_04690_),
    .A1(_03469_),
    .A2(net1764));
 sg13g2_inv_1 _12618_ (.Y(_04691_),
    .A(_04690_));
 sg13g2_nand2_1 _12619_ (.Y(_04692_),
    .A(net1706),
    .B(_04691_));
 sg13g2_nor2_1 _12620_ (.A(net1706),
    .B(_04691_),
    .Y(_04693_));
 sg13g2_xnor2_1 _12621_ (.Y(_04694_),
    .A(net1706),
    .B(_04691_));
 sg13g2_or2_1 _12622_ (.X(_04695_),
    .B(_04694_),
    .A(_04688_));
 sg13g2_o21ai_1 _12623_ (.B1(_04692_),
    .Y(_04696_),
    .A1(_04686_),
    .A2(_04693_));
 sg13g2_o21ai_1 _12624_ (.B1(_04696_),
    .Y(_04697_),
    .A1(_04683_),
    .A2(_04695_));
 sg13g2_xnor2_1 _12625_ (.Y(_04698_),
    .A(net1704),
    .B(_04672_));
 sg13g2_inv_1 _12626_ (.Y(_04699_),
    .A(_04698_));
 sg13g2_a21oi_1 _12627_ (.A1(_04697_),
    .A2(_04699_),
    .Y(_04700_),
    .B1(_04673_));
 sg13g2_or2_1 _12628_ (.X(_04701_),
    .B(net1764),
    .A(_03461_));
 sg13g2_nand2b_1 _12629_ (.Y(_04702_),
    .B(net1764),
    .A_N(_03462_));
 sg13g2_nand2_1 _12630_ (.Y(_04703_),
    .A(_04701_),
    .B(_04702_));
 sg13g2_a221oi_1 _12631_ (.B2(_04702_),
    .C1(_04673_),
    .B1(_04701_),
    .A1(_04697_),
    .Y(_04704_),
    .A2(_04699_));
 sg13g2_nand2_1 _12632_ (.Y(_04705_),
    .A(_03457_),
    .B(net1765));
 sg13g2_o21ai_1 _12633_ (.B1(_04705_),
    .Y(_04706_),
    .A1(_03448_),
    .A2(net1765));
 sg13g2_nor2_1 _12634_ (.A(_03439_),
    .B(net1765),
    .Y(_04707_));
 sg13g2_a21oi_1 _12635_ (.A1(_03438_),
    .A2(net1765),
    .Y(_04708_),
    .B1(_04707_));
 sg13g2_and3_1 _12636_ (.X(_04709_),
    .A(_04704_),
    .B(_04706_),
    .C(_04708_));
 sg13g2_or2_1 _12637_ (.X(_04710_),
    .B(_04709_),
    .A(_04668_));
 sg13g2_xnor2_1 _12638_ (.Y(_04711_),
    .A(_04700_),
    .B(_04703_));
 sg13g2_xnor2_1 _12639_ (.Y(_04712_),
    .A(_04697_),
    .B(_04699_));
 sg13g2_inv_2 _12640_ (.Y(_04713_),
    .A(_04712_));
 sg13g2_nand2_1 _12641_ (.Y(_04714_),
    .A(_04706_),
    .B(_04712_));
 sg13g2_xor2_1 _12642_ (.B(_04682_),
    .A(_04680_),
    .X(_04715_));
 sg13g2_xnor2_1 _12643_ (.Y(_04716_),
    .A(_04683_),
    .B(_04688_));
 sg13g2_nand2_1 _12644_ (.Y(_04717_),
    .A(_04715_),
    .B(net1702));
 sg13g2_o21ai_1 _12645_ (.B1(_04687_),
    .Y(_04718_),
    .A1(_04683_),
    .A2(_04688_));
 sg13g2_xor2_1 _12646_ (.B(_04718_),
    .A(_04694_),
    .X(_04719_));
 sg13g2_xnor2_1 _12647_ (.Y(_04720_),
    .A(_04694_),
    .B(_04718_));
 sg13g2_nand2b_1 _12648_ (.Y(_04721_),
    .B(_04719_),
    .A_N(_04717_));
 sg13g2_nor3_1 _12649_ (.A(_04711_),
    .B(_04714_),
    .C(_04721_),
    .Y(_04722_));
 sg13g2_a21oi_1 _12650_ (.A1(_04704_),
    .A2(_04706_),
    .Y(_04723_),
    .B1(_04708_));
 sg13g2_nor2_1 _12651_ (.A(_04709_),
    .B(_04723_),
    .Y(_04724_));
 sg13g2_or2_1 _12652_ (.X(_04725_),
    .B(_04723_),
    .A(_04709_));
 sg13g2_o21ai_1 _12653_ (.B1(_04710_),
    .Y(_04726_),
    .A1(_04722_),
    .A2(_04724_));
 sg13g2_and2_1 _12654_ (.A(net1696),
    .B(_04726_),
    .X(_04727_));
 sg13g2_nor2_1 _12655_ (.A(net1721),
    .B(_04637_),
    .Y(_04728_));
 sg13g2_nor2_1 _12656_ (.A(net1773),
    .B(_04728_),
    .Y(_04729_));
 sg13g2_o21ai_1 _12657_ (.B1(_04126_),
    .Y(_04730_),
    .A1(_04153_),
    .A2(_04160_));
 sg13g2_a21oi_1 _12658_ (.A1(_04127_),
    .A2(_04161_),
    .Y(_04731_),
    .B1(_04677_));
 sg13g2_xnor2_1 _12659_ (.Y(_04732_),
    .A(_04116_),
    .B(_04162_));
 sg13g2_a22oi_1 _12660_ (.Y(_04733_),
    .B1(_04730_),
    .B2(_04731_),
    .A2(_04115_),
    .A1(net1942));
 sg13g2_a21oi_1 _12661_ (.A1(_04659_),
    .A2(_04733_),
    .Y(_04734_),
    .B1(_04729_));
 sg13g2_inv_1 _12662_ (.Y(_04735_),
    .A(_04734_));
 sg13g2_and3_2 _12663_ (.X(_04736_),
    .A(net1696),
    .B(_04726_),
    .C(_04735_));
 sg13g2_nor2_1 _12664_ (.A(_04596_),
    .B(net1708),
    .Y(_04737_));
 sg13g2_a21oi_1 _12665_ (.A1(_04105_),
    .A2(net1708),
    .Y(_04738_),
    .B1(_04737_));
 sg13g2_nand2_1 _12666_ (.Y(_04739_),
    .A(net1715),
    .B(_04738_));
 sg13g2_nor2_1 _12667_ (.A(net1721),
    .B(_04739_),
    .Y(_04740_));
 sg13g2_nand3_1 _12668_ (.B(_04114_),
    .C(_04163_),
    .A(_04097_),
    .Y(_04741_));
 sg13g2_nand2b_2 _12669_ (.Y(_04742_),
    .B(_04741_),
    .A_N(_04164_));
 sg13g2_a221oi_1 _12670_ (.B2(net1946),
    .C1(net1705),
    .B1(_04742_),
    .A1(net1761),
    .Y(_04743_),
    .A2(_04732_));
 sg13g2_o21ai_1 _12671_ (.B1(_04743_),
    .Y(_04744_),
    .A1(net1773),
    .A2(_04740_));
 sg13g2_inv_1 _12672_ (.Y(_04745_),
    .A(_04744_));
 sg13g2_xnor2_1 _12673_ (.Y(_04746_),
    .A(net1761),
    .B(_04679_));
 sg13g2_xnor2_1 _12674_ (.Y(_04747_),
    .A(_04677_),
    .B(_04679_));
 sg13g2_nor2_2 _12675_ (.A(_04682_),
    .B(_04747_),
    .Y(_04748_));
 sg13g2_nand3_1 _12676_ (.B(_04719_),
    .C(_04748_),
    .A(net1702),
    .Y(_04749_));
 sg13g2_nor3_1 _12677_ (.A(_04711_),
    .B(_04714_),
    .C(_04749_),
    .Y(_04750_));
 sg13g2_o21ai_1 _12678_ (.B1(_04710_),
    .Y(_04751_),
    .A1(_04724_),
    .A2(_04750_));
 sg13g2_and2_1 _12679_ (.A(_04744_),
    .B(_04751_),
    .X(_04752_));
 sg13g2_nor2_1 _12680_ (.A(_04727_),
    .B(_04735_),
    .Y(_04753_));
 sg13g2_a21oi_1 _12681_ (.A1(_04664_),
    .A2(_04727_),
    .Y(_04754_),
    .B1(_04753_));
 sg13g2_inv_2 _12682_ (.Y(_04755_),
    .A(net1687));
 sg13g2_nor3_1 _12683_ (.A(_04664_),
    .B(_04666_),
    .C(_04727_),
    .Y(_04756_));
 sg13g2_xnor2_1 _12684_ (.Y(_04757_),
    .A(_04736_),
    .B(_04752_));
 sg13g2_nor3_1 _12685_ (.A(net1686),
    .B(_04756_),
    .C(_04757_),
    .Y(_04758_));
 sg13g2_a21oi_1 _12686_ (.A1(_04745_),
    .A2(net1686),
    .Y(_04759_),
    .B1(_04758_));
 sg13g2_nand2_1 _12687_ (.Y(_04760_),
    .A(net1690),
    .B(_04759_));
 sg13g2_nand3_1 _12688_ (.B(_04666_),
    .C(_04736_),
    .A(_04664_),
    .Y(_04761_));
 sg13g2_a21oi_1 _12689_ (.A1(_04734_),
    .A2(net1686),
    .Y(_04762_),
    .B1(net1694));
 sg13g2_nor2_1 _12690_ (.A(_04565_),
    .B(net1711),
    .Y(_04763_));
 sg13g2_a21oi_1 _12691_ (.A1(_04570_),
    .A2(net1710),
    .Y(_04764_),
    .B1(_04763_));
 sg13g2_nor2_1 _12692_ (.A(_04577_),
    .B(net1712),
    .Y(_04765_));
 sg13g2_a21oi_1 _12693_ (.A1(_04579_),
    .A2(net1713),
    .Y(_04766_),
    .B1(_04765_));
 sg13g2_nor2_1 _12694_ (.A(net1720),
    .B(_04766_),
    .Y(_04767_));
 sg13g2_a21oi_1 _12695_ (.A1(net1720),
    .A2(_04764_),
    .Y(_04768_),
    .B1(_04767_));
 sg13g2_nand2_1 _12696_ (.Y(_04769_),
    .A(_04560_),
    .B(net1712));
 sg13g2_o21ai_1 _12697_ (.B1(_04769_),
    .Y(_04770_),
    .A1(_04553_),
    .A2(net1712));
 sg13g2_nor2_1 _12698_ (.A(net1718),
    .B(_04770_),
    .Y(_04771_));
 sg13g2_a22oi_1 _12699_ (.Y(_04772_),
    .B1(_04546_),
    .B2(_04460_),
    .A2(_04544_),
    .A1(_04543_));
 sg13g2_nand2_1 _12700_ (.Y(_04773_),
    .A(net1719),
    .B(_04772_));
 sg13g2_nor2_1 _12701_ (.A(net1722),
    .B(_04771_),
    .Y(_04774_));
 sg13g2_nor2_1 _12702_ (.A(_04589_),
    .B(net1707),
    .Y(_04775_));
 sg13g2_a21oi_1 _12703_ (.A1(_04596_),
    .A2(net1708),
    .Y(_04776_),
    .B1(_04775_));
 sg13g2_mux2_1 _12704_ (.A0(_04604_),
    .A1(_04610_),
    .S(net1707),
    .X(_04777_));
 sg13g2_nor2_1 _12705_ (.A(net1720),
    .B(_04777_),
    .Y(_04778_));
 sg13g2_a21oi_1 _12706_ (.A1(net1720),
    .A2(_04776_),
    .Y(_04779_),
    .B1(_04778_));
 sg13g2_nand2_1 _12707_ (.Y(_04780_),
    .A(net1725),
    .B(_04779_));
 sg13g2_o21ai_1 _12708_ (.B1(_04780_),
    .Y(_04781_),
    .A1(net1725),
    .A2(_04661_));
 sg13g2_nor2b_1 _12709_ (.A(_04585_),
    .B_N(_04781_),
    .Y(_04782_));
 sg13g2_a221oi_1 _12710_ (.B2(_04774_),
    .C1(_04782_),
    .B1(_04773_),
    .A1(net1722),
    .Y(_04783_),
    .A2(_04768_));
 sg13g2_nand2b_2 _12711_ (.Y(_04784_),
    .B(_04783_),
    .A_N(_04652_));
 sg13g2_nor2_1 _12712_ (.A(_03444_),
    .B(_03448_),
    .Y(_04785_));
 sg13g2_nand4_1 _12713_ (.B(net1933),
    .C(_03433_),
    .A(_03308_),
    .Y(_04786_),
    .D(_03452_));
 sg13g2_inv_1 _12714_ (.Y(_04787_),
    .A(_04786_));
 sg13g2_nor2_1 _12715_ (.A(_04785_),
    .B(_04787_),
    .Y(_04788_));
 sg13g2_nand2_1 _12716_ (.Y(_04789_),
    .A(net1776),
    .B(_04788_));
 sg13g2_o21ai_1 _12717_ (.B1(_04302_),
    .Y(_04790_),
    .A1(_04784_),
    .A2(_04789_));
 sg13g2_a21oi_1 _12718_ (.A1(net1950),
    .A2(_04787_),
    .Y(_04791_),
    .B1(_03448_));
 sg13g2_nor2_1 _12719_ (.A(_03444_),
    .B(_04791_),
    .Y(_04792_));
 sg13g2_or2_1 _12720_ (.X(_04793_),
    .B(_04792_),
    .A(_03455_));
 sg13g2_or2_1 _12721_ (.X(_04794_),
    .B(_04793_),
    .A(net2197));
 sg13g2_inv_2 _12722_ (.Y(_04795_),
    .A(_04794_));
 sg13g2_nand2b_1 _12723_ (.Y(_04796_),
    .B(_04795_),
    .A_N(_04790_));
 sg13g2_a21oi_1 _12724_ (.A1(_04761_),
    .A2(_04762_),
    .Y(_04797_),
    .B1(net1683));
 sg13g2_a22oi_1 _12725_ (.Y(_04798_),
    .B1(_04760_),
    .B2(_04797_),
    .A2(net2201),
    .A1(net3485));
 sg13g2_inv_1 _12726_ (.Y(_00174_),
    .A(_04798_));
 sg13g2_nand2_1 _12727_ (.Y(_04799_),
    .A(net1708),
    .B(_04635_));
 sg13g2_o21ai_1 _12728_ (.B1(_04799_),
    .Y(_04800_),
    .A1(_04598_),
    .A2(net1708));
 sg13g2_nand2_1 _12729_ (.Y(_04801_),
    .A(net1716),
    .B(_04800_));
 sg13g2_nand3_1 _12730_ (.B(net1715),
    .C(_04800_),
    .A(net1725),
    .Y(_04802_));
 sg13g2_or3_1 _12731_ (.A(_04077_),
    .B(_04096_),
    .C(_04164_),
    .X(_04803_));
 sg13g2_nand2_1 _12732_ (.Y(_04804_),
    .A(_04165_),
    .B(_04803_));
 sg13g2_a21o_1 _12733_ (.A2(_04804_),
    .A1(net1946),
    .B1(net1705),
    .X(_04805_));
 sg13g2_a221oi_1 _12734_ (.B2(net1776),
    .C1(_04805_),
    .B1(_04802_),
    .A1(net1761),
    .Y(_04806_),
    .A2(_04742_));
 sg13g2_nor3_1 _12735_ (.A(_04667_),
    .B(_04709_),
    .C(_04723_),
    .Y(_04807_));
 sg13g2_nor2_1 _12736_ (.A(_04806_),
    .B(net1701),
    .Y(_04808_));
 sg13g2_or3_1 _12737_ (.A(_04736_),
    .B(_04752_),
    .C(_04808_),
    .X(_04809_));
 sg13g2_o21ai_1 _12738_ (.B1(_04808_),
    .Y(_04810_),
    .A1(_04736_),
    .A2(_04752_));
 sg13g2_and2_1 _12739_ (.A(_04809_),
    .B(_04810_),
    .X(_04811_));
 sg13g2_mux2_1 _12740_ (.A0(_04811_),
    .A1(_04806_),
    .S(net1686),
    .X(_04812_));
 sg13g2_or2_1 _12741_ (.X(_04813_),
    .B(_04812_),
    .A(net1695));
 sg13g2_a21oi_1 _12742_ (.A1(net1695),
    .A2(_04759_),
    .Y(_04814_),
    .B1(net1682));
 sg13g2_a22oi_1 _12743_ (.Y(_04815_),
    .B1(_04813_),
    .B2(_04814_),
    .A2(net2201),
    .A1(net3601));
 sg13g2_inv_1 _12744_ (.Y(_00175_),
    .A(_04815_));
 sg13g2_or2_1 _12745_ (.X(_04816_),
    .B(net1702),
    .A(_04715_));
 sg13g2_nor2_1 _12746_ (.A(_04746_),
    .B(_04816_),
    .Y(_04817_));
 sg13g2_inv_1 _12747_ (.Y(_04818_),
    .A(_04817_));
 sg13g2_nor2_1 _12748_ (.A(net1715),
    .B(_04660_),
    .Y(_04819_));
 sg13g2_a21oi_2 _12749_ (.B1(_04819_),
    .Y(_04820_),
    .A2(_04776_),
    .A1(net1715));
 sg13g2_a21o_1 _12750_ (.A2(_04820_),
    .A1(net1725),
    .B1(net1773),
    .X(_04821_));
 sg13g2_nand3_1 _12751_ (.B(_04165_),
    .C(_04167_),
    .A(_04076_),
    .Y(_04822_));
 sg13g2_and2_1 _12752_ (.A(_04168_),
    .B(_04822_),
    .X(_04823_));
 sg13g2_nor2_1 _12753_ (.A(net1950),
    .B(_04823_),
    .Y(_04824_));
 sg13g2_a21oi_1 _12754_ (.A1(net1761),
    .A2(_04804_),
    .Y(_04825_),
    .B1(_04824_));
 sg13g2_nand3_1 _12755_ (.B(_04821_),
    .C(_04825_),
    .A(net1703),
    .Y(_04826_));
 sg13g2_xnor2_1 _12756_ (.Y(_04827_),
    .A(_04704_),
    .B(_04706_));
 sg13g2_and3_2 _12757_ (.X(_04828_),
    .A(_04711_),
    .B(_04713_),
    .C(_04827_));
 sg13g2_nand3_1 _12758_ (.B(_04713_),
    .C(_04827_),
    .A(_04711_),
    .Y(_04829_));
 sg13g2_nor2_2 _12759_ (.A(_04719_),
    .B(_04829_),
    .Y(_04830_));
 sg13g2_nand4_1 _12760_ (.B(_04713_),
    .C(_04720_),
    .A(_04711_),
    .Y(_04831_),
    .D(_04827_));
 sg13g2_and2_1 _12761_ (.A(net1700),
    .B(_04831_),
    .X(_04832_));
 sg13g2_nand2_2 _12762_ (.Y(_04833_),
    .A(net1700),
    .B(_04831_));
 sg13g2_o21ai_1 _12763_ (.B1(net1701),
    .Y(_04834_),
    .A1(_04818_),
    .A2(_04831_));
 sg13g2_and3_1 _12764_ (.X(_04835_),
    .A(_04809_),
    .B(_04826_),
    .C(_04834_));
 sg13g2_a21o_1 _12765_ (.A2(_04834_),
    .A1(_04826_),
    .B1(_04808_),
    .X(_04836_));
 sg13g2_nor3_1 _12766_ (.A(_04736_),
    .B(_04752_),
    .C(_04836_),
    .Y(_04837_));
 sg13g2_nand2_1 _12767_ (.Y(_04838_),
    .A(net1686),
    .B(_04826_));
 sg13g2_o21ai_1 _12768_ (.B1(_04755_),
    .Y(_04839_),
    .A1(_04835_),
    .A2(_04837_));
 sg13g2_a21oi_1 _12769_ (.A1(_04838_),
    .A2(_04839_),
    .Y(_04840_),
    .B1(net1695));
 sg13g2_nor2_1 _12770_ (.A(net1682),
    .B(_04840_),
    .Y(_04841_));
 sg13g2_o21ai_1 _12771_ (.B1(_04841_),
    .Y(_04842_),
    .A1(net1690),
    .A2(_04812_));
 sg13g2_o21ai_1 _12772_ (.B1(_04842_),
    .Y(_00176_),
    .A1(_01139_),
    .A2(_03108_));
 sg13g2_nand2_1 _12773_ (.Y(_04843_),
    .A(net1715),
    .B(_04631_));
 sg13g2_o21ai_1 _12774_ (.B1(_04843_),
    .Y(_04844_),
    .A1(net1715),
    .A2(_04636_));
 sg13g2_o21ai_1 _12775_ (.B1(net1774),
    .Y(_04845_),
    .A1(net1721),
    .A2(_04844_));
 sg13g2_nand2b_1 _12776_ (.Y(_04846_),
    .B(net1761),
    .A_N(_04823_));
 sg13g2_nand3_1 _12777_ (.B(_04168_),
    .C(_04170_),
    .A(_04055_),
    .Y(_04847_));
 sg13g2_nand2_1 _12778_ (.Y(_04848_),
    .A(_04171_),
    .B(_04847_));
 sg13g2_a21oi_1 _12779_ (.A1(net1944),
    .A2(_04848_),
    .Y(_04849_),
    .B1(net1705));
 sg13g2_and3_1 _12780_ (.X(_04850_),
    .A(_04845_),
    .B(_04846_),
    .C(_04849_));
 sg13g2_inv_1 _12781_ (.Y(_04851_),
    .A(_04850_));
 sg13g2_nand2_1 _12782_ (.Y(_04852_),
    .A(_04711_),
    .B(_04827_));
 sg13g2_nand2_2 _12783_ (.Y(_04853_),
    .A(net1699),
    .B(_04852_));
 sg13g2_nand2_2 _12784_ (.Y(_04854_),
    .A(net1699),
    .B(_04829_));
 sg13g2_nand2b_2 _12785_ (.Y(_04855_),
    .B(_04720_),
    .A_N(net1702));
 sg13g2_o21ai_1 _12786_ (.B1(net1699),
    .Y(_04856_),
    .A1(_04715_),
    .A2(_04855_));
 sg13g2_and3_1 _12787_ (.X(_04857_),
    .A(_04851_),
    .B(_04854_),
    .C(_04856_));
 sg13g2_nor4_1 _12788_ (.A(_04736_),
    .B(_04752_),
    .C(_04836_),
    .D(_04857_),
    .Y(_04858_));
 sg13g2_xnor2_1 _12789_ (.Y(_04859_),
    .A(_04837_),
    .B(_04857_));
 sg13g2_nor2_1 _12790_ (.A(net1686),
    .B(_04859_),
    .Y(_04860_));
 sg13g2_a21oi_1 _12791_ (.A1(net1686),
    .A2(_04851_),
    .Y(_04861_),
    .B1(_04860_));
 sg13g2_nor2_1 _12792_ (.A(net1695),
    .B(_04861_),
    .Y(_04862_));
 sg13g2_a21oi_1 _12793_ (.A1(_04838_),
    .A2(_04839_),
    .Y(_04863_),
    .B1(net1690));
 sg13g2_nor3_1 _12794_ (.A(net1682),
    .B(_04862_),
    .C(_04863_),
    .Y(_04864_));
 sg13g2_a21o_1 _12795_ (.A2(net2201),
    .A1(net3649),
    .B1(_04864_),
    .X(_00177_));
 sg13g2_nor2_1 _12796_ (.A(_04610_),
    .B(net1707),
    .Y(_04865_));
 sg13g2_a21oi_1 _12797_ (.A1(_04589_),
    .A2(net1707),
    .Y(_04866_),
    .B1(_04865_));
 sg13g2_mux2_1 _12798_ (.A0(_04738_),
    .A1(_04866_),
    .S(net1715),
    .X(_04867_));
 sg13g2_nand2_1 _12799_ (.Y(_04868_),
    .A(net1725),
    .B(_04867_));
 sg13g2_nand3_1 _12800_ (.B(_04171_),
    .C(_04173_),
    .A(_04037_),
    .Y(_04869_));
 sg13g2_nand2b_2 _12801_ (.Y(_04870_),
    .B(_04869_),
    .A_N(_04174_));
 sg13g2_nand2_1 _12802_ (.Y(_04871_),
    .A(net1944),
    .B(_04870_));
 sg13g2_a221oi_1 _12803_ (.B2(net1774),
    .C1(net1705),
    .B1(_04868_),
    .A1(net1762),
    .Y(_04872_),
    .A2(_04848_));
 sg13g2_and2_1 _12804_ (.A(_04871_),
    .B(_04872_),
    .X(_04873_));
 sg13g2_nor2_1 _12805_ (.A(_04748_),
    .B(_04855_),
    .Y(_04874_));
 sg13g2_nand2_1 _12806_ (.Y(_04875_),
    .A(_04828_),
    .B(_04874_));
 sg13g2_a21o_2 _12807_ (.A2(_04875_),
    .A1(net1700),
    .B1(_04873_),
    .X(_04876_));
 sg13g2_nand2_1 _12808_ (.Y(_04877_),
    .A(_04858_),
    .B(_04876_));
 sg13g2_xnor2_1 _12809_ (.Y(_04878_),
    .A(_04858_),
    .B(_04876_));
 sg13g2_nand2_1 _12810_ (.Y(_04879_),
    .A(net1686),
    .B(_04873_));
 sg13g2_o21ai_1 _12811_ (.B1(_04879_),
    .Y(_04880_),
    .A1(net1689),
    .A2(_04878_));
 sg13g2_inv_1 _12812_ (.Y(_04881_),
    .A(_04880_));
 sg13g2_a21oi_1 _12813_ (.A1(net1690),
    .A2(_04881_),
    .Y(_04882_),
    .B1(net1682));
 sg13g2_o21ai_1 _12814_ (.B1(_04882_),
    .Y(_04883_),
    .A1(net1690),
    .A2(_04861_));
 sg13g2_o21ai_1 _12815_ (.B1(_04883_),
    .Y(_00178_),
    .A1(_01141_),
    .A2(_03108_));
 sg13g2_or2_1 _12816_ (.X(_04884_),
    .B(_04800_),
    .A(net1716));
 sg13g2_nand2_1 _12817_ (.Y(_04885_),
    .A(_04593_),
    .B(net1707));
 sg13g2_o21ai_1 _12818_ (.B1(_04885_),
    .Y(_04886_),
    .A1(_04612_),
    .A2(net1710));
 sg13g2_o21ai_1 _12819_ (.B1(_04884_),
    .Y(_04887_),
    .A1(net1720),
    .A2(_04886_));
 sg13g2_nand2b_1 _12820_ (.Y(_04888_),
    .B(net1726),
    .A_N(_04887_));
 sg13g2_nor2_1 _12821_ (.A(_03998_),
    .B(_03999_),
    .Y(_04889_));
 sg13g2_xor2_1 _12822_ (.B(_04889_),
    .A(_04175_),
    .X(_04890_));
 sg13g2_a22oi_1 _12823_ (.Y(_04891_),
    .B1(_04890_),
    .B2(net1944),
    .A2(_04870_),
    .A1(net1761));
 sg13g2_nand2_1 _12824_ (.Y(_04892_),
    .A(net1703),
    .B(_04891_));
 sg13g2_a21oi_1 _12825_ (.A1(net1775),
    .A2(_04888_),
    .Y(_04893_),
    .B1(_04892_));
 sg13g2_a21oi_1 _12826_ (.A1(net1699),
    .A2(_04855_),
    .Y(_04894_),
    .B1(_04893_));
 sg13g2_and2_1 _12827_ (.A(_04854_),
    .B(_04894_),
    .X(_04895_));
 sg13g2_nand2_1 _12828_ (.Y(_04896_),
    .A(_04854_),
    .B(_04894_));
 sg13g2_nor2_1 _12829_ (.A(_04877_),
    .B(_04895_),
    .Y(_04897_));
 sg13g2_xnor2_1 _12830_ (.Y(_04898_),
    .A(_04877_),
    .B(_04895_));
 sg13g2_nand2_1 _12831_ (.Y(_04899_),
    .A(net1687),
    .B(_04893_));
 sg13g2_o21ai_1 _12832_ (.B1(_04899_),
    .Y(_04900_),
    .A1(net1689),
    .A2(_04898_));
 sg13g2_nor2_1 _12833_ (.A(net1695),
    .B(_04900_),
    .Y(_04901_));
 sg13g2_nor2_1 _12834_ (.A(net1690),
    .B(_04880_),
    .Y(_04902_));
 sg13g2_nor3_1 _12835_ (.A(net1682),
    .B(_04901_),
    .C(_04902_),
    .Y(_04903_));
 sg13g2_a21o_1 _12836_ (.A2(net2201),
    .A1(net3602),
    .B1(_04903_),
    .X(_00179_));
 sg13g2_xnor2_1 _12837_ (.Y(_04904_),
    .A(_04177_),
    .B(_04179_));
 sg13g2_a22oi_1 _12838_ (.Y(_04905_),
    .B1(_04904_),
    .B2(net1944),
    .A2(_04781_),
    .A1(net1774));
 sg13g2_o21ai_1 _12839_ (.B1(_04905_),
    .Y(_04906_),
    .A1(_04677_),
    .A2(_04890_));
 sg13g2_nand2_1 _12840_ (.Y(_04907_),
    .A(net1703),
    .B(_04906_));
 sg13g2_nor2_1 _12841_ (.A(net1702),
    .B(_04829_),
    .Y(_04908_));
 sg13g2_o21ai_1 _12842_ (.B1(net1702),
    .Y(_04909_),
    .A1(_04715_),
    .A2(_04746_));
 sg13g2_nand2_1 _12843_ (.Y(_04910_),
    .A(_04828_),
    .B(_04909_));
 sg13g2_o21ai_1 _12844_ (.B1(net1700),
    .Y(_04911_),
    .A1(_04719_),
    .A2(_04910_));
 sg13g2_nand2_1 _12845_ (.Y(_04912_),
    .A(_04907_),
    .B(_04911_));
 sg13g2_nand4_1 _12846_ (.B(_04876_),
    .C(_04896_),
    .A(_04858_),
    .Y(_04913_),
    .D(_04912_));
 sg13g2_xnor2_1 _12847_ (.Y(_04914_),
    .A(_04897_),
    .B(_04912_));
 sg13g2_mux2_1 _12848_ (.A0(_04907_),
    .A1(_04914_),
    .S(_04755_),
    .X(_04915_));
 sg13g2_a21oi_1 _12849_ (.A1(net1691),
    .A2(_04915_),
    .Y(_04916_),
    .B1(net1682));
 sg13g2_o21ai_1 _12850_ (.B1(_04916_),
    .Y(_04917_),
    .A1(net1690),
    .A2(_04900_));
 sg13g2_o21ai_1 _12851_ (.B1(_04917_),
    .Y(_00180_),
    .A1(_01143_),
    .A2(_03108_));
 sg13g2_xor2_1 _12852_ (.B(_04181_),
    .A(_03948_),
    .X(_04918_));
 sg13g2_a22oi_1 _12853_ (.Y(_04919_),
    .B1(net1763),
    .B2(_04904_),
    .A2(_04640_),
    .A1(net1774));
 sg13g2_o21ai_1 _12854_ (.B1(_04919_),
    .Y(_04920_),
    .A1(net1949),
    .A2(_04918_));
 sg13g2_nand2_1 _12855_ (.Y(_04921_),
    .A(_04717_),
    .B(_04720_));
 sg13g2_nand2_1 _12856_ (.Y(_04922_),
    .A(_04717_),
    .B(_04830_));
 sg13g2_a22oi_1 _12857_ (.Y(_04923_),
    .B1(_04922_),
    .B2(net1699),
    .A2(_04920_),
    .A1(net1703));
 sg13g2_nor2_1 _12858_ (.A(_04913_),
    .B(_04923_),
    .Y(_04924_));
 sg13g2_xor2_1 _12859_ (.B(_04923_),
    .A(_04913_),
    .X(_04925_));
 sg13g2_a21o_1 _12860_ (.A2(_04920_),
    .A1(net1704),
    .B1(_04755_),
    .X(_04926_));
 sg13g2_o21ai_1 _12861_ (.B1(_04926_),
    .Y(_04927_),
    .A1(net1688),
    .A2(_04925_));
 sg13g2_nand2_1 _12862_ (.Y(_04928_),
    .A(net1695),
    .B(_04915_));
 sg13g2_a21oi_1 _12863_ (.A1(net1693),
    .A2(_04927_),
    .Y(_04929_),
    .B1(net1685));
 sg13g2_a22oi_1 _12864_ (.Y(_04930_),
    .B1(_04928_),
    .B2(_04929_),
    .A2(net2199),
    .A1(net3811));
 sg13g2_inv_1 _12865_ (.Y(_00181_),
    .A(_04930_));
 sg13g2_nor2_1 _12866_ (.A(net1773),
    .B(net1721),
    .Y(_04931_));
 sg13g2_nand2_1 _12867_ (.Y(_04932_),
    .A(_04605_),
    .B(net1710));
 sg13g2_o21ai_1 _12868_ (.B1(_04932_),
    .Y(_04933_),
    .A1(_04570_),
    .A2(net1710));
 sg13g2_nand2_1 _12869_ (.Y(_04934_),
    .A(net1717),
    .B(_04933_));
 sg13g2_o21ai_1 _12870_ (.B1(_04934_),
    .Y(_04935_),
    .A1(net1716),
    .A2(_04866_));
 sg13g2_inv_1 _12871_ (.Y(_04936_),
    .A(_04935_));
 sg13g2_nand2b_1 _12872_ (.Y(_04937_),
    .B(_04185_),
    .A_N(_04192_));
 sg13g2_xnor2_1 _12873_ (.Y(_04938_),
    .A(_04185_),
    .B(_04192_));
 sg13g2_a21oi_1 _12874_ (.A1(net1761),
    .A2(_04918_),
    .Y(_04939_),
    .B1(net1705));
 sg13g2_o21ai_1 _12875_ (.B1(_04939_),
    .Y(_04940_),
    .A1(net1949),
    .A2(_04938_));
 sg13g2_a221oi_1 _12876_ (.B2(_04935_),
    .C1(_04940_),
    .B1(_04931_),
    .A1(net1706),
    .Y(_04941_),
    .A2(_04739_));
 sg13g2_and3_1 _12877_ (.X(_04942_),
    .A(net1702),
    .B(_04748_),
    .C(net1700));
 sg13g2_nor3_1 _12878_ (.A(_04832_),
    .B(_04941_),
    .C(_04942_),
    .Y(_04943_));
 sg13g2_nor2b_1 _12879_ (.A(_04924_),
    .B_N(_04943_),
    .Y(_04944_));
 sg13g2_nand2b_1 _12880_ (.Y(_04945_),
    .B(_04924_),
    .A_N(_04943_));
 sg13g2_nor2_1 _12881_ (.A(net1687),
    .B(_04944_),
    .Y(_04946_));
 sg13g2_a22oi_1 _12882_ (.Y(_04947_),
    .B1(_04945_),
    .B2(_04946_),
    .A2(_04941_),
    .A1(net1688));
 sg13g2_nand2_1 _12883_ (.Y(_04948_),
    .A(net1692),
    .B(_04947_));
 sg13g2_a21oi_1 _12884_ (.A1(net1697),
    .A2(_04927_),
    .Y(_04949_),
    .B1(net1685));
 sg13g2_a22oi_1 _12885_ (.Y(_04950_),
    .B1(_04948_),
    .B2(_04949_),
    .A2(net2199),
    .A1(net3861));
 sg13g2_inv_1 _12886_ (.Y(_00182_),
    .A(_04950_));
 sg13g2_nand2_1 _12887_ (.Y(_04951_),
    .A(_04602_),
    .B(net1710));
 sg13g2_o21ai_1 _12888_ (.B1(_04951_),
    .Y(_04952_),
    .A1(_04568_),
    .A2(net1710));
 sg13g2_nand2_1 _12889_ (.Y(_04953_),
    .A(net1717),
    .B(_04952_));
 sg13g2_o21ai_1 _12890_ (.B1(_04953_),
    .Y(_04954_),
    .A1(net1717),
    .A2(_04886_));
 sg13g2_a21oi_1 _12891_ (.A1(net1725),
    .A2(_04954_),
    .Y(_04955_),
    .B1(_04659_));
 sg13g2_and2_1 _12892_ (.A(_04191_),
    .B(_04937_),
    .X(_04956_));
 sg13g2_xor2_1 _12893_ (.B(_04956_),
    .A(_04200_),
    .X(_04957_));
 sg13g2_a221oi_1 _12894_ (.B2(net1944),
    .C1(_04955_),
    .B1(_04957_),
    .A1(net1762),
    .Y(_04958_),
    .A2(_04938_));
 sg13g2_a21o_1 _12895_ (.A2(_04801_),
    .A1(net1706),
    .B1(_04958_),
    .X(_04959_));
 sg13g2_and2_1 _12896_ (.A(_04833_),
    .B(_04959_),
    .X(_04960_));
 sg13g2_or4_1 _12897_ (.A(_04913_),
    .B(_04923_),
    .C(_04943_),
    .D(_04960_),
    .X(_04961_));
 sg13g2_nor2_1 _12898_ (.A(net1688),
    .B(_04961_),
    .Y(_04962_));
 sg13g2_a22oi_1 _12899_ (.Y(_04963_),
    .B1(_04960_),
    .B2(_04945_),
    .A2(_04959_),
    .A1(net1687));
 sg13g2_nand2b_1 _12900_ (.Y(_04964_),
    .B(_04963_),
    .A_N(_04962_));
 sg13g2_a21o_1 _12901_ (.A2(_04947_),
    .A1(net1697),
    .B1(net1684),
    .X(_04965_));
 sg13g2_a21oi_1 _12902_ (.A1(net1693),
    .A2(_04964_),
    .Y(_04966_),
    .B1(_04965_));
 sg13g2_a21o_1 _12903_ (.A2(net2199),
    .A1(net3750),
    .B1(_04966_),
    .X(_00183_));
 sg13g2_nand2_1 _12904_ (.Y(_04967_),
    .A(_04212_),
    .B(_04218_));
 sg13g2_o21ai_1 _12905_ (.B1(_04199_),
    .Y(_04968_),
    .A1(_04200_),
    .A2(_04956_));
 sg13g2_xnor2_1 _12906_ (.Y(_04969_),
    .A(_04967_),
    .B(_04968_));
 sg13g2_nor2_1 _12907_ (.A(net1717),
    .B(_04777_),
    .Y(_04970_));
 sg13g2_a21oi_1 _12908_ (.A1(net1717),
    .A2(_04764_),
    .Y(_04971_),
    .B1(_04970_));
 sg13g2_a22oi_1 _12909_ (.Y(_04972_),
    .B1(_04971_),
    .B2(_04931_),
    .A2(_04957_),
    .A1(net1762));
 sg13g2_nand2_1 _12910_ (.Y(_04973_),
    .A(net1706),
    .B(_04820_));
 sg13g2_nand2_1 _12911_ (.Y(_04974_),
    .A(_04972_),
    .B(_04973_));
 sg13g2_a21oi_1 _12912_ (.A1(net1944),
    .A2(_04969_),
    .Y(_04975_),
    .B1(_04974_));
 sg13g2_a21oi_1 _12913_ (.A1(_04817_),
    .A2(_04828_),
    .Y(_04976_),
    .B1(_04833_));
 sg13g2_nor2b_2 _12914_ (.A(_04976_),
    .B_N(_04975_),
    .Y(_04977_));
 sg13g2_xor2_1 _12915_ (.B(_04975_),
    .A(_04962_),
    .X(_04978_));
 sg13g2_nand2_1 _12916_ (.Y(_04979_),
    .A(net1693),
    .B(_04978_));
 sg13g2_a21oi_1 _12917_ (.A1(net1697),
    .A2(_04964_),
    .Y(_04980_),
    .B1(net1684));
 sg13g2_a22oi_1 _12918_ (.Y(_04981_),
    .B1(_04979_),
    .B2(_04980_),
    .A2(net2199),
    .A1(net3810));
 sg13g2_inv_1 _12919_ (.Y(_00184_),
    .A(_04981_));
 sg13g2_and2_1 _12920_ (.A(net4084),
    .B(net2199),
    .X(_04982_));
 sg13g2_nand2_1 _12921_ (.Y(_04983_),
    .A(net1706),
    .B(_04844_));
 sg13g2_nand2b_1 _12922_ (.Y(_04984_),
    .B(_04214_),
    .A_N(_04207_));
 sg13g2_a21oi_1 _12923_ (.A1(_04218_),
    .A2(_04968_),
    .Y(_04985_),
    .B1(_04213_));
 sg13g2_xnor2_1 _12924_ (.Y(_04986_),
    .A(_04984_),
    .B(_04985_));
 sg13g2_mux2_1 _12925_ (.A0(_04633_),
    .A1(_04642_),
    .S(net1719),
    .X(_04987_));
 sg13g2_a21oi_1 _12926_ (.A1(net1725),
    .A2(_04987_),
    .Y(_04988_),
    .B1(_04659_));
 sg13g2_a21oi_1 _12927_ (.A1(net1762),
    .A2(_04969_),
    .Y(_04989_),
    .B1(_04988_));
 sg13g2_o21ai_1 _12928_ (.B1(_04989_),
    .Y(_04990_),
    .A1(net1949),
    .A2(_04986_));
 sg13g2_nand2_1 _12929_ (.Y(_04991_),
    .A(_04983_),
    .B(_04990_));
 sg13g2_o21ai_1 _12930_ (.B1(_04832_),
    .Y(_04992_),
    .A1(_04816_),
    .A2(_04829_));
 sg13g2_and2_1 _12931_ (.A(_04991_),
    .B(_04992_),
    .X(_04993_));
 sg13g2_nor4_1 _12932_ (.A(net1687),
    .B(_04961_),
    .C(_04977_),
    .D(_04993_),
    .Y(_04994_));
 sg13g2_inv_1 _12933_ (.Y(_04995_),
    .A(_04994_));
 sg13g2_o21ai_1 _12934_ (.B1(_04993_),
    .Y(_04996_),
    .A1(_04961_),
    .A2(_04977_));
 sg13g2_a21oi_1 _12935_ (.A1(net1688),
    .A2(_04991_),
    .Y(_04997_),
    .B1(_04994_));
 sg13g2_nand2_1 _12936_ (.Y(_04998_),
    .A(_04996_),
    .B(_04997_));
 sg13g2_nand2_1 _12937_ (.Y(_04999_),
    .A(net1697),
    .B(_04978_));
 sg13g2_a21oi_1 _12938_ (.A1(net1691),
    .A2(_04998_),
    .Y(_05000_),
    .B1(net1683));
 sg13g2_a21o_1 _12939_ (.A2(_05000_),
    .A1(_04999_),
    .B1(_04982_),
    .X(_00185_));
 sg13g2_nor2_1 _12940_ (.A(_04677_),
    .B(_04986_),
    .Y(_05001_));
 sg13g2_mux2_1 _12941_ (.A0(_04579_),
    .A1(_04565_),
    .S(net1711),
    .X(_05002_));
 sg13g2_mux2_1 _12942_ (.A0(_04933_),
    .A1(_05002_),
    .S(net1717),
    .X(_05003_));
 sg13g2_nor3_1 _12943_ (.A(_04311_),
    .B(net1721),
    .C(_05003_),
    .Y(_05004_));
 sg13g2_nand2_1 _12944_ (.Y(_05005_),
    .A(net1706),
    .B(_04867_));
 sg13g2_nand2_1 _12945_ (.Y(_05006_),
    .A(_04220_),
    .B(_04242_));
 sg13g2_xnor2_1 _12946_ (.Y(_05007_),
    .A(_04220_),
    .B(_04242_));
 sg13g2_o21ai_1 _12947_ (.B1(_05005_),
    .Y(_05008_),
    .A1(net1949),
    .A2(_05007_));
 sg13g2_nor3_1 _12948_ (.A(_05001_),
    .B(_05004_),
    .C(_05008_),
    .Y(_05009_));
 sg13g2_nand2_1 _12949_ (.Y(_05010_),
    .A(_04995_),
    .B(_05009_));
 sg13g2_nor3_1 _12950_ (.A(net1702),
    .B(_04748_),
    .C(_04829_),
    .Y(_05011_));
 sg13g2_o21ai_1 _12951_ (.B1(_05009_),
    .Y(_05012_),
    .A1(_04833_),
    .A2(_05011_));
 sg13g2_nand2_1 _12952_ (.Y(_05013_),
    .A(_04994_),
    .B(_05012_));
 sg13g2_nand2_1 _12953_ (.Y(_05014_),
    .A(_05010_),
    .B(_05013_));
 sg13g2_nand2_1 _12954_ (.Y(_05015_),
    .A(net1695),
    .B(_04998_));
 sg13g2_a21oi_1 _12955_ (.A1(net1691),
    .A2(_05014_),
    .Y(_05016_),
    .B1(net1682));
 sg13g2_a22oi_1 _12956_ (.Y(_05017_),
    .B1(_05015_),
    .B2(_05016_),
    .A2(net2201),
    .A1(net3985));
 sg13g2_inv_1 _12957_ (.Y(_00186_),
    .A(_05017_));
 sg13g2_and2_1 _12958_ (.A(net4080),
    .B(net2201),
    .X(_05018_));
 sg13g2_nand2_1 _12959_ (.Y(_05019_),
    .A(_04663_),
    .B(_04887_));
 sg13g2_a21oi_1 _12960_ (.A1(_04220_),
    .A2(_04242_),
    .Y(_05020_),
    .B1(_04241_));
 sg13g2_xnor2_1 _12961_ (.Y(_05021_),
    .A(_04249_),
    .B(_05020_));
 sg13g2_nor2_1 _12962_ (.A(net1949),
    .B(_05021_),
    .Y(_05022_));
 sg13g2_mux2_1 _12963_ (.A0(_04581_),
    .A1(_04563_),
    .S(net1714),
    .X(_05023_));
 sg13g2_or2_1 _12964_ (.X(_05024_),
    .B(_05023_),
    .A(net1720));
 sg13g2_o21ai_1 _12965_ (.B1(_05024_),
    .Y(_05025_),
    .A1(net1718),
    .A2(_04952_));
 sg13g2_o21ai_1 _12966_ (.B1(_04658_),
    .Y(_05026_),
    .A1(net1722),
    .A2(_05025_));
 sg13g2_o21ai_1 _12967_ (.B1(_05026_),
    .Y(_05027_),
    .A1(_04677_),
    .A2(_05007_));
 sg13g2_o21ai_1 _12968_ (.B1(_05019_),
    .Y(_05028_),
    .A1(_05022_),
    .A2(_05027_));
 sg13g2_o21ai_1 _12969_ (.B1(_05028_),
    .Y(_05029_),
    .A1(_04833_),
    .A2(_04908_));
 sg13g2_nand2_1 _12970_ (.Y(_05030_),
    .A(_05012_),
    .B(_05029_));
 sg13g2_nor2_1 _12971_ (.A(_04995_),
    .B(_05030_),
    .Y(_05031_));
 sg13g2_a21o_1 _12972_ (.A2(_05028_),
    .A1(_05013_),
    .B1(_05031_),
    .X(_05032_));
 sg13g2_nand2_1 _12973_ (.Y(_05033_),
    .A(net1696),
    .B(_05014_));
 sg13g2_a21oi_1 _12974_ (.A1(net1691),
    .A2(_05032_),
    .Y(_05034_),
    .B1(net1682));
 sg13g2_a21o_1 _12975_ (.A2(_05034_),
    .A1(_05033_),
    .B1(_05018_),
    .X(_00187_));
 sg13g2_nor2_1 _12976_ (.A(_04249_),
    .B(_05006_),
    .Y(_05035_));
 sg13g2_nor2b_1 _12977_ (.A(_05035_),
    .B_N(_04253_),
    .Y(_05036_));
 sg13g2_xnor2_1 _12978_ (.Y(_05037_),
    .A(_04227_),
    .B(_05036_));
 sg13g2_a21o_1 _12979_ (.A2(_04768_),
    .A1(net1726),
    .B1(_04659_),
    .X(_05038_));
 sg13g2_a21oi_1 _12980_ (.A1(net1721),
    .A2(_04779_),
    .Y(_05039_),
    .B1(_05038_));
 sg13g2_a221oi_1 _12981_ (.B2(net1944),
    .C1(_05039_),
    .B1(_05037_),
    .A1(net1762),
    .Y(_05040_),
    .A2(_05021_));
 sg13g2_o21ai_1 _12982_ (.B1(_05040_),
    .Y(_05041_),
    .A1(_04662_),
    .A2(net1703));
 sg13g2_inv_1 _12983_ (.Y(_05042_),
    .A(_05041_));
 sg13g2_a21oi_1 _12984_ (.A1(_04832_),
    .A2(_04910_),
    .Y(_05043_),
    .B1(_05042_));
 sg13g2_or3_1 _12985_ (.A(_04995_),
    .B(_05030_),
    .C(_05043_),
    .X(_05044_));
 sg13g2_o21ai_1 _12986_ (.B1(_05044_),
    .Y(_05045_),
    .A1(_05031_),
    .A2(_05042_));
 sg13g2_nand2_1 _12987_ (.Y(_05046_),
    .A(net1695),
    .B(_05032_));
 sg13g2_a21oi_1 _12988_ (.A1(net1690),
    .A2(_05045_),
    .Y(_05047_),
    .B1(_04794_));
 sg13g2_a22oi_1 _12989_ (.Y(_05048_),
    .B1(_05046_),
    .B2(_05047_),
    .A2(net2201),
    .A1(net4032));
 sg13g2_inv_1 _12990_ (.Y(_00188_),
    .A(_05048_));
 sg13g2_o21ai_1 _12991_ (.B1(_04226_),
    .Y(_05049_),
    .A1(_04227_),
    .A2(_05036_));
 sg13g2_xor2_1 _12992_ (.B(_05049_),
    .A(_04234_),
    .X(_05050_));
 sg13g2_nand2_1 _12993_ (.Y(_05051_),
    .A(net1762),
    .B(_05037_));
 sg13g2_nor2_1 _12994_ (.A(net1722),
    .B(_04645_),
    .Y(_05052_));
 sg13g2_a21oi_1 _12995_ (.A1(net1723),
    .A2(_04634_),
    .Y(_05053_),
    .B1(_05052_));
 sg13g2_o21ai_1 _12996_ (.B1(_05051_),
    .Y(_05054_),
    .A1(net1703),
    .A2(_04728_));
 sg13g2_a221oi_1 _12997_ (.B2(_04658_),
    .C1(_05054_),
    .B1(_05053_),
    .A1(net1945),
    .Y(_05055_),
    .A2(_05050_));
 sg13g2_nand2_1 _12998_ (.Y(_05056_),
    .A(_04721_),
    .B(_04828_));
 sg13g2_a21oi_1 _12999_ (.A1(net1700),
    .A2(_05056_),
    .Y(_05057_),
    .B1(_05055_));
 sg13g2_or3_1 _13000_ (.A(_05030_),
    .B(_05043_),
    .C(_05057_),
    .X(_05058_));
 sg13g2_nor4_1 _13001_ (.A(_04961_),
    .B(_04977_),
    .C(_04993_),
    .D(_05058_),
    .Y(_05059_));
 sg13g2_or4_1 _13002_ (.A(_04961_),
    .B(_04977_),
    .C(_04993_),
    .D(_05058_),
    .X(_05060_));
 sg13g2_xor2_1 _13003_ (.B(_05055_),
    .A(_05044_),
    .X(_05061_));
 sg13g2_a21o_1 _13004_ (.A2(_05061_),
    .A1(net1691),
    .B1(net1683),
    .X(_05062_));
 sg13g2_a21oi_1 _13005_ (.A1(net1696),
    .A2(_05045_),
    .Y(_05063_),
    .B1(_05062_));
 sg13g2_a21o_1 _13006_ (.A2(net2201),
    .A1(net3774),
    .B1(_05063_),
    .X(_00189_));
 sg13g2_nor2_1 _13007_ (.A(_04677_),
    .B(_05050_),
    .Y(_05064_));
 sg13g2_nand2_1 _13008_ (.Y(_05065_),
    .A(net1705),
    .B(_04740_));
 sg13g2_xnor2_1 _13009_ (.Y(_05066_),
    .A(_04256_),
    .B(_04278_));
 sg13g2_nor2_1 _13010_ (.A(net1949),
    .B(_05066_),
    .Y(_05067_));
 sg13g2_mux2_1 _13011_ (.A0(_04560_),
    .A1(_04577_),
    .S(net1712),
    .X(_05068_));
 sg13g2_nand2_1 _13012_ (.Y(_05069_),
    .A(_04622_),
    .B(_05002_));
 sg13g2_nand2b_1 _13013_ (.Y(_05070_),
    .B(net1718),
    .A_N(_05068_));
 sg13g2_a22oi_1 _13014_ (.Y(_05071_),
    .B1(_05069_),
    .B2(_05070_),
    .A2(_04936_),
    .A1(net1722));
 sg13g2_o21ai_1 _13015_ (.B1(_05065_),
    .Y(_05072_),
    .A1(_04659_),
    .A2(_05071_));
 sg13g2_nor3_1 _13016_ (.A(_05064_),
    .B(_05067_),
    .C(_05072_),
    .Y(_05073_));
 sg13g2_nand2b_1 _13017_ (.Y(_05074_),
    .B(net1699),
    .A_N(_04749_));
 sg13g2_nand3_1 _13018_ (.B(_05073_),
    .C(_05074_),
    .A(_04854_),
    .Y(_05075_));
 sg13g2_inv_1 _13019_ (.Y(_05076_),
    .A(_05075_));
 sg13g2_nor3_2 _13020_ (.A(net1687),
    .B(_05060_),
    .C(_05076_),
    .Y(_05077_));
 sg13g2_o21ai_1 _13021_ (.B1(_05073_),
    .Y(_05078_),
    .A1(net1687),
    .A2(_05060_));
 sg13g2_nand2b_1 _13022_ (.Y(_05079_),
    .B(_05078_),
    .A_N(_05077_));
 sg13g2_nand2_1 _13023_ (.Y(_05080_),
    .A(net1697),
    .B(_05061_));
 sg13g2_a21oi_1 _13024_ (.A1(net1693),
    .A2(_05079_),
    .Y(_05081_),
    .B1(net1684));
 sg13g2_a22oi_1 _13025_ (.Y(_05082_),
    .B1(_05080_),
    .B2(_05081_),
    .A2(net2199),
    .A1(net3895));
 sg13g2_inv_1 _13026_ (.Y(_00190_),
    .A(_05082_));
 sg13g2_and2_1 _13027_ (.A(net4060),
    .B(net2199),
    .X(_05083_));
 sg13g2_o21ai_1 _13028_ (.B1(_04277_),
    .Y(_05084_),
    .A1(_04256_),
    .A2(_04278_));
 sg13g2_xor2_1 _13029_ (.B(_05084_),
    .A(_04283_),
    .X(_05085_));
 sg13g2_or2_1 _13030_ (.X(_05086_),
    .B(_05066_),
    .A(_04677_));
 sg13g2_o21ai_1 _13031_ (.B1(_05086_),
    .Y(_05087_),
    .A1(net1703),
    .A2(_04802_));
 sg13g2_nand2_1 _13032_ (.Y(_05088_),
    .A(_04576_),
    .B(net1712));
 sg13g2_o21ai_1 _13033_ (.B1(_05088_),
    .Y(_05089_),
    .A1(_04558_),
    .A2(net1712));
 sg13g2_mux2_1 _13034_ (.A0(_05023_),
    .A1(_05089_),
    .S(net1719),
    .X(_05090_));
 sg13g2_o21ai_1 _13035_ (.B1(_05090_),
    .Y(_05091_),
    .A1(net1726),
    .A2(_04954_));
 sg13g2_a221oi_1 _13036_ (.B2(_04658_),
    .C1(_05087_),
    .B1(_05091_),
    .A1(net1945),
    .Y(_05092_),
    .A2(_05085_));
 sg13g2_and2_1 _13037_ (.A(_04854_),
    .B(_05092_),
    .X(_05093_));
 sg13g2_inv_1 _13038_ (.Y(_05094_),
    .A(_05093_));
 sg13g2_mux2_1 _13039_ (.A0(_05092_),
    .A1(_05094_),
    .S(_05077_),
    .X(_05095_));
 sg13g2_nand2_1 _13040_ (.Y(_05096_),
    .A(net1692),
    .B(_05095_));
 sg13g2_a21oi_1 _13041_ (.A1(net1698),
    .A2(_05079_),
    .Y(_05097_),
    .B1(net1684));
 sg13g2_a21o_1 _13042_ (.A2(_05097_),
    .A1(_05096_),
    .B1(_05083_),
    .X(_00191_));
 sg13g2_o21ai_1 _13043_ (.B1(_04289_),
    .Y(_05098_),
    .A1(_04256_),
    .A2(_04284_));
 sg13g2_nand2_1 _13044_ (.Y(_05099_),
    .A(_04262_),
    .B(_05098_));
 sg13g2_xor2_1 _13045_ (.B(_05098_),
    .A(_04262_),
    .X(_05100_));
 sg13g2_nand3_1 _13046_ (.B(net1705),
    .C(_04820_),
    .A(net1726),
    .Y(_05101_));
 sg13g2_mux2_1 _13047_ (.A0(_04766_),
    .A1(_04770_),
    .S(net1718),
    .X(_05102_));
 sg13g2_a21oi_1 _13048_ (.A1(net1722),
    .A2(_04971_),
    .Y(_05103_),
    .B1(_05102_));
 sg13g2_o21ai_1 _13049_ (.B1(_05101_),
    .Y(_05104_),
    .A1(_04659_),
    .A2(_05103_));
 sg13g2_a22oi_1 _13050_ (.Y(_05105_),
    .B1(_05100_),
    .B2(net1945),
    .A2(_05085_),
    .A1(net1763));
 sg13g2_nand2b_1 _13051_ (.Y(_05106_),
    .B(_05105_),
    .A_N(_05104_));
 sg13g2_a21oi_1 _13052_ (.A1(_05077_),
    .A2(_05094_),
    .Y(_05107_),
    .B1(_05106_));
 sg13g2_o21ai_1 _13053_ (.B1(_04853_),
    .Y(_05108_),
    .A1(_04713_),
    .A2(_04856_));
 sg13g2_nor4_2 _13054_ (.A(_04667_),
    .B(_04713_),
    .C(_04725_),
    .Y(_05109_),
    .D(_04747_));
 sg13g2_nor3_1 _13055_ (.A(_05106_),
    .B(_05108_),
    .C(_05109_),
    .Y(_05110_));
 sg13g2_nor2_1 _13056_ (.A(_05093_),
    .B(_05110_),
    .Y(_05111_));
 sg13g2_a21o_1 _13057_ (.A2(_05111_),
    .A1(_05077_),
    .B1(_05107_),
    .X(_05112_));
 sg13g2_and2_1 _13058_ (.A(net1692),
    .B(_05112_),
    .X(_05113_));
 sg13g2_and2_1 _13059_ (.A(net1697),
    .B(_05095_),
    .X(_05114_));
 sg13g2_nor3_1 _13060_ (.A(net1684),
    .B(_05113_),
    .C(_05114_),
    .Y(_05115_));
 sg13g2_a21o_1 _13061_ (.A2(net2199),
    .A1(net3821),
    .B1(_05115_),
    .X(_00192_));
 sg13g2_nand2_1 _13062_ (.Y(_05116_),
    .A(_04261_),
    .B(_05099_));
 sg13g2_xnor2_1 _13063_ (.Y(_05117_),
    .A(_04269_),
    .B(_05116_));
 sg13g2_nor3_1 _13064_ (.A(net1723),
    .B(net1703),
    .C(_04844_),
    .Y(_05118_));
 sg13g2_nor2_1 _13065_ (.A(net1720),
    .B(_04647_),
    .Y(_05119_));
 sg13g2_nor2_1 _13066_ (.A(net1722),
    .B(_05119_),
    .Y(_05120_));
 sg13g2_o21ai_1 _13067_ (.B1(_05120_),
    .Y(_05121_),
    .A1(net1718),
    .A2(_04644_));
 sg13g2_a21oi_1 _13068_ (.A1(net1723),
    .A2(_04987_),
    .Y(_05122_),
    .B1(_04659_));
 sg13g2_a221oi_1 _13069_ (.B2(_05122_),
    .C1(_05118_),
    .B1(_05121_),
    .A1(net1762),
    .Y(_05123_),
    .A2(_05100_));
 sg13g2_o21ai_1 _13070_ (.B1(_05123_),
    .Y(_05124_),
    .A1(net1950),
    .A2(_05117_));
 sg13g2_a21oi_1 _13071_ (.A1(_05077_),
    .A2(_05111_),
    .Y(_05125_),
    .B1(_05124_));
 sg13g2_nor2_1 _13072_ (.A(_05108_),
    .B(_05124_),
    .Y(_05126_));
 sg13g2_nand2b_1 _13073_ (.Y(_05127_),
    .B(_05111_),
    .A_N(_05126_));
 sg13g2_nor4_1 _13074_ (.A(net1687),
    .B(_05060_),
    .C(_05076_),
    .D(_05127_),
    .Y(_05128_));
 sg13g2_nor2_1 _13075_ (.A(_05125_),
    .B(_05128_),
    .Y(_05129_));
 sg13g2_nor2_1 _13076_ (.A(net1697),
    .B(_05129_),
    .Y(_05130_));
 sg13g2_and2_1 _13077_ (.A(net1697),
    .B(_05112_),
    .X(_05131_));
 sg13g2_nor3_1 _13078_ (.A(net1684),
    .B(_05130_),
    .C(_05131_),
    .Y(_05132_));
 sg13g2_a21o_1 _13079_ (.A2(net2200),
    .A1(net3812),
    .B1(_05132_),
    .X(_00193_));
 sg13g2_nand2_1 _13080_ (.Y(_05133_),
    .A(net1763),
    .B(_05117_));
 sg13g2_nand3_1 _13081_ (.B(_04291_),
    .C(_04297_),
    .A(_04286_),
    .Y(_05134_));
 sg13g2_nand2_1 _13082_ (.Y(_05135_),
    .A(_04298_),
    .B(_05134_));
 sg13g2_nand2_1 _13083_ (.Y(_05136_),
    .A(net1945),
    .B(_05135_));
 sg13g2_or2_1 _13084_ (.X(_05137_),
    .B(_05003_),
    .A(net1726));
 sg13g2_nand2_1 _13085_ (.Y(_05138_),
    .A(_04622_),
    .B(_05068_));
 sg13g2_nand2_1 _13086_ (.Y(_05139_),
    .A(_04553_),
    .B(net1712));
 sg13g2_o21ai_1 _13087_ (.B1(_05139_),
    .Y(_05140_),
    .A1(_04546_),
    .A2(net1713));
 sg13g2_nand4_1 _13088_ (.B(_05137_),
    .C(_05138_),
    .A(_04658_),
    .Y(_05141_),
    .D(_05140_));
 sg13g2_nand2_1 _13089_ (.Y(_05142_),
    .A(net1705),
    .B(_04868_));
 sg13g2_nand4_1 _13090_ (.B(_05136_),
    .C(_05141_),
    .A(_05133_),
    .Y(_05143_),
    .D(_05142_));
 sg13g2_nor2b_1 _13091_ (.A(_05128_),
    .B_N(_05143_),
    .Y(_05144_));
 sg13g2_a21o_1 _13092_ (.A2(_04874_),
    .A1(_04853_),
    .B1(_04854_),
    .X(_05145_));
 sg13g2_and2_1 _13093_ (.A(_05143_),
    .B(_05145_),
    .X(_05146_));
 sg13g2_nor2b_1 _13094_ (.A(_05146_),
    .B_N(_05128_),
    .Y(_05147_));
 sg13g2_or2_1 _13095_ (.X(_05148_),
    .B(_05147_),
    .A(_05144_));
 sg13g2_nor2_1 _13096_ (.A(net1692),
    .B(_05129_),
    .Y(_05149_));
 sg13g2_a21oi_1 _13097_ (.A1(net1692),
    .A2(_05148_),
    .Y(_05150_),
    .B1(net1684));
 sg13g2_nor2b_1 _13098_ (.A(_05149_),
    .B_N(_05150_),
    .Y(_05151_));
 sg13g2_a21o_1 _13099_ (.A2(net2200),
    .A1(net3807),
    .B1(_05151_),
    .X(_00194_));
 sg13g2_and2_1 _13100_ (.A(net4053),
    .B(net2200),
    .X(_05152_));
 sg13g2_xnor2_1 _13101_ (.Y(_05153_),
    .A(_03600_),
    .B(_03663_));
 sg13g2_nand2_1 _13102_ (.Y(_05154_),
    .A(_04296_),
    .B(_04298_));
 sg13g2_xor2_1 _13103_ (.B(_05154_),
    .A(_05153_),
    .X(_05155_));
 sg13g2_nand2_1 _13104_ (.Y(_05156_),
    .A(net1945),
    .B(_05155_));
 sg13g2_nand2_1 _13105_ (.Y(_05157_),
    .A(_04551_),
    .B(net1713));
 sg13g2_nand2b_1 _13106_ (.Y(_05158_),
    .B(_04547_),
    .A_N(net1713));
 sg13g2_o21ai_1 _13107_ (.B1(_04658_),
    .Y(_05159_),
    .A1(net1718),
    .A2(_05089_));
 sg13g2_a221oi_1 _13108_ (.B2(_05158_),
    .C1(_05159_),
    .B1(_05157_),
    .A1(net1722),
    .Y(_05160_),
    .A2(_05025_));
 sg13g2_a221oi_1 _13109_ (.B2(net1763),
    .C1(_05160_),
    .B1(_05135_),
    .A1(_04669_),
    .Y(_05161_),
    .A2(_04888_));
 sg13g2_nand2_1 _13110_ (.Y(_05162_),
    .A(_05156_),
    .B(_05161_));
 sg13g2_nand3_1 _13111_ (.B(net1699),
    .C(_04855_),
    .A(_04712_),
    .Y(_05163_));
 sg13g2_nand3_1 _13112_ (.B(_05162_),
    .C(_05163_),
    .A(_04853_),
    .Y(_05164_));
 sg13g2_mux2_1 _13113_ (.A0(_05162_),
    .A1(_05164_),
    .S(_05147_),
    .X(_05165_));
 sg13g2_nand2_1 _13114_ (.Y(_05166_),
    .A(net1692),
    .B(_05165_));
 sg13g2_a21oi_1 _13115_ (.A1(net1698),
    .A2(_05148_),
    .Y(_05167_),
    .B1(net1684));
 sg13g2_a21o_1 _13116_ (.A2(_05167_),
    .A1(_05166_),
    .B1(_05152_),
    .X(_00195_));
 sg13g2_nand2_2 _13117_ (.Y(_05168_),
    .A(\data_to_write[0] ),
    .B(net2279));
 sg13g2_and3_1 _13118_ (.X(_05169_),
    .A(\addr[8] ),
    .B(\addr[7] ),
    .C(\addr[6] ));
 sg13g2_o21ai_1 _13119_ (.B1(\addr[10] ),
    .Y(_05170_),
    .A1(\addr[9] ),
    .A2(_05169_));
 sg13g2_nor4_2 _13120_ (.A(_00947_),
    .B(\i_tinyqv.cpu.data_write_n[0] ),
    .C(net2302),
    .Y(_05171_),
    .D(net2195));
 sg13g2_nand2_1 _13121_ (.Y(_05172_),
    .A(net2386),
    .B(net2388));
 sg13g2_and2_1 _13122_ (.A(\addr[5] ),
    .B(_01921_),
    .X(_05173_));
 sg13g2_inv_1 _13123_ (.Y(_05174_),
    .A(_05173_));
 sg13g2_nand2_2 _13124_ (.Y(_05175_),
    .A(net2385),
    .B(_05173_));
 sg13g2_nor2_2 _13125_ (.A(_05172_),
    .B(_05175_),
    .Y(_05176_));
 sg13g2_or2_1 _13126_ (.X(_05177_),
    .B(_05175_),
    .A(_05172_));
 sg13g2_and2_1 _13127_ (.A(_05171_),
    .B(net2090),
    .X(_05178_));
 sg13g2_nand2_1 _13128_ (.Y(_05179_),
    .A(_05171_),
    .B(net2090));
 sg13g2_nand2_2 _13129_ (.Y(_05180_),
    .A(net2275),
    .B(net2038));
 sg13g2_a22oi_1 _13130_ (.Y(_00196_),
    .B1(_05180_),
    .B2(_05168_),
    .A2(net2038),
    .A1(_01063_));
 sg13g2_o21ai_1 _13131_ (.B1(net2281),
    .Y(_05181_),
    .A1(net3502),
    .A2(net2047));
 sg13g2_a21oi_1 _13132_ (.A1(_00973_),
    .A2(net2047),
    .Y(_00197_),
    .B1(_05181_));
 sg13g2_o21ai_1 _13133_ (.B1(net2276),
    .Y(_05182_),
    .A1(net3586),
    .A2(net2046));
 sg13g2_a21oi_1 _13134_ (.A1(_00972_),
    .A2(net2046),
    .Y(_00198_),
    .B1(_05182_));
 sg13g2_o21ai_1 _13135_ (.B1(net2276),
    .Y(_05183_),
    .A1(net3446),
    .A2(net2046));
 sg13g2_a21oi_1 _13136_ (.A1(_00971_),
    .A2(net2046),
    .Y(_00199_),
    .B1(_05183_));
 sg13g2_o21ai_1 _13137_ (.B1(net2277),
    .Y(_05184_),
    .A1(net3393),
    .A2(net2046));
 sg13g2_a21oi_1 _13138_ (.A1(_00970_),
    .A2(net2046),
    .Y(_00200_),
    .B1(_05184_));
 sg13g2_o21ai_1 _13139_ (.B1(net2276),
    .Y(_05185_),
    .A1(net3487),
    .A2(net2048));
 sg13g2_a21oi_1 _13140_ (.A1(net2352),
    .A2(net2048),
    .Y(_00201_),
    .B1(_05185_));
 sg13g2_o21ai_1 _13141_ (.B1(net2281),
    .Y(_05186_),
    .A1(net3549),
    .A2(net2047));
 sg13g2_a21oi_1 _13142_ (.A1(_00968_),
    .A2(net2047),
    .Y(_00202_),
    .B1(_05186_));
 sg13g2_o21ai_1 _13143_ (.B1(net2281),
    .Y(_05187_),
    .A1(net3511),
    .A2(net2046));
 sg13g2_a21oi_1 _13144_ (.A1(_00967_),
    .A2(net2046),
    .Y(_00203_),
    .B1(_05187_));
 sg13g2_o21ai_1 _13145_ (.B1(net2279),
    .Y(_05188_),
    .A1(\data_to_write[8] ),
    .A2(net2038));
 sg13g2_a21oi_1 _13146_ (.A1(_01062_),
    .A2(net2038),
    .Y(_00204_),
    .B1(_05188_));
 sg13g2_o21ai_1 _13147_ (.B1(net2277),
    .Y(_05189_),
    .A1(net3463),
    .A2(net2041));
 sg13g2_a21oi_1 _13148_ (.A1(_00966_),
    .A2(net2041),
    .Y(_00205_),
    .B1(_05189_));
 sg13g2_o21ai_1 _13149_ (.B1(net2275),
    .Y(_05190_),
    .A1(\data_to_write[10] ),
    .A2(net2038));
 sg13g2_a21oi_1 _13150_ (.A1(_01060_),
    .A2(net2038),
    .Y(_00206_),
    .B1(_05190_));
 sg13g2_o21ai_1 _13151_ (.B1(net2276),
    .Y(_05191_),
    .A1(\data_to_write[11] ),
    .A2(net2039));
 sg13g2_a21oi_1 _13152_ (.A1(_01059_),
    .A2(net2039),
    .Y(_00207_),
    .B1(_05191_));
 sg13g2_o21ai_1 _13153_ (.B1(net2275),
    .Y(_05192_),
    .A1(\data_to_write[12] ),
    .A2(net2039));
 sg13g2_a21oi_1 _13154_ (.A1(_01058_),
    .A2(net2038),
    .Y(_00208_),
    .B1(_05192_));
 sg13g2_o21ai_1 _13155_ (.B1(net2280),
    .Y(_05193_),
    .A1(net3632),
    .A2(net2044));
 sg13g2_a21oi_1 _13156_ (.A1(_00965_),
    .A2(net2044),
    .Y(_00209_),
    .B1(_05193_));
 sg13g2_o21ai_1 _13157_ (.B1(net2278),
    .Y(_05194_),
    .A1(net3370),
    .A2(net2040));
 sg13g2_a21oi_1 _13158_ (.A1(_00964_),
    .A2(net2040),
    .Y(_00210_),
    .B1(_05194_));
 sg13g2_o21ai_1 _13159_ (.B1(net2280),
    .Y(_05195_),
    .A1(\i_peripherals.i_user_peri39.instr[15] ),
    .A2(net2042));
 sg13g2_a21oi_1 _13160_ (.A1(_00963_),
    .A2(net2042),
    .Y(_00211_),
    .B1(_05195_));
 sg13g2_o21ai_1 _13161_ (.B1(net2280),
    .Y(_05196_),
    .A1(\i_peripherals.i_user_peri39.instr[16] ),
    .A2(net2044));
 sg13g2_a21oi_1 _13162_ (.A1(_00962_),
    .A2(net2044),
    .Y(_00212_),
    .B1(_05196_));
 sg13g2_o21ai_1 _13163_ (.B1(net2280),
    .Y(_05197_),
    .A1(\i_peripherals.i_user_peri39.instr[17] ),
    .A2(net2042));
 sg13g2_a21oi_1 _13164_ (.A1(_00961_),
    .A2(net2042),
    .Y(_00213_),
    .B1(_05197_));
 sg13g2_o21ai_1 _13165_ (.B1(net2280),
    .Y(_05198_),
    .A1(\i_peripherals.i_user_peri39.instr[18] ),
    .A2(net2044));
 sg13g2_a21oi_1 _13166_ (.A1(_00960_),
    .A2(net2044),
    .Y(_00214_),
    .B1(_05198_));
 sg13g2_o21ai_1 _13167_ (.B1(net2280),
    .Y(_05199_),
    .A1(\i_peripherals.i_user_peri39.instr[19] ),
    .A2(net2042));
 sg13g2_a21oi_1 _13168_ (.A1(_00959_),
    .A2(net2042),
    .Y(_00215_),
    .B1(_05199_));
 sg13g2_o21ai_1 _13169_ (.B1(net2276),
    .Y(_05200_),
    .A1(\data_to_write[20] ),
    .A2(net2039));
 sg13g2_a21oi_1 _13170_ (.A1(_01056_),
    .A2(net2039),
    .Y(_00216_),
    .B1(_05200_));
 sg13g2_o21ai_1 _13171_ (.B1(net2278),
    .Y(_05201_),
    .A1(net3698),
    .A2(net2048));
 sg13g2_a21oi_1 _13172_ (.A1(_00958_),
    .A2(net2048),
    .Y(_00217_),
    .B1(_05201_));
 sg13g2_o21ai_1 _13173_ (.B1(net2276),
    .Y(_05202_),
    .A1(\i_peripherals.i_user_peri39.instr[22] ),
    .A2(net2048));
 sg13g2_a21oi_1 _13174_ (.A1(_00957_),
    .A2(net2041),
    .Y(_00218_),
    .B1(_05202_));
 sg13g2_o21ai_1 _13175_ (.B1(net2276),
    .Y(_05203_),
    .A1(\i_peripherals.i_user_peri39.instr[23] ),
    .A2(net2048));
 sg13g2_a21oi_1 _13176_ (.A1(_00956_),
    .A2(net2048),
    .Y(_00219_),
    .B1(_05203_));
 sg13g2_o21ai_1 _13177_ (.B1(net2276),
    .Y(_05204_),
    .A1(net3451),
    .A2(net2040));
 sg13g2_a21oi_1 _13178_ (.A1(_00955_),
    .A2(net2040),
    .Y(_00220_),
    .B1(_05204_));
 sg13g2_o21ai_1 _13179_ (.B1(net2280),
    .Y(_05205_),
    .A1(net3341),
    .A2(net2043));
 sg13g2_a21oi_1 _13180_ (.A1(_00954_),
    .A2(net2043),
    .Y(_00221_),
    .B1(_05205_));
 sg13g2_o21ai_1 _13181_ (.B1(net2278),
    .Y(_05206_),
    .A1(\i_peripherals.i_user_peri39.instr[26] ),
    .A2(net2043));
 sg13g2_a21oi_1 _13182_ (.A1(_00953_),
    .A2(net2043),
    .Y(_00222_),
    .B1(_05206_));
 sg13g2_o21ai_1 _13183_ (.B1(net2278),
    .Y(_05207_),
    .A1(net3467),
    .A2(net2040));
 sg13g2_a21oi_1 _13184_ (.A1(_00952_),
    .A2(net2040),
    .Y(_00223_),
    .B1(_05207_));
 sg13g2_o21ai_1 _13185_ (.B1(net2280),
    .Y(_05208_),
    .A1(net3375),
    .A2(net2042));
 sg13g2_a21oi_1 _13186_ (.A1(_00951_),
    .A2(net2042),
    .Y(_00224_),
    .B1(_05208_));
 sg13g2_o21ai_1 _13187_ (.B1(net2278),
    .Y(_05209_),
    .A1(net3372),
    .A2(net2040));
 sg13g2_a21oi_1 _13188_ (.A1(_00950_),
    .A2(net2040),
    .Y(_00225_),
    .B1(_05209_));
 sg13g2_o21ai_1 _13189_ (.B1(net2283),
    .Y(_05210_),
    .A1(net3492),
    .A2(net2044));
 sg13g2_a21oi_1 _13190_ (.A1(_00949_),
    .A2(net2045),
    .Y(_00226_),
    .B1(_05210_));
 sg13g2_o21ai_1 _13191_ (.B1(net2283),
    .Y(_05211_),
    .A1(net3381),
    .A2(net2045));
 sg13g2_a21oi_1 _13192_ (.A1(_00948_),
    .A2(net2044),
    .Y(_00227_),
    .B1(_05211_));
 sg13g2_nand2_1 _13193_ (.Y(_05212_),
    .A(net3763),
    .B(_02362_));
 sg13g2_o21ai_1 _13194_ (.B1(net3982),
    .Y(_05213_),
    .A1(net3532),
    .A2(net2884));
 sg13g2_nand2_1 _13195_ (.Y(_05214_),
    .A(_02362_),
    .B(_05213_));
 sg13g2_nand4_1 _13196_ (.B(_02364_),
    .C(_05212_),
    .A(net2267),
    .Y(_00228_),
    .D(_05213_));
 sg13g2_nand2_2 _13197_ (.Y(_05215_),
    .A(_01921_),
    .B(_01950_));
 sg13g2_nor2_2 _13198_ (.A(net2386),
    .B(net2388),
    .Y(_05216_));
 sg13g2_nor2b_2 _13199_ (.A(_05215_),
    .B_N(_05216_),
    .Y(_05217_));
 sg13g2_nand3_1 _13200_ (.B(net2087),
    .C(net2179),
    .A(_05171_),
    .Y(_05218_));
 sg13g2_nand2_1 _13201_ (.Y(_05219_),
    .A(net2945),
    .B(net2035));
 sg13g2_o21ai_1 _13202_ (.B1(_05219_),
    .Y(_00229_),
    .A1(net2351),
    .A2(net2037));
 sg13g2_nand2_1 _13203_ (.Y(_05220_),
    .A(net3072),
    .B(net2035));
 sg13g2_o21ai_1 _13204_ (.B1(_05220_),
    .Y(_00230_),
    .A1(_00973_),
    .A2(net2036));
 sg13g2_nand2_1 _13205_ (.Y(_05221_),
    .A(net2962),
    .B(net2035));
 sg13g2_o21ai_1 _13206_ (.B1(_05221_),
    .Y(_00231_),
    .A1(_00972_),
    .A2(net2036));
 sg13g2_nand2_1 _13207_ (.Y(_05222_),
    .A(net3124),
    .B(net2035));
 sg13g2_o21ai_1 _13208_ (.B1(_05222_),
    .Y(_00232_),
    .A1(_00971_),
    .A2(net2036));
 sg13g2_nand2_1 _13209_ (.Y(_05223_),
    .A(net3030),
    .B(net2036));
 sg13g2_o21ai_1 _13210_ (.B1(_05223_),
    .Y(_00233_),
    .A1(_00970_),
    .A2(net2032));
 sg13g2_nand2_1 _13211_ (.Y(_05224_),
    .A(net2928),
    .B(net2035));
 sg13g2_o21ai_1 _13212_ (.B1(_05224_),
    .Y(_00234_),
    .A1(net2352),
    .A2(net2035));
 sg13g2_nand2_1 _13213_ (.Y(_05225_),
    .A(net2995),
    .B(net2036));
 sg13g2_o21ai_1 _13214_ (.B1(_05225_),
    .Y(_00235_),
    .A1(_00968_),
    .A2(net2036));
 sg13g2_nand2_1 _13215_ (.Y(_05226_),
    .A(net2922),
    .B(net2031));
 sg13g2_o21ai_1 _13216_ (.B1(_05226_),
    .Y(_00236_),
    .A1(_00967_),
    .A2(net2031));
 sg13g2_mux2_1 _13217_ (.A0(\data_to_write[8] ),
    .A1(net3584),
    .S(net2035),
    .X(_00237_));
 sg13g2_nand2_1 _13218_ (.Y(_05227_),
    .A(net2993),
    .B(net2031));
 sg13g2_o21ai_1 _13219_ (.B1(_05227_),
    .Y(_00238_),
    .A1(_00966_),
    .A2(net2031));
 sg13g2_mux2_1 _13220_ (.A0(\data_to_write[10] ),
    .A1(net3563),
    .S(net2037),
    .X(_00239_));
 sg13g2_mux2_1 _13221_ (.A0(\data_to_write[11] ),
    .A1(net3559),
    .S(net2035),
    .X(_00240_));
 sg13g2_mux2_1 _13222_ (.A0(\data_to_write[12] ),
    .A1(net3634),
    .S(net2036),
    .X(_00241_));
 sg13g2_nand2_1 _13223_ (.Y(_05228_),
    .A(net2977),
    .B(net2033));
 sg13g2_o21ai_1 _13224_ (.B1(_05228_),
    .Y(_00242_),
    .A1(_00965_),
    .A2(net2033));
 sg13g2_nand2_1 _13225_ (.Y(_05229_),
    .A(net3026),
    .B(net2034));
 sg13g2_o21ai_1 _13226_ (.B1(_05229_),
    .Y(_00243_),
    .A1(_00964_),
    .A2(net2034));
 sg13g2_nand2_1 _13227_ (.Y(_05230_),
    .A(net3108),
    .B(net2030));
 sg13g2_o21ai_1 _13228_ (.B1(_05230_),
    .Y(_00244_),
    .A1(_00963_),
    .A2(net2032));
 sg13g2_nand2_1 _13229_ (.Y(_05231_),
    .A(net2926),
    .B(net2033));
 sg13g2_o21ai_1 _13230_ (.B1(_05231_),
    .Y(_00245_),
    .A1(_00962_),
    .A2(net2033));
 sg13g2_nand2_1 _13231_ (.Y(_05232_),
    .A(net3085),
    .B(net2029));
 sg13g2_o21ai_1 _13232_ (.B1(_05232_),
    .Y(_00246_),
    .A1(_00961_),
    .A2(net2029));
 sg13g2_nand2_1 _13233_ (.Y(_05233_),
    .A(net2872),
    .B(net2033));
 sg13g2_o21ai_1 _13234_ (.B1(_05233_),
    .Y(_00247_),
    .A1(_00960_),
    .A2(net2033));
 sg13g2_nand2_1 _13235_ (.Y(_05234_),
    .A(net3001),
    .B(net2030));
 sg13g2_o21ai_1 _13236_ (.B1(_05234_),
    .Y(_00248_),
    .A1(_00959_),
    .A2(net2030));
 sg13g2_mux2_1 _13237_ (.A0(\data_to_write[20] ),
    .A1(net3683),
    .S(net2030),
    .X(_00249_));
 sg13g2_nand2_1 _13238_ (.Y(_05235_),
    .A(net2951),
    .B(net2029));
 sg13g2_o21ai_1 _13239_ (.B1(_05235_),
    .Y(_00250_),
    .A1(_00958_),
    .A2(net2029));
 sg13g2_nand2_1 _13240_ (.Y(_05236_),
    .A(net3150),
    .B(net2029));
 sg13g2_o21ai_1 _13241_ (.B1(_05236_),
    .Y(_00251_),
    .A1(_00957_),
    .A2(net2029));
 sg13g2_nand2_1 _13242_ (.Y(_05237_),
    .A(net3011),
    .B(net2031));
 sg13g2_o21ai_1 _13243_ (.B1(_05237_),
    .Y(_00252_),
    .A1(_00956_),
    .A2(net2031));
 sg13g2_nand2_1 _13244_ (.Y(_05238_),
    .A(net2939),
    .B(net2031));
 sg13g2_o21ai_1 _13245_ (.B1(_05238_),
    .Y(_00253_),
    .A1(_00955_),
    .A2(net2031));
 sg13g2_nand2_1 _13246_ (.Y(_05239_),
    .A(net3206),
    .B(net2032));
 sg13g2_o21ai_1 _13247_ (.B1(_05239_),
    .Y(_00254_),
    .A1(_00954_),
    .A2(net2032));
 sg13g2_nand2_1 _13248_ (.Y(_05240_),
    .A(net2886),
    .B(net2029));
 sg13g2_o21ai_1 _13249_ (.B1(_05240_),
    .Y(_00255_),
    .A1(_00953_),
    .A2(net2029));
 sg13g2_nand2_1 _13250_ (.Y(_05241_),
    .A(net2924),
    .B(net2033));
 sg13g2_o21ai_1 _13251_ (.B1(_05241_),
    .Y(_00256_),
    .A1(_00952_),
    .A2(net2034));
 sg13g2_nand2_1 _13252_ (.Y(_05242_),
    .A(net2979),
    .B(net2030));
 sg13g2_o21ai_1 _13253_ (.B1(_05242_),
    .Y(_00257_),
    .A1(_00951_),
    .A2(net2030));
 sg13g2_nand2_1 _13254_ (.Y(_05243_),
    .A(net2933),
    .B(net2034));
 sg13g2_o21ai_1 _13255_ (.B1(_05243_),
    .Y(_00258_),
    .A1(_00950_),
    .A2(net2034));
 sg13g2_nand2_1 _13256_ (.Y(_05244_),
    .A(net2918),
    .B(net2034));
 sg13g2_o21ai_1 _13257_ (.B1(_05244_),
    .Y(_00259_),
    .A1(_00949_),
    .A2(net2034));
 sg13g2_nand2_1 _13258_ (.Y(_05245_),
    .A(net3051),
    .B(net2033));
 sg13g2_o21ai_1 _13259_ (.B1(_05245_),
    .Y(_00260_),
    .A1(_00948_),
    .A2(net2030));
 sg13g2_nor2b_2 _13260_ (.A(net2386),
    .B_N(net2388),
    .Y(_05246_));
 sg13g2_nor2b_2 _13261_ (.A(_05215_),
    .B_N(_05246_),
    .Y(_05247_));
 sg13g2_nand3_1 _13262_ (.B(net2087),
    .C(net2172),
    .A(_05171_),
    .Y(_05248_));
 sg13g2_nand2_1 _13263_ (.Y(_05249_),
    .A(net3035),
    .B(net2026));
 sg13g2_o21ai_1 _13264_ (.B1(_05249_),
    .Y(_00261_),
    .A1(net2351),
    .A2(net2027));
 sg13g2_nand2_1 _13265_ (.Y(_05250_),
    .A(net3033),
    .B(net2026));
 sg13g2_o21ai_1 _13266_ (.B1(_05250_),
    .Y(_00262_),
    .A1(_00973_),
    .A2(net2028));
 sg13g2_nand2_1 _13267_ (.Y(_05251_),
    .A(net3047),
    .B(net2026));
 sg13g2_o21ai_1 _13268_ (.B1(_05251_),
    .Y(_00263_),
    .A1(_00972_),
    .A2(net2027));
 sg13g2_nand2_1 _13269_ (.Y(_05252_),
    .A(net3036),
    .B(net2026));
 sg13g2_o21ai_1 _13270_ (.B1(_05252_),
    .Y(_00264_),
    .A1(_00971_),
    .A2(net2027));
 sg13g2_nand2_1 _13271_ (.Y(_05253_),
    .A(net3040),
    .B(net2023));
 sg13g2_o21ai_1 _13272_ (.B1(_05253_),
    .Y(_00265_),
    .A1(_00970_),
    .A2(net2023));
 sg13g2_nand2_1 _13273_ (.Y(_05254_),
    .A(net2969),
    .B(net2026));
 sg13g2_o21ai_1 _13274_ (.B1(_05254_),
    .Y(_00266_),
    .A1(net2352),
    .A2(net2026));
 sg13g2_nand2_1 _13275_ (.Y(_05255_),
    .A(net3152),
    .B(net2027));
 sg13g2_o21ai_1 _13276_ (.B1(_05255_),
    .Y(_00267_),
    .A1(_00968_),
    .A2(net2027));
 sg13g2_nand2_1 _13277_ (.Y(_05256_),
    .A(net2904),
    .B(net2022));
 sg13g2_o21ai_1 _13278_ (.B1(_05256_),
    .Y(_00268_),
    .A1(_00967_),
    .A2(net2022));
 sg13g2_mux2_1 _13279_ (.A0(\data_to_write[8] ),
    .A1(net3609),
    .S(net2026),
    .X(_00269_));
 sg13g2_nand2_1 _13280_ (.Y(_05257_),
    .A(net2970),
    .B(net2022));
 sg13g2_o21ai_1 _13281_ (.B1(_05257_),
    .Y(_00270_),
    .A1(_00966_),
    .A2(net2022));
 sg13g2_mux2_1 _13282_ (.A0(\data_to_write[10] ),
    .A1(net3556),
    .S(net2027),
    .X(_00271_));
 sg13g2_mux2_1 _13283_ (.A0(\data_to_write[11] ),
    .A1(net3588),
    .S(net2026),
    .X(_00272_));
 sg13g2_mux2_1 _13284_ (.A0(\data_to_write[12] ),
    .A1(net3668),
    .S(net2027),
    .X(_00273_));
 sg13g2_nand2_1 _13285_ (.Y(_05258_),
    .A(net3028),
    .B(net2024));
 sg13g2_o21ai_1 _13286_ (.B1(_05258_),
    .Y(_00274_),
    .A1(_00965_),
    .A2(net2024));
 sg13g2_nand2_1 _13287_ (.Y(_05259_),
    .A(net2964),
    .B(net2025));
 sg13g2_o21ai_1 _13288_ (.B1(_05259_),
    .Y(_00275_),
    .A1(_00964_),
    .A2(net2025));
 sg13g2_nand2_1 _13289_ (.Y(_05260_),
    .A(net3066),
    .B(net2021));
 sg13g2_o21ai_1 _13290_ (.B1(_05260_),
    .Y(_00276_),
    .A1(_00963_),
    .A2(net2023));
 sg13g2_nand2_1 _13291_ (.Y(_05261_),
    .A(net2822),
    .B(net2024));
 sg13g2_o21ai_1 _13292_ (.B1(_05261_),
    .Y(_00277_),
    .A1(_00962_),
    .A2(net2024));
 sg13g2_nand2_1 _13293_ (.Y(_05262_),
    .A(net2865),
    .B(net2020));
 sg13g2_o21ai_1 _13294_ (.B1(_05262_),
    .Y(_00278_),
    .A1(_00961_),
    .A2(net2020));
 sg13g2_nand2_1 _13295_ (.Y(_05263_),
    .A(net2960),
    .B(net2024));
 sg13g2_o21ai_1 _13296_ (.B1(_05263_),
    .Y(_00279_),
    .A1(_00960_),
    .A2(net2024));
 sg13g2_nand2_1 _13297_ (.Y(_05264_),
    .A(net2981),
    .B(net2021));
 sg13g2_o21ai_1 _13298_ (.B1(_05264_),
    .Y(_00280_),
    .A1(_00959_),
    .A2(net2021));
 sg13g2_mux2_1 _13299_ (.A0(\data_to_write[20] ),
    .A1(net3735),
    .S(net2021),
    .X(_00281_));
 sg13g2_nand2_1 _13300_ (.Y(_05265_),
    .A(net2911),
    .B(net2020));
 sg13g2_o21ai_1 _13301_ (.B1(_05265_),
    .Y(_00282_),
    .A1(_00958_),
    .A2(net2020));
 sg13g2_nand2_1 _13302_ (.Y(_05266_),
    .A(net2983),
    .B(net2020));
 sg13g2_o21ai_1 _13303_ (.B1(_05266_),
    .Y(_00283_),
    .A1(_00957_),
    .A2(net2020));
 sg13g2_nand2_1 _13304_ (.Y(_05267_),
    .A(net3013),
    .B(net2022));
 sg13g2_o21ai_1 _13305_ (.B1(_05267_),
    .Y(_00284_),
    .A1(_00956_),
    .A2(net2022));
 sg13g2_nand2_1 _13306_ (.Y(_05268_),
    .A(net2849),
    .B(net2022));
 sg13g2_o21ai_1 _13307_ (.B1(_05268_),
    .Y(_00285_),
    .A1(_00955_),
    .A2(net2022));
 sg13g2_nand2_1 _13308_ (.Y(_05269_),
    .A(net2817),
    .B(net2023));
 sg13g2_o21ai_1 _13309_ (.B1(_05269_),
    .Y(_00286_),
    .A1(_00954_),
    .A2(net2023));
 sg13g2_nand2_1 _13310_ (.Y(_05270_),
    .A(net2972),
    .B(net2020));
 sg13g2_o21ai_1 _13311_ (.B1(_05270_),
    .Y(_00287_),
    .A1(_00953_),
    .A2(net2021));
 sg13g2_nand2_1 _13312_ (.Y(_05271_),
    .A(net2900),
    .B(net2025));
 sg13g2_o21ai_1 _13313_ (.B1(_05271_),
    .Y(_00288_),
    .A1(_00952_),
    .A2(net2024));
 sg13g2_nand2_1 _13314_ (.Y(_05272_),
    .A(net2955),
    .B(net2021));
 sg13g2_o21ai_1 _13315_ (.B1(_05272_),
    .Y(_00289_),
    .A1(_00951_),
    .A2(net2020));
 sg13g2_nand2_1 _13316_ (.Y(_05273_),
    .A(net2987),
    .B(net2025));
 sg13g2_o21ai_1 _13317_ (.B1(_05273_),
    .Y(_00290_),
    .A1(_00950_),
    .A2(net2025));
 sg13g2_nand2_1 _13318_ (.Y(_05274_),
    .A(net2853),
    .B(net2025));
 sg13g2_o21ai_1 _13319_ (.B1(_05274_),
    .Y(_00291_),
    .A1(_00949_),
    .A2(net2025));
 sg13g2_nand2_1 _13320_ (.Y(_05275_),
    .A(net2898),
    .B(net2024));
 sg13g2_o21ai_1 _13321_ (.B1(_05275_),
    .Y(_00292_),
    .A1(_00948_),
    .A2(net2021));
 sg13g2_nor3_2 _13322_ (.A(net4171),
    .B(net4164),
    .C(net3022),
    .Y(_05276_));
 sg13g2_nor3_1 _13323_ (.A(net3022),
    .B(_05180_),
    .C(_05276_),
    .Y(_00293_));
 sg13g2_nand3_1 _13324_ (.B(_01054_),
    .C(_01055_),
    .A(\i_peripherals.i_user_peri39.busy_counter[2] ),
    .Y(_05277_));
 sg13g2_nand2_1 _13325_ (.Y(_05278_),
    .A(net3702),
    .B(net3022));
 sg13g2_a21oi_1 _13326_ (.A1(_05277_),
    .A2(_05278_),
    .Y(_00294_),
    .B1(_05180_));
 sg13g2_nor2_2 _13327_ (.A(_02577_),
    .B(_02639_),
    .Y(_05279_));
 sg13g2_nor2_1 _13328_ (.A(net2346),
    .B(_05279_),
    .Y(_05280_));
 sg13g2_nand2_2 _13329_ (.Y(_05281_),
    .A(net2494),
    .B(_05279_));
 sg13g2_nor2_1 _13330_ (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .B(net1760),
    .Y(_05282_));
 sg13g2_a21oi_1 _13331_ (.A1(_01089_),
    .A2(_05280_),
    .Y(_00295_),
    .B1(_05282_));
 sg13g2_nor2_1 _13332_ (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .B(net1760),
    .Y(_05283_));
 sg13g2_a21oi_1 _13333_ (.A1(_01093_),
    .A2(_05280_),
    .Y(_00296_),
    .B1(_05283_));
 sg13g2_nor2_1 _13334_ (.A(net1753),
    .B(net1752),
    .Y(_05284_));
 sg13g2_a21oi_2 _13335_ (.B1(_02805_),
    .Y(_05285_),
    .A2(_02803_),
    .A1(net2438));
 sg13g2_nand2_1 _13336_ (.Y(_05286_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .B(net2439));
 sg13g2_xnor2_1 _13337_ (.Y(_05287_),
    .A(\i_tinyqv.cpu.pc[1] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[1] ));
 sg13g2_nand2_1 _13338_ (.Y(_05288_),
    .A(net2406),
    .B(_05287_));
 sg13g2_o21ai_1 _13339_ (.B1(_05288_),
    .Y(_05289_),
    .A1(net2406),
    .A2(\i_tinyqv.cpu.instr_write_offset[1] ));
 sg13g2_nor3_1 _13340_ (.A(_02803_),
    .B(_02805_),
    .C(_02810_),
    .Y(_05290_));
 sg13g2_a22oi_1 _13341_ (.Y(_05291_),
    .B1(net1747),
    .B2(net3199),
    .A2(net2062),
    .A1(net3163));
 sg13g2_o21ai_1 _13342_ (.B1(_05291_),
    .Y(_00297_),
    .A1(_05285_),
    .A2(_05289_));
 sg13g2_nand2_1 _13343_ (.Y(_05292_),
    .A(\i_tinyqv.cpu.pc[2] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sg13g2_xnor2_1 _13344_ (.Y(_05293_),
    .A(\i_tinyqv.cpu.pc[2] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[2] ));
 sg13g2_xnor2_1 _13345_ (.Y(_05294_),
    .A(_05286_),
    .B(_05293_));
 sg13g2_nand2_1 _13346_ (.Y(_05295_),
    .A(net2406),
    .B(_05294_));
 sg13g2_o21ai_1 _13347_ (.B1(_05295_),
    .Y(_05296_),
    .A1(net2408),
    .A2(\i_tinyqv.cpu.instr_write_offset[2] ));
 sg13g2_a22oi_1 _13348_ (.Y(_05297_),
    .B1(net1746),
    .B2(net3291),
    .A2(net2062),
    .A1(net2388));
 sg13g2_o21ai_1 _13349_ (.B1(net3292),
    .Y(_00298_),
    .A1(_05285_),
    .A2(_05296_));
 sg13g2_xnor2_1 _13350_ (.Y(_05298_),
    .A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[3] ));
 sg13g2_o21ai_1 _13351_ (.B1(_05292_),
    .Y(_05299_),
    .A1(_05286_),
    .A2(_05293_));
 sg13g2_nor2b_1 _13352_ (.A(_05298_),
    .B_N(_05299_),
    .Y(_05300_));
 sg13g2_xnor2_1 _13353_ (.Y(_05301_),
    .A(_05298_),
    .B(_05299_));
 sg13g2_xnor2_1 _13354_ (.Y(_05302_),
    .A(\i_tinyqv.cpu.instr_data_start[3] ),
    .B(\i_tinyqv.cpu.instr_write_offset[3] ));
 sg13g2_nor2_1 _13355_ (.A(net2406),
    .B(_05302_),
    .Y(_05303_));
 sg13g2_a21oi_1 _13356_ (.A1(net2406),
    .A2(_05301_),
    .Y(_05304_),
    .B1(_05303_));
 sg13g2_a22oi_1 _13357_ (.Y(_05305_),
    .B1(net1746),
    .B2(net3212),
    .A2(net2062),
    .A1(\addr[3] ));
 sg13g2_o21ai_1 _13358_ (.B1(net3213),
    .Y(_00299_),
    .A1(_05285_),
    .A2(_05304_));
 sg13g2_nor2b_2 _13359_ (.A(net2388),
    .B_N(net2386),
    .Y(_05306_));
 sg13g2_nor2b_1 _13360_ (.A(_05215_),
    .B_N(_05306_),
    .Y(_05307_));
 sg13g2_or4_1 _13361_ (.A(\addr[10] ),
    .B(\addr[9] ),
    .C(\addr[8] ),
    .D(_01922_),
    .X(_05308_));
 sg13g2_nor2_2 _13362_ (.A(\addr[6] ),
    .B(_05308_),
    .Y(_05309_));
 sg13g2_and2_1 _13363_ (.A(net2165),
    .B(_05309_),
    .X(_05310_));
 sg13g2_nor3_1 _13364_ (.A(\addr[6] ),
    .B(_02430_),
    .C(_05308_),
    .Y(_05311_));
 sg13g2_nand2_1 _13365_ (.Y(_05312_),
    .A(net2165),
    .B(_05311_));
 sg13g2_a21oi_1 _13366_ (.A1(net3897),
    .A2(net2084),
    .Y(_05313_),
    .B1(net2246));
 sg13g2_o21ai_1 _13367_ (.B1(_05313_),
    .Y(_00300_),
    .A1(net2351),
    .A2(net2084));
 sg13g2_a21oi_1 _13368_ (.A1(net3938),
    .A2(net2082),
    .Y(_05314_),
    .B1(net2249));
 sg13g2_o21ai_1 _13369_ (.B1(_05314_),
    .Y(_00301_),
    .A1(_00973_),
    .A2(net2082));
 sg13g2_o21ai_1 _13370_ (.B1(net2279),
    .Y(_05315_),
    .A1(net2396),
    .A2(net2082));
 sg13g2_a21oi_1 _13371_ (.A1(_01052_),
    .A2(net2082),
    .Y(_00302_),
    .B1(_05315_));
 sg13g2_a21oi_1 _13372_ (.A1(net3934),
    .A2(net2083),
    .Y(_05316_),
    .B1(net2253));
 sg13g2_o21ai_1 _13373_ (.B1(_05316_),
    .Y(_00303_),
    .A1(_00971_),
    .A2(net2083));
 sg13g2_o21ai_1 _13374_ (.B1(net2279),
    .Y(_05317_),
    .A1(net2392),
    .A2(net2082));
 sg13g2_a21oi_1 _13375_ (.A1(_01050_),
    .A2(net2082),
    .Y(_00304_),
    .B1(_05317_));
 sg13g2_a21oi_1 _13376_ (.A1(net3860),
    .A2(net2083),
    .Y(_05318_),
    .B1(net2249));
 sg13g2_o21ai_1 _13377_ (.B1(_05318_),
    .Y(_00305_),
    .A1(net2352),
    .A2(net2083));
 sg13g2_a221oi_1 _13378_ (.B2(_01048_),
    .C1(net2249),
    .B1(net2082),
    .A1(_02436_),
    .Y(_00306_),
    .A2(net2085));
 sg13g2_o21ai_1 _13379_ (.B1(net2279),
    .Y(_05319_),
    .A1(\data_to_write[7] ),
    .A2(net2083));
 sg13g2_a21oi_1 _13380_ (.A1(_01047_),
    .A2(net2083),
    .Y(_00307_),
    .B1(_05319_));
 sg13g2_nor2_1 _13381_ (.A(net2196),
    .B(_05276_),
    .Y(_05320_));
 sg13g2_nor2_1 _13382_ (.A(_02613_),
    .B(_05320_),
    .Y(_05321_));
 sg13g2_nor2b_1 _13383_ (.A(_05180_),
    .B_N(_05321_),
    .Y(_00308_));
 sg13g2_and2_1 _13384_ (.A(net2174),
    .B(_05309_),
    .X(_05322_));
 sg13g2_nor3_1 _13385_ (.A(_01095_),
    .B(net4100),
    .C(_02613_),
    .Y(_05323_));
 sg13g2_nor2b_1 _13386_ (.A(net3835),
    .B_N(\i_peripherals.i_uart.i_uart_rx.fsm_state[1] ),
    .Y(_05324_));
 sg13g2_and2_1 _13387_ (.A(net3448),
    .B(_05324_),
    .X(_05325_));
 sg13g2_nand2_1 _13388_ (.Y(_05326_),
    .A(net3448),
    .B(_05324_));
 sg13g2_nand3_1 _13389_ (.B(net3976),
    .C(net2481),
    .A(net3448),
    .Y(_05327_));
 sg13g2_nand2_1 _13390_ (.Y(_05328_),
    .A(net2481),
    .B(_05325_));
 sg13g2_a221oi_1 _13391_ (.B2(_01095_),
    .C1(net2248),
    .B1(_05328_),
    .A1(net2081),
    .Y(_00309_),
    .A2(_05323_));
 sg13g2_nor2_1 _13392_ (.A(_05172_),
    .B(_05215_),
    .Y(_05329_));
 sg13g2_nand2_1 _13393_ (.Y(_05330_),
    .A(_05311_),
    .B(_05329_));
 sg13g2_o21ai_1 _13394_ (.B1(net2272),
    .Y(_05331_),
    .A1(net2399),
    .A2(_05330_));
 sg13g2_a21oi_1 _13395_ (.A1(_01046_),
    .A2(_05330_),
    .Y(_00310_),
    .B1(_05331_));
 sg13g2_nand2b_1 _13396_ (.Y(_05332_),
    .B(\i_peripherals.i_uart.baud_divider[6] ),
    .A_N(\i_peripherals.i_uart.i_uart_tx.cycle_counter[6] ));
 sg13g2_nand2_1 _13397_ (.Y(_05333_),
    .A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[5] ),
    .B(_01049_));
 sg13g2_nand2_1 _13398_ (.Y(_05334_),
    .A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[3] ),
    .B(_01051_));
 sg13g2_a22oi_1 _13399_ (.Y(_05335_),
    .B1(\i_peripherals.i_uart.baud_divider[0] ),
    .B2(_01045_),
    .A2(\i_peripherals.i_uart.baud_divider[1] ),
    .A1(_01044_));
 sg13g2_a221oi_1 _13400_ (.B2(\i_peripherals.i_uart.i_uart_tx.cycle_counter[1] ),
    .C1(_05335_),
    .B1(_01053_),
    .A1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[2] ),
    .Y(_05336_),
    .A2(_01052_));
 sg13g2_nor2_1 _13401_ (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[2] ),
    .B(_01052_),
    .Y(_05337_));
 sg13g2_o21ai_1 _13402_ (.B1(_05334_),
    .Y(_05338_),
    .A1(_05336_),
    .A2(_05337_));
 sg13g2_a22oi_1 _13403_ (.Y(_05339_),
    .B1(\i_peripherals.i_uart.baud_divider[3] ),
    .B2(_01043_),
    .A2(\i_peripherals.i_uart.baud_divider[4] ),
    .A1(_01042_));
 sg13g2_a22oi_1 _13404_ (.Y(_05340_),
    .B1(_05338_),
    .B2(_05339_),
    .A2(_01050_),
    .A1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[4] ));
 sg13g2_o21ai_1 _13405_ (.B1(_05332_),
    .Y(_05341_),
    .A1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[5] ),
    .A2(_01049_));
 sg13g2_a21oi_1 _13406_ (.A1(_05333_),
    .A2(_05340_),
    .Y(_05342_),
    .B1(_05341_));
 sg13g2_a221oi_1 _13407_ (.B2(\i_peripherals.i_uart.i_uart_tx.cycle_counter[6] ),
    .C1(_05342_),
    .B1(_01048_),
    .A1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[7] ),
    .Y(_05343_),
    .A2(_01047_));
 sg13g2_nand2b_1 _13408_ (.Y(_05344_),
    .B(\i_peripherals.i_uart.baud_divider[7] ),
    .A_N(\i_peripherals.i_uart.i_uart_tx.cycle_counter[7] ));
 sg13g2_o21ai_1 _13409_ (.B1(_05344_),
    .Y(_05345_),
    .A1(_00990_),
    .A2(\i_peripherals.i_uart.i_uart_tx.cycle_counter[8] ));
 sg13g2_nor2_1 _13410_ (.A(_05343_),
    .B(_05345_),
    .Y(_05346_));
 sg13g2_a221oi_1 _13411_ (.B2(_00990_),
    .C1(_05346_),
    .B1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[8] ),
    .A1(_00989_),
    .Y(_05347_),
    .A2(\i_peripherals.i_uart.i_uart_tx.cycle_counter[9] ));
 sg13g2_nand2b_1 _13412_ (.Y(_05348_),
    .B(\i_peripherals.i_uart.baud_divider[9] ),
    .A_N(\i_peripherals.i_uart.i_uart_tx.cycle_counter[9] ));
 sg13g2_o21ai_1 _13413_ (.B1(_05348_),
    .Y(_05349_),
    .A1(_00988_),
    .A2(\i_peripherals.i_uart.i_uart_tx.cycle_counter[10] ));
 sg13g2_a22oi_1 _13414_ (.Y(_05350_),
    .B1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[10] ),
    .B2(_00988_),
    .A2(\i_peripherals.i_uart.i_uart_tx.cycle_counter[11] ),
    .A1(_00987_));
 sg13g2_o21ai_1 _13415_ (.B1(_05350_),
    .Y(_05351_),
    .A1(_05347_),
    .A2(_05349_));
 sg13g2_a22oi_1 _13416_ (.Y(_05352_),
    .B1(_01041_),
    .B2(\i_peripherals.i_uart.baud_divider[11] ),
    .A2(_01040_),
    .A1(\i_peripherals.i_uart.baud_divider[12] ));
 sg13g2_a22oi_1 _13417_ (.Y(_05353_),
    .B1(_05351_),
    .B2(_05352_),
    .A2(\i_peripherals.i_uart.i_uart_tx.cycle_counter[12] ),
    .A1(_00986_));
 sg13g2_nor2_1 _13418_ (.A(_05214_),
    .B(_05353_),
    .Y(_05354_));
 sg13g2_and3_2 _13419_ (.X(_05355_),
    .A(_02363_),
    .B(_02429_),
    .C(net2081));
 sg13g2_or2_1 _13420_ (.X(_05356_),
    .B(net2019),
    .A(_05354_));
 sg13g2_nor2b_1 _13421_ (.A(net2019),
    .B_N(net3449),
    .Y(_05357_));
 sg13g2_a21oi_1 _13422_ (.A1(net2399),
    .A2(net2019),
    .Y(_05358_),
    .B1(_05357_));
 sg13g2_o21ai_1 _13423_ (.B1(net2262),
    .Y(_05359_),
    .A1(net3763),
    .A2(_05356_));
 sg13g2_a21oi_1 _13424_ (.A1(_05356_),
    .A2(_05358_),
    .Y(_00311_),
    .B1(_05359_));
 sg13g2_nor2b_1 _13425_ (.A(net2018),
    .B_N(net3299),
    .Y(_05360_));
 sg13g2_a21oi_1 _13426_ (.A1(net2397),
    .A2(net2018),
    .Y(_05361_),
    .B1(_05360_));
 sg13g2_o21ai_1 _13427_ (.B1(net2259),
    .Y(_05362_),
    .A1(net3449),
    .A2(net1896));
 sg13g2_a21oi_1 _13428_ (.A1(net1896),
    .A2(_05361_),
    .Y(_00312_),
    .B1(_05362_));
 sg13g2_nor2b_1 _13429_ (.A(net2017),
    .B_N(\i_peripherals.i_uart.i_uart_tx.data_to_send[3] ),
    .Y(_05363_));
 sg13g2_a21oi_1 _13430_ (.A1(net2395),
    .A2(net2017),
    .Y(_05364_),
    .B1(_05363_));
 sg13g2_o21ai_1 _13431_ (.B1(net2259),
    .Y(_05365_),
    .A1(net3299),
    .A2(net1896));
 sg13g2_a21oi_1 _13432_ (.A1(net1895),
    .A2(_05364_),
    .Y(_00313_),
    .B1(_05365_));
 sg13g2_nor2b_1 _13433_ (.A(net2017),
    .B_N(net3414),
    .Y(_05366_));
 sg13g2_a21oi_1 _13434_ (.A1(net2393),
    .A2(net2017),
    .Y(_05367_),
    .B1(_05366_));
 sg13g2_o21ai_1 _13435_ (.B1(net2259),
    .Y(_05368_),
    .A1(net3547),
    .A2(net1896));
 sg13g2_a21oi_1 _13436_ (.A1(net1895),
    .A2(_05367_),
    .Y(_00314_),
    .B1(_05368_));
 sg13g2_nor2b_1 _13437_ (.A(net2018),
    .B_N(net3389),
    .Y(_05369_));
 sg13g2_a21oi_1 _13438_ (.A1(net2391),
    .A2(net2018),
    .Y(_05370_),
    .B1(_05369_));
 sg13g2_o21ai_1 _13439_ (.B1(net2259),
    .Y(_05371_),
    .A1(net3414),
    .A2(net1896));
 sg13g2_a21oi_1 _13440_ (.A1(net1895),
    .A2(_05370_),
    .Y(_00315_),
    .B1(_05371_));
 sg13g2_nor2b_1 _13441_ (.A(net2017),
    .B_N(\i_peripherals.i_uart.i_uart_tx.data_to_send[6] ),
    .Y(_05372_));
 sg13g2_a21oi_1 _13442_ (.A1(net2389),
    .A2(net2017),
    .Y(_05373_),
    .B1(_05372_));
 sg13g2_o21ai_1 _13443_ (.B1(net2259),
    .Y(_05374_),
    .A1(net3389),
    .A2(net1895));
 sg13g2_a21oi_1 _13444_ (.A1(net1895),
    .A2(_05373_),
    .Y(_00316_),
    .B1(_05374_));
 sg13g2_nand2_1 _13445_ (.Y(_05375_),
    .A(_00968_),
    .B(net2018));
 sg13g2_o21ai_1 _13446_ (.B1(net2259),
    .Y(_05376_),
    .A1(net3400),
    .A2(net1895));
 sg13g2_o21ai_1 _13447_ (.B1(_05375_),
    .Y(_05377_),
    .A1(\i_peripherals.i_uart.i_uart_tx.data_to_send[7] ),
    .A2(net2017));
 sg13g2_a21oi_1 _13448_ (.A1(net1895),
    .A2(_05377_),
    .Y(_00317_),
    .B1(_05376_));
 sg13g2_nand2_1 _13449_ (.Y(_05378_),
    .A(\data_to_write[7] ),
    .B(net2018));
 sg13g2_o21ai_1 _13450_ (.B1(net2259),
    .Y(_05379_),
    .A1(net3458),
    .A2(net2017));
 sg13g2_a21oi_1 _13451_ (.A1(net1895),
    .A2(_05378_),
    .Y(_00318_),
    .B1(_05379_));
 sg13g2_nand2_2 _13452_ (.Y(_05380_),
    .A(net2267),
    .B(_05353_));
 sg13g2_nor2_1 _13453_ (.A(net3216),
    .B(_02364_),
    .Y(_05381_));
 sg13g2_nor2_1 _13454_ (.A(_01045_),
    .B(_02363_),
    .Y(_05382_));
 sg13g2_nor3_1 _13455_ (.A(net1900),
    .B(net3217),
    .C(_05382_),
    .Y(_00319_));
 sg13g2_nor3_2 _13456_ (.A(_01044_),
    .B(_01045_),
    .C(_02363_),
    .Y(_05383_));
 sg13g2_nor2_1 _13457_ (.A(net3337),
    .B(_05382_),
    .Y(_05384_));
 sg13g2_nor3_1 _13458_ (.A(net1900),
    .B(_05383_),
    .C(_05384_),
    .Y(_00320_));
 sg13g2_xnor2_1 _13459_ (.Y(_05385_),
    .A(net3756),
    .B(_05383_));
 sg13g2_nor2_1 _13460_ (.A(net1900),
    .B(_05385_),
    .Y(_00321_));
 sg13g2_and3_1 _13461_ (.X(_05386_),
    .A(net3068),
    .B(net4170),
    .C(_05383_));
 sg13g2_a21oi_1 _13462_ (.A1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[2] ),
    .A2(_05383_),
    .Y(_05387_),
    .B1(net3068));
 sg13g2_nor3_1 _13463_ (.A(net1900),
    .B(_05386_),
    .C(net3069),
    .Y(_00322_));
 sg13g2_and2_1 _13464_ (.A(net3350),
    .B(_05386_),
    .X(_05388_));
 sg13g2_nor2_1 _13465_ (.A(net3350),
    .B(_05386_),
    .Y(_05389_));
 sg13g2_nor3_1 _13466_ (.A(net1900),
    .B(_05388_),
    .C(net3351),
    .Y(_00323_));
 sg13g2_and2_1 _13467_ (.A(net3249),
    .B(_05388_),
    .X(_05390_));
 sg13g2_nor2_1 _13468_ (.A(net3249),
    .B(_05388_),
    .Y(_05391_));
 sg13g2_nor3_1 _13469_ (.A(net1900),
    .B(_05390_),
    .C(net3250),
    .Y(_00324_));
 sg13g2_and2_1 _13470_ (.A(net3335),
    .B(_05390_),
    .X(_05392_));
 sg13g2_nor2_1 _13471_ (.A(net3335),
    .B(_05390_),
    .Y(_05393_));
 sg13g2_nor3_1 _13472_ (.A(net1900),
    .B(_05392_),
    .C(net3336),
    .Y(_00325_));
 sg13g2_and2_1 _13473_ (.A(net3288),
    .B(_05392_),
    .X(_05394_));
 sg13g2_nor2_1 _13474_ (.A(net3288),
    .B(_05392_),
    .Y(_05395_));
 sg13g2_nor3_1 _13475_ (.A(net1900),
    .B(_05394_),
    .C(net3289),
    .Y(_00326_));
 sg13g2_and2_1 _13476_ (.A(net3307),
    .B(_05394_),
    .X(_05396_));
 sg13g2_nor2_1 _13477_ (.A(net3307),
    .B(_05394_),
    .Y(_05397_));
 sg13g2_nor3_1 _13478_ (.A(net1901),
    .B(_05396_),
    .C(net3308),
    .Y(_00327_));
 sg13g2_and2_1 _13479_ (.A(net3272),
    .B(_05396_),
    .X(_05398_));
 sg13g2_nor2_1 _13480_ (.A(net3272),
    .B(_05396_),
    .Y(_05399_));
 sg13g2_nor3_1 _13481_ (.A(net1901),
    .B(_05398_),
    .C(net3273),
    .Y(_00328_));
 sg13g2_and2_1 _13482_ (.A(net3402),
    .B(_05398_),
    .X(_05400_));
 sg13g2_nor2_1 _13483_ (.A(net3402),
    .B(_05398_),
    .Y(_05401_));
 sg13g2_nor3_1 _13484_ (.A(net1901),
    .B(_05400_),
    .C(_05401_),
    .Y(_00329_));
 sg13g2_xnor2_1 _13485_ (.Y(_05402_),
    .A(net3648),
    .B(_05400_));
 sg13g2_nor2_1 _13486_ (.A(net1901),
    .B(_05402_),
    .Y(_00330_));
 sg13g2_a21oi_1 _13487_ (.A1(\i_peripherals.i_uart.i_uart_tx.cycle_counter[11] ),
    .A2(_05400_),
    .Y(_05403_),
    .B1(net2909));
 sg13g2_nor2_1 _13488_ (.A(net1901),
    .B(net2910),
    .Y(_00331_));
 sg13g2_nand2_1 _13489_ (.Y(_05404_),
    .A(_02364_),
    .B(_05353_));
 sg13g2_nor2b_1 _13490_ (.A(net3532),
    .B_N(net3982),
    .Y(_05405_));
 sg13g2_a21oi_1 _13491_ (.A1(net2884),
    .A2(_05405_),
    .Y(_05406_),
    .B1(net3758));
 sg13g2_a21o_1 _13492_ (.A2(_05406_),
    .A1(_02362_),
    .B1(_05355_),
    .X(_05407_));
 sg13g2_nand3_1 _13493_ (.B(_05404_),
    .C(_05407_),
    .A(net2268),
    .Y(_05408_));
 sg13g2_o21ai_1 _13494_ (.B1(_05408_),
    .Y(_00332_),
    .A1(_01039_),
    .A2(_05380_));
 sg13g2_a21oi_1 _13495_ (.A1(_02364_),
    .A2(_05353_),
    .Y(_05409_),
    .B1(_05406_));
 sg13g2_o21ai_1 _13496_ (.B1(net2268),
    .Y(_05410_),
    .A1(net2884),
    .A2(_05409_));
 sg13g2_a21oi_1 _13497_ (.A1(net2884),
    .A2(_05409_),
    .Y(_00333_),
    .B1(_05410_));
 sg13g2_nor3_1 _13498_ (.A(_01038_),
    .B(_01039_),
    .C(_05353_),
    .Y(_05411_));
 sg13g2_nor2_1 _13499_ (.A(net3532),
    .B(_05411_),
    .Y(_05412_));
 sg13g2_and2_1 _13500_ (.A(net3532),
    .B(_05411_),
    .X(_05413_));
 sg13g2_nor3_1 _13501_ (.A(net2246),
    .B(net3533),
    .C(_05413_),
    .Y(_00334_));
 sg13g2_nand4_1 _13502_ (.B(_01039_),
    .C(_05404_),
    .A(net2884),
    .Y(_05414_),
    .D(_05405_));
 sg13g2_xor2_1 _13503_ (.B(_05413_),
    .A(net3982),
    .X(_05415_));
 sg13g2_and3_1 _13504_ (.X(_00335_),
    .A(net2268),
    .B(_05414_),
    .C(_05415_));
 sg13g2_nor2_1 _13505_ (.A(_00990_),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[8] ),
    .Y(_05416_));
 sg13g2_nor2_1 _13506_ (.A(_01047_),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[7] ),
    .Y(_05417_));
 sg13g2_nand2_1 _13507_ (.Y(_05418_),
    .A(_01053_),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ));
 sg13g2_nor2b_1 _13508_ (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[0] ),
    .B_N(\i_peripherals.i_uart.baud_divider[0] ),
    .Y(_05419_));
 sg13g2_nor2_1 _13509_ (.A(_01053_),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ),
    .Y(_05420_));
 sg13g2_a221oi_1 _13510_ (.B2(_05419_),
    .C1(_05420_),
    .B1(_05418_),
    .A1(\i_peripherals.i_uart.baud_divider[2] ),
    .Y(_05421_),
    .A2(_01099_));
 sg13g2_a221oi_1 _13511_ (.B2(_01051_),
    .C1(_05421_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[3] ),
    .A1(_01052_),
    .Y(_05422_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[2] ));
 sg13g2_a221oi_1 _13512_ (.B2(\i_peripherals.i_uart.baud_divider[4] ),
    .C1(_05422_),
    .B1(_01101_),
    .A1(\i_peripherals.i_uart.baud_divider[3] ),
    .Y(_05423_),
    .A2(_01100_));
 sg13g2_a21o_1 _13513_ (.A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[4] ),
    .A1(_01050_),
    .B1(_05423_),
    .X(_05424_));
 sg13g2_o21ai_1 _13514_ (.B1(_05424_),
    .Y(_05425_),
    .A1(_01049_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ));
 sg13g2_a22oi_1 _13515_ (.Y(_05426_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[6] ),
    .B2(_01048_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ),
    .A1(_01049_));
 sg13g2_a221oi_1 _13516_ (.B2(_05426_),
    .C1(_05417_),
    .B1(_05425_),
    .A1(\i_peripherals.i_uart.baud_divider[6] ),
    .Y(_05427_),
    .A2(_01102_));
 sg13g2_a221oi_1 _13517_ (.B2(_00990_),
    .C1(_05427_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[8] ),
    .A1(_01047_),
    .Y(_05428_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[7] ));
 sg13g2_nand2_1 _13518_ (.Y(_05429_),
    .A(_00989_),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[9] ));
 sg13g2_o21ai_1 _13519_ (.B1(_05429_),
    .Y(_05430_),
    .A1(_05416_),
    .A2(_05428_));
 sg13g2_a22oi_1 _13520_ (.Y(_05431_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[11] ),
    .B2(_00987_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[10] ),
    .A1(_00988_));
 sg13g2_nand2_1 _13521_ (.Y(_05432_),
    .A(\i_peripherals.i_uart.baud_divider[11] ),
    .B(_01105_));
 sg13g2_a22oi_1 _13522_ (.Y(_05433_),
    .B1(_01104_),
    .B2(\i_peripherals.i_uart.baud_divider[10] ),
    .A2(_01103_),
    .A1(\i_peripherals.i_uart.baud_divider[9] ));
 sg13g2_nand4_1 _13523_ (.B(_05431_),
    .C(_05432_),
    .A(_05430_),
    .Y(_05434_),
    .D(_05433_));
 sg13g2_nor2b_1 _13524_ (.A(_05431_),
    .B_N(_05432_),
    .Y(_05435_));
 sg13g2_a21oi_1 _13525_ (.A1(_00986_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[12] ),
    .Y(_05436_),
    .B1(_05435_));
 sg13g2_a22oi_1 _13526_ (.Y(_05437_),
    .B1(_05434_),
    .B2(_05436_),
    .A2(_01106_),
    .A1(\i_peripherals.i_uart.baud_divider[12] ));
 sg13g2_or3_1 _13527_ (.A(net3448),
    .B(net3835),
    .C(net3976),
    .X(_05438_));
 sg13g2_o21ai_1 _13528_ (.B1(\i_peripherals.i_uart.i_uart_rx.fsm_state[3] ),
    .Y(_05439_),
    .A1(\i_peripherals.i_uart.i_uart_rx.fsm_state[2] ),
    .A2(\i_peripherals.i_uart.i_uart_rx.fsm_state[1] ));
 sg13g2_nand3_1 _13529_ (.B(_05438_),
    .C(_05439_),
    .A(_05437_),
    .Y(_05440_));
 sg13g2_mux2_1 _13530_ (.A0(net3126),
    .A1(net3104),
    .S(_05440_),
    .X(_00336_));
 sg13g2_mux2_1 _13531_ (.A0(net3396),
    .A1(net3126),
    .S(_05440_),
    .X(_00337_));
 sg13g2_mux2_1 _13532_ (.A0(net3359),
    .A1(\i_peripherals.i_uart.i_uart_rx.recieved_data[2] ),
    .S(_05440_),
    .X(_00338_));
 sg13g2_mux2_1 _13533_ (.A0(net3426),
    .A1(net3359),
    .S(_05440_),
    .X(_00339_));
 sg13g2_mux2_1 _13534_ (.A0(\i_peripherals.i_uart.i_uart_rx.recieved_data[5] ),
    .A1(net3426),
    .S(_05440_),
    .X(_00340_));
 sg13g2_mux2_1 _13535_ (.A0(net3406),
    .A1(net3486),
    .S(_05440_),
    .X(_00341_));
 sg13g2_mux2_1 _13536_ (.A0(net3123),
    .A1(net3406),
    .S(_05440_),
    .X(_00342_));
 sg13g2_mux2_1 _13537_ (.A0(net2896),
    .A1(net3123),
    .S(_05440_),
    .X(_00343_));
 sg13g2_xnor2_1 _13538_ (.Y(_05441_),
    .A(\i_peripherals.i_uart.baud_divider[8] ),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[7] ));
 sg13g2_nor2b_1 _13539_ (.A(\i_peripherals.i_uart.baud_divider[1] ),
    .B_N(\i_peripherals.i_uart.i_uart_rx.cycle_counter[0] ),
    .Y(_05442_));
 sg13g2_a22oi_1 _13540_ (.Y(_05443_),
    .B1(_01101_),
    .B2(\i_peripherals.i_uart.baud_divider[5] ),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[2] ),
    .A1(_01051_));
 sg13g2_nor2_1 _13541_ (.A(_01048_),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ),
    .Y(_05444_));
 sg13g2_nor2_1 _13542_ (.A(\i_peripherals.i_uart.baud_divider[11] ),
    .B(_01104_),
    .Y(_05445_));
 sg13g2_nand2b_1 _13543_ (.Y(_05446_),
    .B(\i_peripherals.i_uart.baud_divider[9] ),
    .A_N(\i_peripherals.i_uart.i_uart_rx.cycle_counter[8] ));
 sg13g2_nor2_1 _13544_ (.A(_01053_),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[0] ),
    .Y(_05447_));
 sg13g2_a221oi_1 _13545_ (.B2(_00988_),
    .C1(_05445_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[9] ),
    .A1(_01049_),
    .Y(_05448_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[4] ));
 sg13g2_a22oi_1 _13546_ (.Y(_05449_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[8] ),
    .B2(_00989_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ),
    .A1(_01052_));
 sg13g2_o21ai_1 _13547_ (.B1(_05446_),
    .Y(_05450_),
    .A1(_01052_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ));
 sg13g2_a21oi_1 _13548_ (.A1(_01047_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[6] ),
    .Y(_05451_),
    .B1(_05450_));
 sg13g2_a221oi_1 _13549_ (.B2(\i_peripherals.i_uart.baud_divider[10] ),
    .C1(_05442_),
    .B1(_01103_),
    .A1(\i_peripherals.i_uart.baud_divider[3] ),
    .Y(_05452_),
    .A2(_01099_));
 sg13g2_and4_1 _13550_ (.A(_05448_),
    .B(_05449_),
    .C(_05451_),
    .D(_05452_),
    .X(_05453_));
 sg13g2_a22oi_1 _13551_ (.Y(_05454_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[11] ),
    .B2(_00986_),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ),
    .A1(_01048_));
 sg13g2_xnor2_1 _13552_ (.Y(_05455_),
    .A(\i_peripherals.i_uart.baud_divider[4] ),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[3] ));
 sg13g2_a22oi_1 _13553_ (.Y(_05456_),
    .B1(_01105_),
    .B2(\i_peripherals.i_uart.baud_divider[12] ),
    .A2(_01102_),
    .A1(\i_peripherals.i_uart.baud_divider[7] ));
 sg13g2_nand3_1 _13554_ (.B(_05443_),
    .C(_05456_),
    .A(_05441_),
    .Y(_05457_));
 sg13g2_a21oi_1 _13555_ (.A1(\i_peripherals.i_uart.baud_divider[11] ),
    .A2(_01104_),
    .Y(_05458_),
    .B1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[12] ));
 sg13g2_nand4_1 _13556_ (.B(_05454_),
    .C(_05455_),
    .A(_05453_),
    .Y(_05459_),
    .D(_05458_));
 sg13g2_or4_1 _13557_ (.A(_05444_),
    .B(_05447_),
    .C(_05457_),
    .D(_05459_),
    .X(_05460_));
 sg13g2_nor2b_1 _13558_ (.A(net2896),
    .B_N(_05460_),
    .Y(_05461_));
 sg13g2_mux2_1 _13559_ (.A0(\i_peripherals.i_uart.ui_in[7] ),
    .A1(\i_peripherals.i_uart.ui_in[3] ),
    .S(\i_peripherals.i_uart.rxd_select ),
    .X(_05462_));
 sg13g2_inv_1 _13560_ (.Y(_05463_),
    .A(_05462_));
 sg13g2_nor2_1 _13561_ (.A(_05460_),
    .B(_05462_),
    .Y(_05464_));
 sg13g2_nor3_1 _13562_ (.A(net2248),
    .B(_05461_),
    .C(_05464_),
    .Y(_00344_));
 sg13g2_nor2_2 _13563_ (.A(\i_peripherals.i_uart.uart_rx_buffered ),
    .B(net2248),
    .Y(_05465_));
 sg13g2_a21o_1 _13564_ (.A2(_05438_),
    .A1(net4088),
    .B1(net2248),
    .X(_00345_));
 sg13g2_nor2_1 _13565_ (.A(net2481),
    .B(_05438_),
    .Y(_05466_));
 sg13g2_nor2_1 _13566_ (.A(_05325_),
    .B(_05466_),
    .Y(_05467_));
 sg13g2_nand2b_2 _13567_ (.Y(_05468_),
    .B(_05467_),
    .A_N(_05437_));
 sg13g2_nand2_1 _13568_ (.Y(_05469_),
    .A(net2481),
    .B(_05326_));
 sg13g2_nor4_1 _13569_ (.A(net2481),
    .B(_05326_),
    .C(_05460_),
    .D(_05463_),
    .Y(_05470_));
 sg13g2_nand3_1 _13570_ (.B(\i_peripherals.i_uart.uart_rx_buffered ),
    .C(_05325_),
    .A(net2481),
    .Y(_05471_));
 sg13g2_a21oi_1 _13571_ (.A1(_05463_),
    .A2(_05466_),
    .Y(_05472_),
    .B1(_05467_));
 sg13g2_nand2_1 _13572_ (.Y(_05473_),
    .A(_05471_),
    .B(_05472_));
 sg13g2_o21ai_1 _13573_ (.B1(_05469_),
    .Y(_05474_),
    .A1(_05470_),
    .A2(_05473_));
 sg13g2_o21ai_1 _13574_ (.B1(net2274),
    .Y(_05475_),
    .A1(_05468_),
    .A2(_05474_));
 sg13g2_a21oi_1 _13575_ (.A1(_05468_),
    .A2(_05474_),
    .Y(_00346_),
    .B1(_05475_));
 sg13g2_or3_1 _13576_ (.A(net4023),
    .B(_05326_),
    .C(_05464_),
    .X(_05476_));
 sg13g2_nand3_1 _13577_ (.B(_05471_),
    .C(_05476_),
    .A(_05468_),
    .Y(_05477_));
 sg13g2_xor2_1 _13578_ (.B(net4023),
    .A(net3976),
    .X(_05478_));
 sg13g2_a21oi_1 _13579_ (.A1(_05326_),
    .A2(_05478_),
    .Y(_05479_),
    .B1(_05477_));
 sg13g2_o21ai_1 _13580_ (.B1(net2274),
    .Y(_05480_),
    .A1(net3976),
    .A2(_05468_));
 sg13g2_nor2_1 _13581_ (.A(_05479_),
    .B(_05480_),
    .Y(_00347_));
 sg13g2_nand3_1 _13582_ (.B(net2481),
    .C(_05437_),
    .A(\i_peripherals.i_uart.i_uart_rx.fsm_state[1] ),
    .Y(_05481_));
 sg13g2_xor2_1 _13583_ (.B(_05481_),
    .A(net3835),
    .X(_05482_));
 sg13g2_nor4_1 _13584_ (.A(net2248),
    .B(_05325_),
    .C(_05466_),
    .D(net3836),
    .Y(_00348_));
 sg13g2_a21oi_1 _13585_ (.A1(net3976),
    .A2(net2481),
    .Y(_05483_),
    .B1(net3448));
 sg13g2_nor2_1 _13586_ (.A(_05324_),
    .B(_05483_),
    .Y(_05484_));
 sg13g2_a21oi_1 _13587_ (.A1(net3977),
    .A2(_05484_),
    .Y(_05485_),
    .B1(_05477_));
 sg13g2_o21ai_1 _13588_ (.B1(net2274),
    .Y(_05486_),
    .A1(net3448),
    .A2(_05468_));
 sg13g2_nor2_1 _13589_ (.A(net3978),
    .B(_05486_),
    .Y(_00349_));
 sg13g2_mux2_1 _13590_ (.A0(\i_peripherals.i_uart.uart_rx_buf_data[0] ),
    .A1(net3104),
    .S(_05465_),
    .X(_00350_));
 sg13g2_mux2_1 _13591_ (.A0(net3144),
    .A1(net3126),
    .S(_05465_),
    .X(_00351_));
 sg13g2_mux2_1 _13592_ (.A0(net3252),
    .A1(\i_peripherals.i_uart.i_uart_rx.recieved_data[2] ),
    .S(_05465_),
    .X(_00352_));
 sg13g2_mux2_1 _13593_ (.A0(net3297),
    .A1(\i_peripherals.i_uart.i_uart_rx.recieved_data[3] ),
    .S(_05465_),
    .X(_00353_));
 sg13g2_mux2_1 _13594_ (.A0(net3247),
    .A1(\i_peripherals.i_uart.i_uart_rx.recieved_data[4] ),
    .S(_05465_),
    .X(_00354_));
 sg13g2_mux2_1 _13595_ (.A0(net3178),
    .A1(\i_peripherals.i_uart.i_uart_rx.recieved_data[5] ),
    .S(_05465_),
    .X(_00355_));
 sg13g2_mux2_1 _13596_ (.A0(net3415),
    .A1(net3406),
    .S(_05465_),
    .X(_00356_));
 sg13g2_mux2_1 _13597_ (.A0(net3356),
    .A1(net3123),
    .S(_05465_),
    .X(_00357_));
 sg13g2_nand2_1 _13598_ (.Y(_05487_),
    .A(net2274),
    .B(_05328_));
 sg13g2_or3_1 _13599_ (.A(_05437_),
    .B(_05466_),
    .C(_05487_),
    .X(_05488_));
 sg13g2_nor2_1 _13600_ (.A(net2750),
    .B(net1893),
    .Y(_00358_));
 sg13g2_xnor2_1 _13601_ (.Y(_05489_),
    .A(net2750),
    .B(net3775));
 sg13g2_nor2_1 _13602_ (.A(net1893),
    .B(_05489_),
    .Y(_00359_));
 sg13g2_and3_1 _13603_ (.X(_05490_),
    .A(net2750),
    .B(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ),
    .C(net2974));
 sg13g2_a21oi_1 _13604_ (.A1(net2750),
    .A2(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ),
    .Y(_05491_),
    .B1(net2974));
 sg13g2_nor3_1 _13605_ (.A(net1893),
    .B(_05490_),
    .C(net2975),
    .Y(_00360_));
 sg13g2_and2_1 _13606_ (.A(net3568),
    .B(_05490_),
    .X(_05492_));
 sg13g2_nor2_1 _13607_ (.A(net3568),
    .B(_05490_),
    .Y(_05493_));
 sg13g2_nor3_1 _13608_ (.A(net1893),
    .B(_05492_),
    .C(net3569),
    .Y(_00361_));
 sg13g2_and2_1 _13609_ (.A(net3518),
    .B(_05492_),
    .X(_05494_));
 sg13g2_nor2_1 _13610_ (.A(net3518),
    .B(_05492_),
    .Y(_05495_));
 sg13g2_nor3_1 _13611_ (.A(net1893),
    .B(_05494_),
    .C(net3519),
    .Y(_00362_));
 sg13g2_xnor2_1 _13612_ (.Y(_05496_),
    .A(net3867),
    .B(_05494_));
 sg13g2_nor2_1 _13613_ (.A(net1893),
    .B(_05496_),
    .Y(_00363_));
 sg13g2_a21oi_1 _13614_ (.A1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ),
    .A2(_05494_),
    .Y(_05497_),
    .B1(net3191));
 sg13g2_and3_1 _13615_ (.X(_05498_),
    .A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ),
    .B(net3191),
    .C(_05494_));
 sg13g2_nor3_1 _13616_ (.A(net1893),
    .B(net3192),
    .C(_05498_),
    .Y(_00364_));
 sg13g2_nor2_1 _13617_ (.A(net3751),
    .B(_05498_),
    .Y(_05499_));
 sg13g2_and2_1 _13618_ (.A(net3751),
    .B(_05498_),
    .X(_05500_));
 sg13g2_nor3_1 _13619_ (.A(net1893),
    .B(net3752),
    .C(_05500_),
    .Y(_00365_));
 sg13g2_and2_1 _13620_ (.A(net3534),
    .B(_05500_),
    .X(_05501_));
 sg13g2_nor2_1 _13621_ (.A(net3534),
    .B(_05500_),
    .Y(_05502_));
 sg13g2_nor3_1 _13622_ (.A(net1894),
    .B(_05501_),
    .C(net3535),
    .Y(_00366_));
 sg13g2_xnor2_1 _13623_ (.Y(_05503_),
    .A(net3770),
    .B(_05501_));
 sg13g2_nor2_1 _13624_ (.A(net1894),
    .B(_05503_),
    .Y(_00367_));
 sg13g2_and3_2 _13625_ (.X(_05504_),
    .A(net3770),
    .B(net3015),
    .C(_05501_));
 sg13g2_a21oi_1 _13626_ (.A1(\i_peripherals.i_uart.i_uart_rx.cycle_counter[9] ),
    .A2(_05501_),
    .Y(_05505_),
    .B1(net3015));
 sg13g2_nor3_1 _13627_ (.A(net1894),
    .B(_05504_),
    .C(net3016),
    .Y(_00368_));
 sg13g2_nand2_1 _13628_ (.Y(_05506_),
    .A(net3740),
    .B(_05504_));
 sg13g2_xnor2_1 _13629_ (.Y(_05507_),
    .A(net3740),
    .B(_05504_));
 sg13g2_nor2_1 _13630_ (.A(net1894),
    .B(net3741),
    .Y(_00369_));
 sg13g2_xnor2_1 _13631_ (.Y(_05508_),
    .A(_01106_),
    .B(_05506_));
 sg13g2_nor2_1 _13632_ (.A(net1894),
    .B(_05508_),
    .Y(_00370_));
 sg13g2_nor2_2 _13633_ (.A(\addr[7] ),
    .B(_05308_),
    .Y(_05509_));
 sg13g2_nand2b_2 _13634_ (.Y(_05510_),
    .B(_00941_),
    .A_N(_05308_));
 sg13g2_nor2_1 _13635_ (.A(_02430_),
    .B(_05510_),
    .Y(_05511_));
 sg13g2_nand2_1 _13636_ (.Y(_05512_),
    .A(_02429_),
    .B(net2158));
 sg13g2_nand2_2 _13637_ (.Y(_05513_),
    .A(net2173),
    .B(_05511_));
 sg13g2_o21ai_1 _13638_ (.B1(net2267),
    .Y(_05514_),
    .A1(net2399),
    .A2(net2015));
 sg13g2_a21oi_1 _13639_ (.A1(_01037_),
    .A2(net2015),
    .Y(_00371_),
    .B1(_05514_));
 sg13g2_o21ai_1 _13640_ (.B1(net2268),
    .Y(_05515_),
    .A1(net2398),
    .A2(net2016));
 sg13g2_a21oi_1 _13641_ (.A1(_01036_),
    .A2(net2016),
    .Y(_00372_),
    .B1(_05515_));
 sg13g2_o21ai_1 _13642_ (.B1(net2266),
    .Y(_05516_),
    .A1(net2396),
    .A2(net2015));
 sg13g2_a21oi_1 _13643_ (.A1(_01035_),
    .A2(net2015),
    .Y(_00373_),
    .B1(_05516_));
 sg13g2_o21ai_1 _13644_ (.B1(net2268),
    .Y(_05517_),
    .A1(net2394),
    .A2(net2016));
 sg13g2_a21oi_1 _13645_ (.A1(_01034_),
    .A2(net2016),
    .Y(_00374_),
    .B1(_05517_));
 sg13g2_o21ai_1 _13646_ (.B1(net2265),
    .Y(_05518_),
    .A1(net2392),
    .A2(net2015));
 sg13g2_a21oi_1 _13647_ (.A1(_01033_),
    .A2(net2015),
    .Y(_00375_),
    .B1(_05518_));
 sg13g2_o21ai_1 _13648_ (.B1(net2266),
    .Y(_05519_),
    .A1(net2389),
    .A2(net2015));
 sg13g2_a21oi_1 _13649_ (.A1(_01032_),
    .A2(net2015),
    .Y(_00376_),
    .B1(_05519_));
 sg13g2_o21ai_1 _13650_ (.B1(net2270),
    .Y(_05520_),
    .A1(\data_to_write[6] ),
    .A2(net2016));
 sg13g2_a21oi_1 _13651_ (.A1(_01031_),
    .A2(net2016),
    .Y(_00377_),
    .B1(_05520_));
 sg13g2_o21ai_1 _13652_ (.B1(net2272),
    .Y(_05521_),
    .A1(\data_to_write[7] ),
    .A2(net2016));
 sg13g2_a21oi_1 _13653_ (.A1(_01030_),
    .A2(net2016),
    .Y(_00378_),
    .B1(_05521_));
 sg13g2_nor3_2 _13654_ (.A(net2385),
    .B(_02430_),
    .C(_05174_),
    .Y(_05522_));
 sg13g2_nand3_1 _13655_ (.B(net2158),
    .C(_05522_),
    .A(_05216_),
    .Y(_05523_));
 sg13g2_nand3_1 _13656_ (.B(net2158),
    .C(_05522_),
    .A(_05216_),
    .Y(_05524_));
 sg13g2_o21ai_1 _13657_ (.B1(net2265),
    .Y(_05525_),
    .A1(net2399),
    .A2(net2014));
 sg13g2_a21oi_1 _13658_ (.A1(_01029_),
    .A2(net2014),
    .Y(_00379_),
    .B1(_05525_));
 sg13g2_a21oi_1 _13659_ (.A1(net3417),
    .A2(net2014),
    .Y(_05526_),
    .B1(net2247));
 sg13g2_o21ai_1 _13660_ (.B1(_05526_),
    .Y(_00380_),
    .A1(_00973_),
    .A2(_05523_));
 sg13g2_o21ai_1 _13661_ (.B1(net2265),
    .Y(_05527_),
    .A1(net2396),
    .A2(_05524_));
 sg13g2_a21oi_1 _13662_ (.A1(_01028_),
    .A2(net2014),
    .Y(_00381_),
    .B1(_05527_));
 sg13g2_o21ai_1 _13663_ (.B1(net2265),
    .Y(_05528_),
    .A1(net2394),
    .A2(net2014));
 sg13g2_a21oi_1 _13664_ (.A1(_01027_),
    .A2(_05524_),
    .Y(_00382_),
    .B1(_05528_));
 sg13g2_o21ai_1 _13665_ (.B1(net2265),
    .Y(_05529_),
    .A1(net2392),
    .A2(net2014));
 sg13g2_a21oi_1 _13666_ (.A1(_01026_),
    .A2(_05524_),
    .Y(_00383_),
    .B1(_05529_));
 sg13g2_o21ai_1 _13667_ (.B1(net2265),
    .Y(_05530_),
    .A1(net2390),
    .A2(net2014));
 sg13g2_a21oi_1 _13668_ (.A1(_01025_),
    .A2(net2014),
    .Y(_00384_),
    .B1(_05530_));
 sg13g2_nor4_2 _13669_ (.A(net3331),
    .B(_02613_),
    .C(net2041),
    .Y(_05531_),
    .D(_05320_));
 sg13g2_nand3b_1 _13670_ (.B(net2038),
    .C(_05321_),
    .Y(_05532_),
    .A_N(net3331));
 sg13g2_a21oi_1 _13671_ (.A1(\i_peripherals.i_user_peri39._GEN[32] ),
    .A2(net2170),
    .Y(_05533_),
    .B1(net2093));
 sg13g2_and4_1 _13672_ (.A(_00943_),
    .B(net2385),
    .C(_01921_),
    .D(_05216_),
    .X(_05534_));
 sg13g2_nand2_1 _13673_ (.Y(_05535_),
    .A(\i_peripherals.i_user_peri39._GEN[64] ),
    .B(net2191));
 sg13g2_a22oi_1 _13674_ (.Y(_05536_),
    .B1(net2162),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[0] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[0] ));
 sg13g2_nand3_1 _13675_ (.B(_05535_),
    .C(_05536_),
    .A(_05533_),
    .Y(_05537_));
 sg13g2_o21ai_1 _13676_ (.B1(_05537_),
    .Y(_05538_),
    .A1(\i_peripherals.i_user_peri39.instr[0] ),
    .A2(net2089));
 sg13g2_a22oi_1 _13677_ (.Y(_05539_),
    .B1(_05329_),
    .B2(\i_peripherals.i_uart.rxd_select ),
    .A2(net2165),
    .A1(\i_peripherals.i_uart.baud_divider[0] ));
 sg13g2_nand2b_1 _13678_ (.Y(_05540_),
    .B(_05539_),
    .A_N(net2167));
 sg13g2_nand2b_1 _13679_ (.Y(_05541_),
    .B(_05309_),
    .A_N(net2174));
 sg13g2_a21oi_1 _13680_ (.A1(_02363_),
    .A2(net2167),
    .Y(_05542_),
    .B1(_05541_));
 sg13g2_a221oi_1 _13681_ (.B2(_05542_),
    .C1(net2159),
    .B1(_05540_),
    .A1(\i_peripherals.i_uart.uart_rx_buf_data[0] ),
    .Y(_05543_),
    .A2(net2081));
 sg13g2_o21ai_1 _13682_ (.B1(_05543_),
    .Y(_05544_),
    .A1(net2195),
    .A2(_05538_));
 sg13g2_a221oi_1 _13683_ (.B2(\i_peripherals.i_uart.ui_in[0] ),
    .C1(_05510_),
    .B1(net2166),
    .A1(net3054),
    .Y(_05545_),
    .A2(net2173));
 sg13g2_inv_1 _13684_ (.Y(_05546_),
    .A(_05545_));
 sg13g2_a21oi_1 _13685_ (.A1(_05544_),
    .A2(_05546_),
    .Y(_05547_),
    .B1(net1980));
 sg13g2_o21ai_1 _13686_ (.B1(net2270),
    .Y(_05548_),
    .A1(net3625),
    .A2(net1986));
 sg13g2_nor2_1 _13687_ (.A(_05547_),
    .B(_05548_),
    .Y(_00385_));
 sg13g2_a21oi_1 _13688_ (.A1(\i_peripherals.i_user_peri39._GEN[1] ),
    .A2(net2177),
    .Y(_05549_),
    .B1(net2093));
 sg13g2_nand2_1 _13689_ (.Y(_05550_),
    .A(\i_peripherals.i_user_peri39._GEN[65] ),
    .B(net2191));
 sg13g2_a22oi_1 _13690_ (.Y(_05551_),
    .B1(net2161),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[1] ),
    .A2(net2169),
    .A1(\i_peripherals.i_user_peri39._GEN[33] ));
 sg13g2_nand3_1 _13691_ (.B(_05550_),
    .C(_05551_),
    .A(_05549_),
    .Y(_05552_));
 sg13g2_o21ai_1 _13692_ (.B1(_05552_),
    .Y(_05553_),
    .A1(\i_peripherals.i_user_peri39.instr[1] ),
    .A2(net2088));
 sg13g2_a22oi_1 _13693_ (.Y(_05554_),
    .B1(net2165),
    .B2(\i_peripherals.i_uart.baud_divider[1] ),
    .A2(net2167),
    .A1(\i_peripherals.i_uart.uart_rx_buffered ));
 sg13g2_o21ai_1 _13694_ (.B1(_05510_),
    .Y(_05555_),
    .A1(_05541_),
    .A2(_05554_));
 sg13g2_a21oi_1 _13695_ (.A1(net3144),
    .A2(net2081),
    .Y(_05556_),
    .B1(_05555_));
 sg13g2_o21ai_1 _13696_ (.B1(_05556_),
    .Y(_05557_),
    .A1(net2195),
    .A2(_05553_));
 sg13g2_a221oi_1 _13697_ (.B2(\i_peripherals.i_uart.ui_in[1] ),
    .C1(_05510_),
    .B1(net2166),
    .A1(\i_peripherals.gpio_out[1] ),
    .Y(_05558_),
    .A2(net2173));
 sg13g2_nor2_1 _13698_ (.A(net1980),
    .B(_05558_),
    .Y(_05559_));
 sg13g2_a22oi_1 _13699_ (.Y(_05560_),
    .B1(_05557_),
    .B2(_05559_),
    .A2(net1985),
    .A1(net3271));
 sg13g2_nor2_1 _13700_ (.A(net2248),
    .B(_05560_),
    .Y(_00386_));
 sg13g2_a21oi_1 _13701_ (.A1(\i_peripherals.i_user_peri39.math_result_reg[2] ),
    .A2(net2161),
    .Y(_05561_),
    .B1(net2093));
 sg13g2_nand2_1 _13702_ (.Y(_05562_),
    .A(\i_peripherals.i_user_peri39._GEN[66] ),
    .B(net2191));
 sg13g2_a22oi_1 _13703_ (.Y(_05563_),
    .B1(net2169),
    .B2(\i_peripherals.i_user_peri39._GEN[34] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[2] ));
 sg13g2_nand3_1 _13704_ (.B(_05562_),
    .C(_05563_),
    .A(_05561_),
    .Y(_05564_));
 sg13g2_o21ai_1 _13705_ (.B1(_05564_),
    .Y(_05565_),
    .A1(\i_peripherals.i_user_peri39.instr[2] ),
    .A2(net2088));
 sg13g2_a221oi_1 _13706_ (.B2(net3252),
    .C1(net2159),
    .B1(net2081),
    .A1(\i_peripherals.i_uart.baud_divider[2] ),
    .Y(_05566_),
    .A2(net2085));
 sg13g2_o21ai_1 _13707_ (.B1(_05566_),
    .Y(_05567_),
    .A1(net2195),
    .A2(_05565_));
 sg13g2_a22oi_1 _13708_ (.Y(_05568_),
    .B1(net2166),
    .B2(\i_peripherals.i_uart.ui_in[2] ),
    .A2(net2173),
    .A1(\i_peripherals.gpio_out[2] ));
 sg13g2_nand2_1 _13709_ (.Y(_05569_),
    .A(_05509_),
    .B(_05568_));
 sg13g2_a21oi_1 _13710_ (.A1(_05567_),
    .A2(_05569_),
    .Y(_05570_),
    .B1(net1985));
 sg13g2_o21ai_1 _13711_ (.B1(net2274),
    .Y(_05571_),
    .A1(net3477),
    .A2(net1986));
 sg13g2_nor2_1 _13712_ (.A(_05570_),
    .B(_05571_),
    .Y(_00387_));
 sg13g2_a21oi_1 _13713_ (.A1(\i_peripherals.i_user_peri39._GEN[35] ),
    .A2(net2169),
    .Y(_05572_),
    .B1(net2093));
 sg13g2_nand2_1 _13714_ (.Y(_05573_),
    .A(\i_peripherals.i_user_peri39._GEN[67] ),
    .B(net2191));
 sg13g2_a22oi_1 _13715_ (.Y(_05574_),
    .B1(net2161),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[3] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[3] ));
 sg13g2_nand3_1 _13716_ (.B(_05573_),
    .C(_05574_),
    .A(_05572_),
    .Y(_05575_));
 sg13g2_o21ai_1 _13717_ (.B1(_05575_),
    .Y(_05576_),
    .A1(\i_peripherals.i_user_peri39.instr[3] ),
    .A2(net2088));
 sg13g2_a221oi_1 _13718_ (.B2(net3297),
    .C1(net2159),
    .B1(net2081),
    .A1(\i_peripherals.i_uart.baud_divider[3] ),
    .Y(_05577_),
    .A2(net2085));
 sg13g2_o21ai_1 _13719_ (.B1(_05577_),
    .Y(_05578_),
    .A1(net2195),
    .A2(_05576_));
 sg13g2_a221oi_1 _13720_ (.B2(\i_peripherals.i_uart.ui_in[3] ),
    .C1(_05510_),
    .B1(net2166),
    .A1(\i_peripherals.gpio_out[3] ),
    .Y(_05579_),
    .A2(net2173));
 sg13g2_nor2_1 _13721_ (.A(net1985),
    .B(_05579_),
    .Y(_05580_));
 sg13g2_a22oi_1 _13722_ (.Y(_05581_),
    .B1(_05578_),
    .B2(_05580_),
    .A2(net1985),
    .A1(net3573));
 sg13g2_nor2_1 _13723_ (.A(net2249),
    .B(net3574),
    .Y(_00388_));
 sg13g2_a21oi_1 _13724_ (.A1(\i_peripherals.i_user_peri39._GEN[36] ),
    .A2(net2171),
    .Y(_05582_),
    .B1(net2095));
 sg13g2_nand2_1 _13725_ (.Y(_05583_),
    .A(\i_peripherals.i_user_peri39._GEN[68] ),
    .B(net2191));
 sg13g2_a22oi_1 _13726_ (.Y(_05584_),
    .B1(net2162),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[4] ),
    .A2(net2178),
    .A1(\i_peripherals.i_user_peri39._GEN[100] ));
 sg13g2_nand3_1 _13727_ (.B(_05583_),
    .C(_05584_),
    .A(_05582_),
    .Y(_05585_));
 sg13g2_o21ai_1 _13728_ (.B1(_05585_),
    .Y(_05586_),
    .A1(\i_peripherals.i_user_peri39.instr[4] ),
    .A2(net2088));
 sg13g2_a221oi_1 _13729_ (.B2(net3247),
    .C1(net2159),
    .B1(net2081),
    .A1(\i_peripherals.i_uart.baud_divider[4] ),
    .Y(_05587_),
    .A2(net2085));
 sg13g2_o21ai_1 _13730_ (.B1(_05587_),
    .Y(_05588_),
    .A1(net2196),
    .A2(_05586_));
 sg13g2_a221oi_1 _13731_ (.B2(\i_peripherals.i_uart.ui_in[4] ),
    .C1(_05510_),
    .B1(net2166),
    .A1(net3136),
    .Y(_05589_),
    .A2(net2173));
 sg13g2_nor2_1 _13732_ (.A(net1980),
    .B(_05589_),
    .Y(_05590_));
 sg13g2_a22oi_1 _13733_ (.Y(_05591_),
    .B1(_05588_),
    .B2(_05590_),
    .A2(net1980),
    .A1(net3419));
 sg13g2_nor2_1 _13734_ (.A(net2246),
    .B(net3420),
    .Y(_00389_));
 sg13g2_a21oi_1 _13735_ (.A1(\i_peripherals.i_user_peri39.math_result_reg[5] ),
    .A2(net2161),
    .Y(_05592_),
    .B1(net2093));
 sg13g2_nand2_1 _13736_ (.Y(_05593_),
    .A(\i_peripherals.i_user_peri39._GEN[69] ),
    .B(net2192));
 sg13g2_a22oi_1 _13737_ (.Y(_05594_),
    .B1(net2169),
    .B2(\i_peripherals.i_user_peri39._GEN[37] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[101] ));
 sg13g2_nand3_1 _13738_ (.B(_05593_),
    .C(_05594_),
    .A(_05592_),
    .Y(_05595_));
 sg13g2_o21ai_1 _13739_ (.B1(_05595_),
    .Y(_05596_),
    .A1(\i_peripherals.i_user_peri39.instr[5] ),
    .A2(net2088));
 sg13g2_a221oi_1 _13740_ (.B2(net3178),
    .C1(net2159),
    .B1(net2081),
    .A1(\i_peripherals.i_uart.baud_divider[5] ),
    .Y(_05597_),
    .A2(net2085));
 sg13g2_o21ai_1 _13741_ (.B1(_05597_),
    .Y(_05598_),
    .A1(net2195),
    .A2(_05596_));
 sg13g2_a221oi_1 _13742_ (.B2(\i_peripherals.i_uart.ui_in[5] ),
    .C1(_05510_),
    .B1(net2166),
    .A1(\i_peripherals.gpio_out[5] ),
    .Y(_05599_),
    .A2(net2173));
 sg13g2_nor2_1 _13743_ (.A(net1985),
    .B(_05599_),
    .Y(_05600_));
 sg13g2_a22oi_1 _13744_ (.Y(_05601_),
    .B1(_05598_),
    .B2(_05600_),
    .A2(net1980),
    .A1(net3194));
 sg13g2_nor2_1 _13745_ (.A(net2248),
    .B(net3195),
    .Y(_00390_));
 sg13g2_a21oi_1 _13746_ (.A1(\i_peripherals.i_user_peri39._GEN[38] ),
    .A2(net2168),
    .Y(_05602_),
    .B1(net2092));
 sg13g2_nand2_1 _13747_ (.Y(_05603_),
    .A(\i_peripherals.i_user_peri39._GEN[70] ),
    .B(net2191));
 sg13g2_a22oi_1 _13748_ (.Y(_05604_),
    .B1(net2162),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[6] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[102] ));
 sg13g2_nand3_1 _13749_ (.B(_05603_),
    .C(_05604_),
    .A(_05602_),
    .Y(_05605_));
 sg13g2_o21ai_1 _13750_ (.B1(_05605_),
    .Y(_05606_),
    .A1(\i_peripherals.i_user_peri39.instr[6] ),
    .A2(net2088));
 sg13g2_a221oi_1 _13751_ (.B2(\i_peripherals.i_uart.uart_rx_buf_data[6] ),
    .C1(_05509_),
    .B1(_05322_),
    .A1(\i_peripherals.i_uart.baud_divider[6] ),
    .Y(_05607_),
    .A2(net2085));
 sg13g2_o21ai_1 _13752_ (.B1(_05607_),
    .Y(_05608_),
    .A1(net2195),
    .A2(_05606_));
 sg13g2_a22oi_1 _13753_ (.Y(_05609_),
    .B1(net2166),
    .B2(\i_peripherals.i_uart.ui_in[6] ),
    .A2(net2173),
    .A1(net3187));
 sg13g2_nand2_1 _13754_ (.Y(_05610_),
    .A(net2159),
    .B(_05609_));
 sg13g2_a21oi_1 _13755_ (.A1(_05608_),
    .A2(_05610_),
    .Y(_05611_),
    .B1(net1980));
 sg13g2_o21ai_1 _13756_ (.B1(net2270),
    .Y(_05612_),
    .A1(net3474),
    .A2(net1986));
 sg13g2_nor2_1 _13757_ (.A(_05611_),
    .B(_05612_),
    .Y(_00391_));
 sg13g2_a21oi_1 _13758_ (.A1(\i_peripherals.i_user_peri39.math_result_reg[7] ),
    .A2(net2162),
    .Y(_05613_),
    .B1(net2095));
 sg13g2_nand2_1 _13759_ (.Y(_05614_),
    .A(\i_peripherals.i_user_peri39._GEN[71] ),
    .B(net2190));
 sg13g2_a22oi_1 _13760_ (.Y(_05615_),
    .B1(net2168),
    .B2(\i_peripherals.i_user_peri39._GEN[39] ),
    .A2(net2175),
    .A1(\i_peripherals.i_user_peri39._GEN[103] ));
 sg13g2_nand3_1 _13761_ (.B(_05614_),
    .C(_05615_),
    .A(_05613_),
    .Y(_05616_));
 sg13g2_o21ai_1 _13762_ (.B1(_05616_),
    .Y(_05617_),
    .A1(\i_peripherals.i_user_peri39.instr[7] ),
    .A2(net2087));
 sg13g2_a221oi_1 _13763_ (.B2(\i_peripherals.i_uart.uart_rx_buf_data[7] ),
    .C1(net2159),
    .B1(_05322_),
    .A1(\i_peripherals.i_uart.baud_divider[7] ),
    .Y(_05618_),
    .A2(net2085));
 sg13g2_o21ai_1 _13764_ (.B1(_05618_),
    .Y(_05619_),
    .A1(net2195),
    .A2(_05617_));
 sg13g2_a221oi_1 _13765_ (.B2(\i_peripherals.i_uart.ui_in[7] ),
    .C1(_05510_),
    .B1(net2166),
    .A1(net2946),
    .Y(_05620_),
    .A2(net2174));
 sg13g2_nor2_1 _13766_ (.A(net1980),
    .B(_05620_),
    .Y(_05621_));
 sg13g2_a22oi_1 _13767_ (.Y(_05622_),
    .B1(_05619_),
    .B2(_05621_),
    .A2(net1980),
    .A1(net3333));
 sg13g2_nor2_1 _13768_ (.A(net2246),
    .B(net3334),
    .Y(_00392_));
 sg13g2_a21oi_1 _13769_ (.A1(\i_peripherals.i_user_peri39.math_result_reg[8] ),
    .A2(net2161),
    .Y(_05623_),
    .B1(net2093));
 sg13g2_nand2_1 _13770_ (.Y(_05624_),
    .A(\i_peripherals.i_user_peri39._GEN[72] ),
    .B(net2192));
 sg13g2_a22oi_1 _13771_ (.Y(_05625_),
    .B1(net2169),
    .B2(\i_peripherals.i_user_peri39._GEN[40] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[104] ));
 sg13g2_nand3_1 _13772_ (.B(_05624_),
    .C(_05625_),
    .A(_05623_),
    .Y(_05626_));
 sg13g2_a21oi_1 _13773_ (.A1(_01062_),
    .A2(net2090),
    .Y(_05627_),
    .B1(net2196));
 sg13g2_a221oi_1 _13774_ (.B2(_05627_),
    .C1(net1984),
    .B1(_05626_),
    .A1(\i_peripherals.i_uart.baud_divider[8] ),
    .Y(_05628_),
    .A2(net2085));
 sg13g2_o21ai_1 _13775_ (.B1(net2274),
    .Y(_05629_),
    .A1(net3352),
    .A2(net1986));
 sg13g2_nor2_1 _13776_ (.A(_05628_),
    .B(_05629_),
    .Y(_00393_));
 sg13g2_a21oi_1 _13777_ (.A1(net2970),
    .A2(net2172),
    .Y(_05630_),
    .B1(net2090));
 sg13g2_nand2_1 _13778_ (.Y(_05631_),
    .A(net3582),
    .B(net2190));
 sg13g2_a22oi_1 _13779_ (.Y(_05632_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[9] ),
    .A2(net2179),
    .A1(net2993));
 sg13g2_nand3_1 _13780_ (.B(_05631_),
    .C(_05632_),
    .A(_05630_),
    .Y(_05633_));
 sg13g2_a21oi_1 _13781_ (.A1(_01061_),
    .A2(net2090),
    .Y(_05634_),
    .B1(net2196));
 sg13g2_a221oi_1 _13782_ (.B2(_05634_),
    .C1(net1984),
    .B1(_05633_),
    .A1(\i_peripherals.i_uart.baud_divider[9] ),
    .Y(_05635_),
    .A2(net2086));
 sg13g2_o21ai_1 _13783_ (.B1(net2275),
    .Y(_05636_),
    .A1(net3738),
    .A2(net1986));
 sg13g2_nor2_1 _13784_ (.A(_05635_),
    .B(_05636_),
    .Y(_00394_));
 sg13g2_a21oi_1 _13785_ (.A1(\i_peripherals.i_user_peri39._GEN[42] ),
    .A2(net2169),
    .Y(_05637_),
    .B1(net2094));
 sg13g2_nand2_1 _13786_ (.Y(_05638_),
    .A(\i_peripherals.i_user_peri39._GEN[74] ),
    .B(net2192));
 sg13g2_a22oi_1 _13787_ (.Y(_05639_),
    .B1(net2161),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[10] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[106] ));
 sg13g2_nand3_1 _13788_ (.B(_05638_),
    .C(_05639_),
    .A(_05637_),
    .Y(_05640_));
 sg13g2_a21oi_1 _13789_ (.A1(_01060_),
    .A2(net2090),
    .Y(_05641_),
    .B1(net2196));
 sg13g2_a221oi_1 _13790_ (.B2(_05641_),
    .C1(net1984),
    .B1(_05640_),
    .A1(\i_peripherals.i_uart.baud_divider[10] ),
    .Y(_05642_),
    .A2(net2086));
 sg13g2_o21ai_1 _13791_ (.B1(net2275),
    .Y(_05643_),
    .A1(net3605),
    .A2(net1986));
 sg13g2_nor2_1 _13792_ (.A(_05642_),
    .B(_05643_),
    .Y(_00395_));
 sg13g2_a21oi_1 _13793_ (.A1(\i_peripherals.i_user_peri39.math_result_reg[11] ),
    .A2(net2161),
    .Y(_05644_),
    .B1(net2093));
 sg13g2_nand2_1 _13794_ (.Y(_05645_),
    .A(\i_peripherals.i_user_peri39._GEN[75] ),
    .B(net2192));
 sg13g2_a22oi_1 _13795_ (.Y(_05646_),
    .B1(net2169),
    .B2(\i_peripherals.i_user_peri39._GEN[43] ),
    .A2(net2178),
    .A1(\i_peripherals.i_user_peri39._GEN[107] ));
 sg13g2_nand3_1 _13796_ (.B(_05645_),
    .C(_05646_),
    .A(_05644_),
    .Y(_05647_));
 sg13g2_a21oi_1 _13797_ (.A1(_01059_),
    .A2(net2090),
    .Y(_05648_),
    .B1(net2196));
 sg13g2_a221oi_1 _13798_ (.B2(_05648_),
    .C1(net1984),
    .B1(_05647_),
    .A1(\i_peripherals.i_uart.baud_divider[11] ),
    .Y(_05649_),
    .A2(net2086));
 sg13g2_o21ai_1 _13799_ (.B1(net2275),
    .Y(_05650_),
    .A1(net3822),
    .A2(net1986));
 sg13g2_nor2_1 _13800_ (.A(_05649_),
    .B(_05650_),
    .Y(_00396_));
 sg13g2_a21oi_1 _13801_ (.A1(\i_peripherals.i_user_peri39.math_result_reg[12] ),
    .A2(net2161),
    .Y(_05651_),
    .B1(net2093));
 sg13g2_nand2_1 _13802_ (.Y(_05652_),
    .A(\i_peripherals.i_user_peri39._GEN[76] ),
    .B(net2191));
 sg13g2_a22oi_1 _13803_ (.Y(_05653_),
    .B1(net2169),
    .B2(\i_peripherals.i_user_peri39._GEN[44] ),
    .A2(net2176),
    .A1(\i_peripherals.i_user_peri39._GEN[108] ));
 sg13g2_nand3_1 _13804_ (.B(_05652_),
    .C(_05653_),
    .A(_05651_),
    .Y(_05654_));
 sg13g2_a21oi_1 _13805_ (.A1(_01058_),
    .A2(net2090),
    .Y(_05655_),
    .B1(net2196));
 sg13g2_a221oi_1 _13806_ (.B2(_05655_),
    .C1(net1984),
    .B1(_05654_),
    .A1(net3784),
    .Y(_05656_),
    .A2(net2086));
 sg13g2_o21ai_1 _13807_ (.B1(net2279),
    .Y(_05657_),
    .A1(net3870),
    .A2(_05531_));
 sg13g2_nor2_1 _13808_ (.A(_05656_),
    .B(_05657_),
    .Y(_00397_));
 sg13g2_nor2_2 _13809_ (.A(_05170_),
    .B(net1982),
    .Y(_05658_));
 sg13g2_a22oi_1 _13810_ (.Y(_05659_),
    .B1(net2163),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[13] ),
    .A2(net2177),
    .A1(net2977));
 sg13g2_a22oi_1 _13811_ (.Y(_05660_),
    .B1(net2193),
    .B2(net3020),
    .A2(net2170),
    .A1(\i_peripherals.i_user_peri39._GEN[45] ));
 sg13g2_nand2_1 _13812_ (.Y(_05661_),
    .A(\i_peripherals.i_user_peri39.instr[13] ),
    .B(net2094));
 sg13g2_nand3_1 _13813_ (.B(_05660_),
    .C(_05661_),
    .A(_05659_),
    .Y(_05662_));
 sg13g2_a22oi_1 _13814_ (.Y(_05663_),
    .B1(net1956),
    .B2(_05662_),
    .A2(net1981),
    .A1(net3243));
 sg13g2_nor2_1 _13815_ (.A(net2250),
    .B(net3244),
    .Y(_00398_));
 sg13g2_a22oi_1 _13816_ (.Y(_05664_),
    .B1(net2160),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[14] ),
    .A2(net2177),
    .A1(\i_peripherals.i_user_peri39._GEN[110] ));
 sg13g2_inv_1 _13817_ (.Y(_05665_),
    .A(_05664_));
 sg13g2_a221oi_1 _13818_ (.B2(\i_peripherals.i_user_peri39._GEN[78] ),
    .C1(_05665_),
    .B1(net2193),
    .A1(\i_peripherals.i_user_peri39._GEN[46] ),
    .Y(_05666_),
    .A2(net2170));
 sg13g2_nor2_1 _13819_ (.A(\i_peripherals.i_user_peri39.instr[14] ),
    .B(net2089),
    .Y(_05667_));
 sg13g2_a21oi_1 _13820_ (.A1(net2087),
    .A2(_05666_),
    .Y(_05668_),
    .B1(_05667_));
 sg13g2_a22oi_1 _13821_ (.Y(_05669_),
    .B1(net1957),
    .B2(_05668_),
    .A2(net1983),
    .A1(net3260));
 sg13g2_nor2_1 _13822_ (.A(net2250),
    .B(net3261),
    .Y(_00399_));
 sg13g2_a22oi_1 _13823_ (.Y(_05670_),
    .B1(net2160),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[15] ),
    .A2(net2175),
    .A1(net3108));
 sg13g2_a22oi_1 _13824_ (.Y(_05671_),
    .B1(net2189),
    .B2(net2878),
    .A2(net2168),
    .A1(net3066));
 sg13g2_nand2_1 _13825_ (.Y(_05672_),
    .A(\i_peripherals.i_user_peri39.instr[15] ),
    .B(net2092));
 sg13g2_nand3_1 _13826_ (.B(_05671_),
    .C(_05672_),
    .A(_05670_),
    .Y(_05673_));
 sg13g2_a22oi_1 _13827_ (.Y(_05674_),
    .B1(net1956),
    .B2(_05673_),
    .A2(net1983),
    .A1(net3204));
 sg13g2_nor2_1 _13828_ (.A(net2250),
    .B(net3205),
    .Y(_00400_));
 sg13g2_a22oi_1 _13829_ (.Y(_05675_),
    .B1(net2170),
    .B2(net2822),
    .A2(net2177),
    .A1(net2926));
 sg13g2_nand2_1 _13830_ (.Y(_05676_),
    .A(net2902),
    .B(net2193));
 sg13g2_a22oi_1 _13831_ (.Y(_05677_),
    .B1(net2160),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[16] ),
    .A2(net2094),
    .A1(\i_peripherals.i_user_peri39.instr[16] ));
 sg13g2_nand3_1 _13832_ (.B(_05676_),
    .C(_05677_),
    .A(_05675_),
    .Y(_05678_));
 sg13g2_a22oi_1 _13833_ (.Y(_05679_),
    .B1(net1956),
    .B2(_05678_),
    .A2(net1981),
    .A1(net3313));
 sg13g2_nor2_1 _13834_ (.A(net2252),
    .B(net3314),
    .Y(_00401_));
 sg13g2_a22oi_1 _13835_ (.Y(_05680_),
    .B1(net2172),
    .B2(net2865),
    .A2(net2175),
    .A1(net3085));
 sg13g2_nand2_1 _13836_ (.Y(_05681_),
    .A(net2847),
    .B(net2189));
 sg13g2_a22oi_1 _13837_ (.Y(_05682_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[17] ),
    .A2(net2092),
    .A1(\i_peripherals.i_user_peri39.instr[17] ));
 sg13g2_nand3_1 _13838_ (.B(_05681_),
    .C(_05682_),
    .A(_05680_),
    .Y(_05683_));
 sg13g2_a22oi_1 _13839_ (.Y(_05684_),
    .B1(net1956),
    .B2(_05683_),
    .A2(net1981),
    .A1(net3226));
 sg13g2_nor2_1 _13840_ (.A(net2250),
    .B(net3227),
    .Y(_00402_));
 sg13g2_nand2_1 _13841_ (.Y(_05685_),
    .A(net2953),
    .B(net2193));
 sg13g2_a22oi_1 _13842_ (.Y(_05686_),
    .B1(net2168),
    .B2(net2960),
    .A2(net2175),
    .A1(net2872));
 sg13g2_a22oi_1 _13843_ (.Y(_05687_),
    .B1(net2160),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[18] ),
    .A2(net2092),
    .A1(\i_peripherals.i_user_peri39.instr[18] ));
 sg13g2_nand3_1 _13844_ (.B(_05686_),
    .C(_05687_),
    .A(_05685_),
    .Y(_05688_));
 sg13g2_a22oi_1 _13845_ (.Y(_05689_),
    .B1(net1957),
    .B2(_05688_),
    .A2(net1981),
    .A1(net3284));
 sg13g2_nor2_1 _13846_ (.A(net2252),
    .B(net3285),
    .Y(_00403_));
 sg13g2_nand2_1 _13847_ (.Y(_05690_),
    .A(net2981),
    .B(net2168));
 sg13g2_a22oi_1 _13848_ (.Y(_05691_),
    .B1(net2189),
    .B2(net2880),
    .A2(net2175),
    .A1(net3001));
 sg13g2_a22oi_1 _13849_ (.Y(_05692_),
    .B1(net2160),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[19] ),
    .A2(net2092),
    .A1(\i_peripherals.i_user_peri39.instr[19] ));
 sg13g2_nand3_1 _13850_ (.B(_05691_),
    .C(_05692_),
    .A(_05690_),
    .Y(_05693_));
 sg13g2_a22oi_1 _13851_ (.Y(_05694_),
    .B1(net1956),
    .B2(_05693_),
    .A2(net1981),
    .A1(net3301));
 sg13g2_nor2_1 _13852_ (.A(net2250),
    .B(net3302),
    .Y(_00404_));
 sg13g2_a22oi_1 _13853_ (.Y(_05695_),
    .B1(net2172),
    .B2(\i_peripherals.i_user_peri39._GEN[52] ),
    .A2(net2179),
    .A1(\i_peripherals.i_user_peri39._GEN[116] ));
 sg13g2_nand2_1 _13854_ (.Y(_05696_),
    .A(\i_peripherals.i_user_peri39._GEN[84] ),
    .B(net2189));
 sg13g2_a22oi_1 _13855_ (.Y(_05697_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[20] ),
    .A2(net2091),
    .A1(\i_peripherals.i_user_peri39.instr[20] ));
 sg13g2_nand3_1 _13856_ (.B(_05696_),
    .C(_05697_),
    .A(_05695_),
    .Y(_05698_));
 sg13g2_a22oi_1 _13857_ (.Y(_05699_),
    .B1(_05658_),
    .B2(_05698_),
    .A2(net1981),
    .A1(net3286));
 sg13g2_nor2_1 _13858_ (.A(net2252),
    .B(net3287),
    .Y(_00405_));
 sg13g2_a22oi_1 _13859_ (.Y(_05700_),
    .B1(net2189),
    .B2(net2841),
    .A2(net2179),
    .A1(net2951));
 sg13g2_nand2_1 _13860_ (.Y(_05701_),
    .A(net2911),
    .B(net2172));
 sg13g2_a22oi_1 _13861_ (.Y(_05702_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[21] ),
    .A2(net2091),
    .A1(\i_peripherals.i_user_peri39.instr[21] ));
 sg13g2_nand3_1 _13862_ (.B(_05701_),
    .C(_05702_),
    .A(_05700_),
    .Y(_05703_));
 sg13g2_a22oi_1 _13863_ (.Y(_05704_),
    .B1(net1956),
    .B2(_05703_),
    .A2(net1981),
    .A1(net3221));
 sg13g2_nor2_1 _13864_ (.A(net2252),
    .B(net3222),
    .Y(_00406_));
 sg13g2_a22oi_1 _13865_ (.Y(_05705_),
    .B1(net2189),
    .B2(net2913),
    .A2(net2179),
    .A1(net3150));
 sg13g2_nand2_1 _13866_ (.Y(_05706_),
    .A(net2983),
    .B(net2172));
 sg13g2_a22oi_1 _13867_ (.Y(_05707_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[22] ),
    .A2(net2091),
    .A1(\i_peripherals.i_user_peri39.instr[22] ));
 sg13g2_nand3_1 _13868_ (.B(_05706_),
    .C(_05707_),
    .A(_05705_),
    .Y(_05708_));
 sg13g2_a22oi_1 _13869_ (.Y(_05709_),
    .B1(net1957),
    .B2(_05708_),
    .A2(net1982),
    .A1(net3258));
 sg13g2_nor2_1 _13870_ (.A(net2252),
    .B(net3259),
    .Y(_00407_));
 sg13g2_nand2_1 _13871_ (.Y(_05710_),
    .A(net3049),
    .B(net2190));
 sg13g2_a22oi_1 _13872_ (.Y(_05711_),
    .B1(net2171),
    .B2(net3013),
    .A2(net2178),
    .A1(net3011));
 sg13g2_a22oi_1 _13873_ (.Y(_05712_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[23] ),
    .A2(net2091),
    .A1(\i_peripherals.i_user_peri39.instr[23] ));
 sg13g2_nand3_1 _13874_ (.B(_05711_),
    .C(_05712_),
    .A(_05710_),
    .Y(_05713_));
 sg13g2_a22oi_1 _13875_ (.Y(_05714_),
    .B1(net1957),
    .B2(_05713_),
    .A2(net1982),
    .A1(net3315));
 sg13g2_nor2_1 _13876_ (.A(net2251),
    .B(net3316),
    .Y(_00408_));
 sg13g2_a22oi_1 _13877_ (.Y(_05715_),
    .B1(net2162),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[24] ),
    .A2(net2178),
    .A1(\i_peripherals.i_user_peri39._GEN[120] ));
 sg13g2_inv_1 _13878_ (.Y(_05716_),
    .A(_05715_));
 sg13g2_a221oi_1 _13879_ (.B2(\i_peripherals.i_user_peri39._GEN[88] ),
    .C1(_05716_),
    .B1(net2191),
    .A1(\i_peripherals.i_user_peri39._GEN[56] ),
    .Y(_05717_),
    .A2(net2171));
 sg13g2_nor2_1 _13880_ (.A(\i_peripherals.i_user_peri39.instr[24] ),
    .B(net2087),
    .Y(_05718_));
 sg13g2_a21oi_1 _13881_ (.A1(net2087),
    .A2(_05717_),
    .Y(_05719_),
    .B1(_05718_));
 sg13g2_a22oi_1 _13882_ (.Y(_05720_),
    .B1(net1957),
    .B2(_05719_),
    .A2(net1982),
    .A1(net3368));
 sg13g2_nor2_1 _13883_ (.A(net2250),
    .B(net3369),
    .Y(_00409_));
 sg13g2_a22oi_1 _13884_ (.Y(_05721_),
    .B1(net2168),
    .B2(net2817),
    .A2(net2175),
    .A1(net3206));
 sg13g2_nand2_1 _13885_ (.Y(_05722_),
    .A(net2807),
    .B(net2190));
 sg13g2_a22oi_1 _13886_ (.Y(_05723_),
    .B1(net2160),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[25] ),
    .A2(net2092),
    .A1(\i_peripherals.i_user_peri39.instr[25] ));
 sg13g2_nand3_1 _13887_ (.B(_05722_),
    .C(_05723_),
    .A(_05721_),
    .Y(_05724_));
 sg13g2_a22oi_1 _13888_ (.Y(_05725_),
    .B1(net1956),
    .B2(_05724_),
    .A2(net1981),
    .A1(net3256));
 sg13g2_nor2_1 _13889_ (.A(net2250),
    .B(net3257),
    .Y(_00410_));
 sg13g2_nand2_1 _13890_ (.Y(_05726_),
    .A(net2972),
    .B(net2172));
 sg13g2_a22oi_1 _13891_ (.Y(_05727_),
    .B1(net2189),
    .B2(net2826),
    .A2(net2179),
    .A1(net2886));
 sg13g2_a22oi_1 _13892_ (.Y(_05728_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[26] ),
    .A2(net2091),
    .A1(\i_peripherals.i_user_peri39.instr[26] ));
 sg13g2_nand3_1 _13893_ (.B(_05727_),
    .C(_05728_),
    .A(_05726_),
    .Y(_05729_));
 sg13g2_a22oi_1 _13894_ (.Y(_05730_),
    .B1(_05658_),
    .B2(_05729_),
    .A2(net1983),
    .A1(net3269));
 sg13g2_nor2_1 _13895_ (.A(net2251),
    .B(net3270),
    .Y(_00411_));
 sg13g2_a22oi_1 _13896_ (.Y(_05731_),
    .B1(net2163),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[27] ),
    .A2(net2177),
    .A1(\i_peripherals.i_user_peri39._GEN[123] ));
 sg13g2_inv_1 _13897_ (.Y(_05732_),
    .A(_05731_));
 sg13g2_a221oi_1 _13898_ (.B2(\i_peripherals.i_user_peri39._GEN[91] ),
    .C1(_05732_),
    .B1(net2193),
    .A1(\i_peripherals.i_user_peri39._GEN[59] ),
    .Y(_05733_),
    .A2(net2170));
 sg13g2_nor2_1 _13899_ (.A(\i_peripherals.i_user_peri39.instr[27] ),
    .B(net2087),
    .Y(_05734_));
 sg13g2_a21oi_1 _13900_ (.A1(net2087),
    .A2(_05733_),
    .Y(_05735_),
    .B1(_05734_));
 sg13g2_a22oi_1 _13901_ (.Y(_05736_),
    .B1(net1957),
    .B2(_05735_),
    .A2(net1982),
    .A1(net3282));
 sg13g2_nor2_1 _13902_ (.A(net2251),
    .B(net3283),
    .Y(_00412_));
 sg13g2_a22oi_1 _13903_ (.Y(_05737_),
    .B1(net2168),
    .B2(net2955),
    .A2(net2175),
    .A1(net2979));
 sg13g2_nand2_1 _13904_ (.Y(_05738_),
    .A(net2874),
    .B(net2190));
 sg13g2_a22oi_1 _13905_ (.Y(_05739_),
    .B1(net2164),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[28] ),
    .A2(net2092),
    .A1(\i_peripherals.i_user_peri39.instr[28] ));
 sg13g2_nand3_1 _13906_ (.B(_05738_),
    .C(_05739_),
    .A(_05737_),
    .Y(_05740_));
 sg13g2_a22oi_1 _13907_ (.Y(_05741_),
    .B1(_05658_),
    .B2(_05740_),
    .A2(net1983),
    .A1(net3323));
 sg13g2_nor2_1 _13908_ (.A(net2251),
    .B(net3324),
    .Y(_00413_));
 sg13g2_nand2_1 _13909_ (.Y(_05742_),
    .A(\i_peripherals.i_user_peri39._GEN[93] ),
    .B(net2193));
 sg13g2_a22oi_1 _13910_ (.Y(_05743_),
    .B1(net2170),
    .B2(\i_peripherals.i_user_peri39._GEN[61] ),
    .A2(net2177),
    .A1(\i_peripherals.i_user_peri39._GEN[125] ));
 sg13g2_a21oi_1 _13911_ (.A1(\i_peripherals.i_user_peri39.math_result_reg[29] ),
    .A2(net2160),
    .Y(_05744_),
    .B1(net2094));
 sg13g2_nand3_1 _13912_ (.B(_05743_),
    .C(_05744_),
    .A(_05742_),
    .Y(_05745_));
 sg13g2_o21ai_1 _13913_ (.B1(_05745_),
    .Y(_05746_),
    .A1(net3372),
    .A2(net2089));
 sg13g2_o21ai_1 _13914_ (.B1(_05531_),
    .Y(_05747_),
    .A1(_05170_),
    .A2(_05746_));
 sg13g2_o21ai_1 _13915_ (.B1(net2278),
    .Y(_05748_),
    .A1(net3619),
    .A2(_05531_));
 sg13g2_nor2b_1 _13916_ (.A(_05748_),
    .B_N(_05747_),
    .Y(_00414_));
 sg13g2_a22oi_1 _13917_ (.Y(_05749_),
    .B1(net2170),
    .B2(net2853),
    .A2(net2177),
    .A1(net2918));
 sg13g2_nand2_1 _13918_ (.Y(_05750_),
    .A(net3134),
    .B(net2193));
 sg13g2_a22oi_1 _13919_ (.Y(_05751_),
    .B1(net2163),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[30] ),
    .A2(net2094),
    .A1(\i_peripherals.i_user_peri39.instr[30] ));
 sg13g2_nand3_1 _13920_ (.B(_05750_),
    .C(_05751_),
    .A(_05749_),
    .Y(_05752_));
 sg13g2_a22oi_1 _13921_ (.Y(_05753_),
    .B1(net1956),
    .B2(_05752_),
    .A2(net1982),
    .A1(net3305));
 sg13g2_nor2_1 _13922_ (.A(net2250),
    .B(net3306),
    .Y(_00415_));
 sg13g2_a22oi_1 _13923_ (.Y(_05754_),
    .B1(net2193),
    .B2(net3005),
    .A2(net2175),
    .A1(net3051));
 sg13g2_nand2_1 _13924_ (.Y(_05755_),
    .A(net2898),
    .B(net2168));
 sg13g2_a22oi_1 _13925_ (.Y(_05756_),
    .B1(net2160),
    .B2(\i_peripherals.i_user_peri39.math_result_reg[31] ),
    .A2(net2092),
    .A1(\i_peripherals.i_user_peri39.instr[31] ));
 sg13g2_nand3_1 _13926_ (.B(_05755_),
    .C(_05756_),
    .A(_05754_),
    .Y(_05757_));
 sg13g2_a22oi_1 _13927_ (.Y(_05758_),
    .B1(net1957),
    .B2(_05757_),
    .A2(net1982),
    .A1(net3234));
 sg13g2_nor2_1 _13928_ (.A(net2251),
    .B(net3235),
    .Y(_00416_));
 sg13g2_nand3_1 _13929_ (.B(_01433_),
    .C(net2300),
    .A(\i_tinyqv.cpu.is_load ),
    .Y(_05759_));
 sg13g2_a21oi_1 _13930_ (.A1(net3331),
    .A2(_05759_),
    .Y(_05760_),
    .B1(net1986));
 sg13g2_nor2_1 _13931_ (.A(net2248),
    .B(net3332),
    .Y(_00417_));
 sg13g2_nand2_1 _13932_ (.Y(_05761_),
    .A(net3694),
    .B(_02064_));
 sg13g2_o21ai_1 _13933_ (.B1(net3365),
    .Y(_05762_),
    .A1(\i_debug_uart_tx.fsm_state[2] ),
    .A2(net3182));
 sg13g2_nand4_1 _13934_ (.B(_02066_),
    .C(net3695),
    .A(net2256),
    .Y(_00418_),
    .D(_05762_));
 sg13g2_nand3_1 _13935_ (.B(net3203),
    .C(\i_debug_uart_tx.cycle_counter[0] ),
    .A(net3354),
    .Y(_05763_));
 sg13g2_nor3_2 _13936_ (.A(net2744),
    .B(_01024_),
    .C(_05763_),
    .Y(_05764_));
 sg13g2_and3_2 _13937_ (.X(_05765_),
    .A(_02064_),
    .B(_05762_),
    .C(_05764_));
 sg13g2_nand3_1 _13938_ (.B(_05762_),
    .C(_05764_),
    .A(_02064_),
    .Y(_05766_));
 sg13g2_and2_1 _13939_ (.A(\i_debug_uart_tx.data_to_send[0] ),
    .B(_05766_),
    .X(_05767_));
 sg13g2_a21oi_1 _13940_ (.A1(net3294),
    .A2(_05765_),
    .Y(_05768_),
    .B1(_05767_));
 sg13g2_a21oi_1 _13941_ (.A1(_01926_),
    .A2(_01932_),
    .Y(_05769_),
    .B1(_02430_));
 sg13g2_and3_1 _13942_ (.X(_05770_),
    .A(\addr[4] ),
    .B(_01935_),
    .C(_02065_));
 sg13g2_nand4_1 _13943_ (.B(_01932_),
    .C(_05769_),
    .A(\addr[3] ),
    .Y(_05771_),
    .D(_05770_));
 sg13g2_inv_2 _13944_ (.Y(_05772_),
    .A(net1978));
 sg13g2_o21ai_1 _13945_ (.B1(net2255),
    .Y(_05773_),
    .A1(net2399),
    .A2(net1979));
 sg13g2_a21oi_1 _13946_ (.A1(net3295),
    .A2(net1979),
    .Y(_00419_),
    .B1(_05773_));
 sg13g2_and2_1 _13947_ (.A(net3294),
    .B(_05766_),
    .X(_05774_));
 sg13g2_a21oi_1 _13948_ (.A1(net3545),
    .A2(_05765_),
    .Y(_05775_),
    .B1(_05774_));
 sg13g2_o21ai_1 _13949_ (.B1(net2255),
    .Y(_05776_),
    .A1(net2397),
    .A2(net1978));
 sg13g2_a21oi_1 _13950_ (.A1(net1978),
    .A2(_05775_),
    .Y(_00420_),
    .B1(_05776_));
 sg13g2_and2_1 _13951_ (.A(\i_debug_uart_tx.data_to_send[2] ),
    .B(_05766_),
    .X(_05777_));
 sg13g2_a21oi_1 _13952_ (.A1(net3472),
    .A2(_05765_),
    .Y(_05778_),
    .B1(_05777_));
 sg13g2_o21ai_1 _13953_ (.B1(net2255),
    .Y(_05779_),
    .A1(net2395),
    .A2(net1978));
 sg13g2_a21oi_1 _13954_ (.A1(net1978),
    .A2(net3473),
    .Y(_00421_),
    .B1(_05779_));
 sg13g2_and2_1 _13955_ (.A(net3472),
    .B(_05766_),
    .X(_05780_));
 sg13g2_a21oi_1 _13956_ (.A1(net3671),
    .A2(_05765_),
    .Y(_05781_),
    .B1(_05780_));
 sg13g2_o21ai_1 _13957_ (.B1(net2255),
    .Y(_05782_),
    .A1(net2393),
    .A2(net1978));
 sg13g2_a21oi_1 _13958_ (.A1(net1978),
    .A2(_05781_),
    .Y(_00422_),
    .B1(_05782_));
 sg13g2_and2_1 _13959_ (.A(net3671),
    .B(_05766_),
    .X(_05783_));
 sg13g2_a21oi_1 _13960_ (.A1(net3796),
    .A2(_05765_),
    .Y(_05784_),
    .B1(_05783_));
 sg13g2_o21ai_1 _13961_ (.B1(net2255),
    .Y(_05785_),
    .A1(net2391),
    .A2(net1979));
 sg13g2_a21oi_1 _13962_ (.A1(net1979),
    .A2(_05784_),
    .Y(_00423_),
    .B1(_05785_));
 sg13g2_mux2_1 _13963_ (.A0(net4141),
    .A1(net3796),
    .S(_05766_),
    .X(_05786_));
 sg13g2_o21ai_1 _13964_ (.B1(net2255),
    .Y(_05787_),
    .A1(_05772_),
    .A2(_05786_));
 sg13g2_a21oi_1 _13965_ (.A1(net2352),
    .A2(_05772_),
    .Y(_00424_),
    .B1(_05787_));
 sg13g2_mux2_1 _13966_ (.A0(net2794),
    .A1(\i_debug_uart_tx.data_to_send[6] ),
    .S(_05766_),
    .X(_05788_));
 sg13g2_o21ai_1 _13967_ (.B1(net2256),
    .Y(_05789_),
    .A1(_05772_),
    .A2(_05788_));
 sg13g2_a21oi_1 _13968_ (.A1(_00968_),
    .A2(_05772_),
    .Y(_00425_),
    .B1(_05789_));
 sg13g2_nand2_1 _13969_ (.Y(_05790_),
    .A(net2794),
    .B(_05766_));
 sg13g2_o21ai_1 _13970_ (.B1(net2255),
    .Y(_05791_),
    .A1(\data_to_write[7] ),
    .A2(net1978));
 sg13g2_a21oi_1 _13971_ (.A1(net1979),
    .A2(_05790_),
    .Y(_00426_),
    .B1(_05791_));
 sg13g2_and2_1 _13972_ (.A(net3201),
    .B(_02066_),
    .X(_05792_));
 sg13g2_nand2b_2 _13973_ (.Y(_05793_),
    .B(net2257),
    .A_N(_05764_));
 sg13g2_nor2_1 _13974_ (.A(net3201),
    .B(_02066_),
    .Y(_05794_));
 sg13g2_nor3_1 _13975_ (.A(_05792_),
    .B(_05793_),
    .C(net3202),
    .Y(_00427_));
 sg13g2_nor2_1 _13976_ (.A(net3203),
    .B(_05792_),
    .Y(_05795_));
 sg13g2_and2_1 _13977_ (.A(net3203),
    .B(_05792_),
    .X(_05796_));
 sg13g2_nor3_1 _13978_ (.A(_05793_),
    .B(_05795_),
    .C(_05796_),
    .Y(_00428_));
 sg13g2_nor2_1 _13979_ (.A(net3354),
    .B(_05796_),
    .Y(_05797_));
 sg13g2_and2_1 _13980_ (.A(net3354),
    .B(_05796_),
    .X(_05798_));
 sg13g2_nor3_1 _13981_ (.A(_05793_),
    .B(_05797_),
    .C(_05798_),
    .Y(_00429_));
 sg13g2_xnor2_1 _13982_ (.Y(_05799_),
    .A(net3553),
    .B(_05798_));
 sg13g2_nor2_1 _13983_ (.A(_05793_),
    .B(_05799_),
    .Y(_00430_));
 sg13g2_nand2_1 _13984_ (.Y(_05800_),
    .A(net2744),
    .B(net2257));
 sg13g2_a21oi_1 _13985_ (.A1(\i_debug_uart_tx.cycle_counter[3] ),
    .A2(_05798_),
    .Y(_00431_),
    .B1(_05800_));
 sg13g2_nor2b_1 _13986_ (.A(\i_debug_uart_tx.fsm_state[2] ),
    .B_N(\i_debug_uart_tx.fsm_state[3] ),
    .Y(_05801_));
 sg13g2_a21oi_1 _13987_ (.A1(net3182),
    .A2(_05801_),
    .Y(_05802_),
    .B1(net3988));
 sg13g2_a21oi_1 _13988_ (.A1(_02064_),
    .A2(_05802_),
    .Y(_05803_),
    .B1(_05772_));
 sg13g2_nor2_1 _13989_ (.A(_02065_),
    .B(_05764_),
    .Y(_05804_));
 sg13g2_or3_1 _13990_ (.A(net2247),
    .B(_05803_),
    .C(_05804_),
    .X(_05805_));
 sg13g2_o21ai_1 _13991_ (.B1(_05805_),
    .Y(_00432_),
    .A1(_01023_),
    .A2(_05793_));
 sg13g2_nor3_1 _13992_ (.A(_01022_),
    .B(_05802_),
    .C(_05804_),
    .Y(_05806_));
 sg13g2_a21oi_1 _13993_ (.A1(\i_debug_uart_tx.fsm_state[0] ),
    .A2(_05764_),
    .Y(_05807_),
    .B1(net3182));
 sg13g2_nor3_1 _13994_ (.A(net2247),
    .B(_05806_),
    .C(net3183),
    .Y(_00433_));
 sg13g2_and3_1 _13995_ (.X(_05808_),
    .A(net3182),
    .B(\i_debug_uart_tx.fsm_state[0] ),
    .C(_05764_));
 sg13g2_nand2_1 _13996_ (.Y(_05809_),
    .A(net3956),
    .B(_05808_));
 sg13g2_o21ai_1 _13997_ (.B1(net2255),
    .Y(_05810_),
    .A1(net3956),
    .A2(_05808_));
 sg13g2_nor2b_1 _13998_ (.A(net3957),
    .B_N(_05809_),
    .Y(_00434_));
 sg13g2_nor2b_1 _13999_ (.A(net3365),
    .B_N(_05809_),
    .Y(_05811_));
 sg13g2_xnor2_1 _14000_ (.Y(_05812_),
    .A(\i_debug_uart_tx.fsm_state[2] ),
    .B(\i_debug_uart_tx.fsm_state[0] ));
 sg13g2_and4_1 _14001_ (.A(net3365),
    .B(net3182),
    .C(_05764_),
    .D(_05812_),
    .X(_05813_));
 sg13g2_nor3_1 _14002_ (.A(net2247),
    .B(net3366),
    .C(_05813_),
    .Y(_00435_));
 sg13g2_nor2_2 _14003_ (.A(_01990_),
    .B(_02018_),
    .Y(_05814_));
 sg13g2_and2_1 _14004_ (.A(net2245),
    .B(_05814_),
    .X(_05815_));
 sg13g2_nand2_2 _14005_ (.Y(_05816_),
    .A(net2245),
    .B(_05814_));
 sg13g2_nor2_1 _14006_ (.A(_02732_),
    .B(_05816_),
    .Y(_05817_));
 sg13g2_o21ai_1 _14007_ (.B1(net1994),
    .Y(_05818_),
    .A1(net3471),
    .A2(_05817_));
 sg13g2_nor2b_2 _14008_ (.A(_02737_),
    .B_N(net2374),
    .Y(_05819_));
 sg13g2_a21oi_1 _14009_ (.A1(_05817_),
    .A2(_05819_),
    .Y(_00436_),
    .B1(_05818_));
 sg13g2_nor3_2 _14010_ (.A(_01261_),
    .B(_01268_),
    .C(_02706_),
    .Y(_05820_));
 sg13g2_o21ai_1 _14011_ (.B1(net2855),
    .Y(_05821_),
    .A1(_05816_),
    .A2(_05820_));
 sg13g2_o21ai_1 _14012_ (.B1(net2373),
    .Y(_05822_),
    .A1(net2371),
    .A2(_01419_));
 sg13g2_nor2b_2 _14013_ (.A(_01269_),
    .B_N(_05822_),
    .Y(_05823_));
 sg13g2_nand2_1 _14014_ (.Y(_05824_),
    .A(_05815_),
    .B(_05823_));
 sg13g2_a21oi_1 _14015_ (.A1(_05821_),
    .A2(_05824_),
    .Y(_00437_),
    .B1(net1993));
 sg13g2_nor2_2 _14016_ (.A(_01305_),
    .B(_02706_),
    .Y(_05825_));
 sg13g2_o21ai_1 _14017_ (.B1(net2894),
    .Y(_05826_),
    .A1(_05816_),
    .A2(_05825_));
 sg13g2_and2_1 _14018_ (.A(_01305_),
    .B(_05822_),
    .X(_05827_));
 sg13g2_nand2_1 _14019_ (.Y(_05828_),
    .A(_05815_),
    .B(_05827_));
 sg13g2_a21oi_1 _14020_ (.A1(_05826_),
    .A2(_05828_),
    .Y(_00438_),
    .B1(net1993));
 sg13g2_nor2_2 _14021_ (.A(_01341_),
    .B(_02706_),
    .Y(_05829_));
 sg13g2_o21ai_1 _14022_ (.B1(net3236),
    .Y(_05830_),
    .A1(_05816_),
    .A2(_05829_));
 sg13g2_and2_1 _14023_ (.A(_01341_),
    .B(_05822_),
    .X(_05831_));
 sg13g2_nand2_1 _14024_ (.Y(_05832_),
    .A(_05815_),
    .B(_05831_));
 sg13g2_a21oi_1 _14025_ (.A1(_05830_),
    .A2(_05832_),
    .Y(_00439_),
    .B1(net1993));
 sg13g2_nand2_2 _14026_ (.Y(_05833_),
    .A(net2244),
    .B(_05814_));
 sg13g2_nor2_1 _14027_ (.A(_02732_),
    .B(_05833_),
    .Y(_05834_));
 sg13g2_o21ai_1 _14028_ (.B1(net1994),
    .Y(_05835_),
    .A1(net3460),
    .A2(_05834_));
 sg13g2_a21oi_1 _14029_ (.A1(_05819_),
    .A2(_05834_),
    .Y(_00440_),
    .B1(_05835_));
 sg13g2_nor2_1 _14030_ (.A(_05820_),
    .B(_05833_),
    .Y(_05836_));
 sg13g2_o21ai_1 _14031_ (.B1(net1994),
    .Y(_05837_),
    .A1(net3809),
    .A2(_05836_));
 sg13g2_nor3_1 _14032_ (.A(_05820_),
    .B(_05823_),
    .C(_05833_),
    .Y(_05838_));
 sg13g2_nor2_1 _14033_ (.A(_05837_),
    .B(_05838_),
    .Y(_00441_));
 sg13g2_nor2_1 _14034_ (.A(_05825_),
    .B(_05833_),
    .Y(_05839_));
 sg13g2_o21ai_1 _14035_ (.B1(net1994),
    .Y(_05840_),
    .A1(net3710),
    .A2(_05839_));
 sg13g2_nor3_1 _14036_ (.A(_05825_),
    .B(_05827_),
    .C(_05833_),
    .Y(_05841_));
 sg13g2_nor2_1 _14037_ (.A(_05840_),
    .B(_05841_),
    .Y(_00442_));
 sg13g2_o21ai_1 _14038_ (.B1(net3110),
    .Y(_05842_),
    .A1(_05829_),
    .A2(_05833_));
 sg13g2_nand3_1 _14039_ (.B(_05814_),
    .C(_05831_),
    .A(net2244),
    .Y(_05843_));
 sg13g2_a21oi_1 _14040_ (.A1(_05842_),
    .A2(_05843_),
    .Y(_00443_),
    .B1(net1993));
 sg13g2_nand2_2 _14041_ (.Y(_05844_),
    .A(net2242),
    .B(_05814_));
 sg13g2_nor2_1 _14042_ (.A(_02732_),
    .B(_05844_),
    .Y(_05845_));
 sg13g2_o21ai_1 _14043_ (.B1(net1995),
    .Y(_05846_),
    .A1(net3808),
    .A2(_05845_));
 sg13g2_a21oi_1 _14044_ (.A1(_05819_),
    .A2(_05845_),
    .Y(_00444_),
    .B1(_05846_));
 sg13g2_nor2_1 _14045_ (.A(_05820_),
    .B(_05844_),
    .Y(_05847_));
 sg13g2_o21ai_1 _14046_ (.B1(net1995),
    .Y(_05848_),
    .A1(net3865),
    .A2(_05847_));
 sg13g2_nor3_1 _14047_ (.A(_05820_),
    .B(_05823_),
    .C(_05844_),
    .Y(_05849_));
 sg13g2_nor2_1 _14048_ (.A(_05848_),
    .B(_05849_),
    .Y(_00445_));
 sg13g2_nor2_1 _14049_ (.A(_05825_),
    .B(_05844_),
    .Y(_05850_));
 sg13g2_o21ai_1 _14050_ (.B1(net1995),
    .Y(_05851_),
    .A1(net3908),
    .A2(_05850_));
 sg13g2_nor3_1 _14051_ (.A(_05825_),
    .B(_05827_),
    .C(_05844_),
    .Y(_05852_));
 sg13g2_nor2_1 _14052_ (.A(_05851_),
    .B(_05852_),
    .Y(_00446_));
 sg13g2_o21ai_1 _14053_ (.B1(net3310),
    .Y(_05853_),
    .A1(_05829_),
    .A2(_05844_));
 sg13g2_nand3_1 _14054_ (.B(_05814_),
    .C(_05831_),
    .A(net2242),
    .Y(_05854_));
 sg13g2_a21oi_1 _14055_ (.A1(_05853_),
    .A2(_05854_),
    .Y(_00447_),
    .B1(net1993));
 sg13g2_nor4_1 _14056_ (.A(_01344_),
    .B(_01990_),
    .C(_02018_),
    .D(_02732_),
    .Y(_05855_));
 sg13g2_o21ai_1 _14057_ (.B1(net1995),
    .Y(_05856_),
    .A1(net3920),
    .A2(_05855_));
 sg13g2_a21oi_1 _14058_ (.A1(_05819_),
    .A2(_05855_),
    .Y(_00448_),
    .B1(_05856_));
 sg13g2_nor3_1 _14059_ (.A(net2380),
    .B(net2336),
    .C(_01990_),
    .Y(_05857_));
 sg13g2_a21o_2 _14060_ (.A2(_05857_),
    .A1(_02007_),
    .B1(net2244),
    .X(_05858_));
 sg13g2_nand2_1 _14061_ (.Y(_05859_),
    .A(net2241),
    .B(_05825_));
 sg13g2_a21oi_1 _14062_ (.A1(\i_peripherals.i_uart.ui_in[1] ),
    .A2(_01138_),
    .Y(_05860_),
    .B1(net3122));
 sg13g2_nor2_1 _14063_ (.A(net2241),
    .B(_05860_),
    .Y(_05861_));
 sg13g2_a21oi_1 _14064_ (.A1(net2241),
    .A2(_05827_),
    .Y(_05862_),
    .B1(_05861_));
 sg13g2_and3_1 _14065_ (.X(_05863_),
    .A(_05858_),
    .B(_05859_),
    .C(_05862_));
 sg13g2_a21oi_1 _14066_ (.A1(_05858_),
    .A2(_05859_),
    .Y(_05864_),
    .B1(net3122));
 sg13g2_nor3_1 _14067_ (.A(net1993),
    .B(_05863_),
    .C(_05864_),
    .Y(_00449_));
 sg13g2_nand2_1 _14068_ (.Y(_05865_),
    .A(net2241),
    .B(_05829_));
 sg13g2_a21oi_1 _14069_ (.A1(_05858_),
    .A2(_05865_),
    .Y(_05866_),
    .B1(net3409));
 sg13g2_a21oi_1 _14070_ (.A1(\i_peripherals.i_uart.ui_in[0] ),
    .A2(_01137_),
    .Y(_05867_),
    .B1(net3409));
 sg13g2_nor2_1 _14071_ (.A(net2241),
    .B(_05867_),
    .Y(_05868_));
 sg13g2_a21oi_1 _14072_ (.A1(net2241),
    .A2(_05831_),
    .Y(_05869_),
    .B1(_05868_));
 sg13g2_and3_1 _14073_ (.X(_05870_),
    .A(_05858_),
    .B(_05865_),
    .C(_05869_));
 sg13g2_nor3_1 _14074_ (.A(net1993),
    .B(_05866_),
    .C(_05870_),
    .Y(_00450_));
 sg13g2_nand2_2 _14075_ (.Y(_05871_),
    .A(net2231),
    .B(_05814_));
 sg13g2_nor2_1 _14076_ (.A(_02732_),
    .B(_05871_),
    .Y(_05872_));
 sg13g2_o21ai_1 _14077_ (.B1(net1995),
    .Y(_05873_),
    .A1(net3484),
    .A2(_05872_));
 sg13g2_a21oi_1 _14078_ (.A1(_05819_),
    .A2(_05872_),
    .Y(_00451_),
    .B1(_05873_));
 sg13g2_nor2_1 _14079_ (.A(_05820_),
    .B(_05871_),
    .Y(_05874_));
 sg13g2_o21ai_1 _14080_ (.B1(net1994),
    .Y(_05875_),
    .A1(net3665),
    .A2(_05874_));
 sg13g2_nor3_1 _14081_ (.A(_05820_),
    .B(_05823_),
    .C(_05871_),
    .Y(_05876_));
 sg13g2_nor2_1 _14082_ (.A(_05875_),
    .B(_05876_),
    .Y(_00452_));
 sg13g2_nor2_1 _14083_ (.A(_05825_),
    .B(_05871_),
    .Y(_05877_));
 sg13g2_o21ai_1 _14084_ (.B1(net1994),
    .Y(_05878_),
    .A1(net3627),
    .A2(_05877_));
 sg13g2_nor3_1 _14085_ (.A(_05825_),
    .B(_05827_),
    .C(_05871_),
    .Y(_05879_));
 sg13g2_nor2_1 _14086_ (.A(_05878_),
    .B(_05879_),
    .Y(_00453_));
 sg13g2_nor2_1 _14087_ (.A(_05829_),
    .B(_05871_),
    .Y(_05880_));
 sg13g2_o21ai_1 _14088_ (.B1(net1994),
    .Y(_05881_),
    .A1(net3805),
    .A2(_05880_));
 sg13g2_nor3_1 _14089_ (.A(_05829_),
    .B(_05831_),
    .C(_05871_),
    .Y(_05882_));
 sg13g2_nor2_1 _14090_ (.A(_05881_),
    .B(_05882_),
    .Y(_00454_));
 sg13g2_o21ai_1 _14091_ (.B1(_02595_),
    .Y(_05883_),
    .A1(net2350),
    .A2(net3753));
 sg13g2_nand3b_1 _14092_ (.B(_05883_),
    .C(net2269),
    .Y(_05884_),
    .A_N(net3967));
 sg13g2_nor2_1 _14093_ (.A(_02596_),
    .B(net1731),
    .Y(_00455_));
 sg13g2_nand3_1 _14094_ (.B(_01939_),
    .C(_05769_),
    .A(_01933_),
    .Y(_05885_));
 sg13g2_nand3_1 _14095_ (.B(net3863),
    .C(_05885_),
    .A(net2267),
    .Y(_05886_));
 sg13g2_nand2_1 _14096_ (.Y(_05887_),
    .A(net2246),
    .B(net3));
 sg13g2_o21ai_1 _14097_ (.B1(_05887_),
    .Y(_05888_),
    .A1(_05168_),
    .A2(_05885_));
 sg13g2_nand2b_1 _14098_ (.Y(_00456_),
    .B(_05886_),
    .A_N(_05888_));
 sg13g2_nor3_1 _14099_ (.A(\i_tinyqv.cpu.instr_write_offset[2] ),
    .B(\i_tinyqv.cpu.instr_write_offset[1] ),
    .C(_02641_),
    .Y(_05889_));
 sg13g2_mux2_1 _14100_ (.A0(net3465),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net1741),
    .X(_00457_));
 sg13g2_mux2_1 _14101_ (.A0(net3490),
    .A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .S(net1741),
    .X(_00458_));
 sg13g2_nor2_1 _14102_ (.A(net3119),
    .B(net1739),
    .Y(_05890_));
 sg13g2_a21oi_1 _14103_ (.A1(_01118_),
    .A2(net1739),
    .Y(_00459_),
    .B1(_05890_));
 sg13g2_mux2_1 _14104_ (.A0(net3461),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(net1740),
    .X(_00460_));
 sg13g2_mux2_1 _14105_ (.A0(net3363),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net1738),
    .X(_00461_));
 sg13g2_nor2_1 _14106_ (.A(net3083),
    .B(net1738),
    .Y(_05891_));
 sg13g2_a21oi_1 _14107_ (.A1(_01134_),
    .A2(net1738),
    .Y(_00462_),
    .B1(_05891_));
 sg13g2_nand2_1 _14108_ (.Y(_05892_),
    .A(net2422),
    .B(net1738));
 sg13g2_o21ai_1 _14109_ (.B1(_05892_),
    .Y(_00463_),
    .A1(_01096_),
    .A2(net1738));
 sg13g2_nor2_1 _14110_ (.A(net3145),
    .B(net1738),
    .Y(_05893_));
 sg13g2_a21oi_1 _14111_ (.A1(_01124_),
    .A2(net1738),
    .Y(_00464_),
    .B1(_05893_));
 sg13g2_nor2_1 _14112_ (.A(net3081),
    .B(net1739),
    .Y(_05894_));
 sg13g2_a21oi_1 _14113_ (.A1(net2330),
    .A2(net1739),
    .Y(_00465_),
    .B1(_05894_));
 sg13g2_nor2_1 _14114_ (.A(net3117),
    .B(net1740),
    .Y(_05895_));
 sg13g2_a21oi_1 _14115_ (.A1(_01133_),
    .A2(net1738),
    .Y(_00466_),
    .B1(_05895_));
 sg13g2_mux2_1 _14116_ (.A0(net3597),
    .A1(net2420),
    .S(net1739),
    .X(_00467_));
 sg13g2_nor2_1 _14117_ (.A(net3147),
    .B(net1740),
    .Y(_05896_));
 sg13g2_a21oi_1 _14118_ (.A1(_01125_),
    .A2(net1740),
    .Y(_00468_),
    .B1(_05896_));
 sg13g2_nor2_1 _14119_ (.A(net3160),
    .B(net1741),
    .Y(_05897_));
 sg13g2_a21oi_1 _14120_ (.A1(_01129_),
    .A2(net1741),
    .Y(_00469_),
    .B1(net3161));
 sg13g2_mux2_1 _14121_ (.A0(net3412),
    .A1(net2419),
    .S(net1741),
    .X(_00470_));
 sg13g2_mux2_1 _14122_ (.A0(\i_tinyqv.cpu.instr_data_in[2] ),
    .A1(net3407),
    .S(net1760),
    .X(_00471_));
 sg13g2_mux2_1 _14123_ (.A0(\i_tinyqv.cpu.instr_data_in[3] ),
    .A1(net3571),
    .S(net1760),
    .X(_00472_));
 sg13g2_nand2_1 _14124_ (.Y(_05898_),
    .A(net2813),
    .B(net1759));
 sg13g2_o21ai_1 _14125_ (.B1(_05898_),
    .Y(_00473_),
    .A1(_01118_),
    .A2(net1759));
 sg13g2_mux2_1 _14126_ (.A0(\i_tinyqv.cpu.instr_data_in[5] ),
    .A1(net3653),
    .S(net1759),
    .X(_00474_));
 sg13g2_mux2_1 _14127_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(net3361),
    .S(net1758),
    .X(_00475_));
 sg13g2_nand2_1 _14128_ (.Y(_05899_),
    .A(net2830),
    .B(net1758));
 sg13g2_o21ai_1 _14129_ (.B1(_05899_),
    .Y(_00476_),
    .A1(_01134_),
    .A2(net1758));
 sg13g2_mux2_1 _14130_ (.A0(net2422),
    .A1(net3525),
    .S(net1758),
    .X(_00477_));
 sg13g2_nand2_1 _14131_ (.Y(_05900_),
    .A(net2863),
    .B(net1758));
 sg13g2_o21ai_1 _14132_ (.B1(_05900_),
    .Y(_00478_),
    .A1(_01124_),
    .A2(net1758));
 sg13g2_nand2_1 _14133_ (.Y(_05901_),
    .A(net2798),
    .B(net1759));
 sg13g2_o21ai_1 _14134_ (.B1(_05901_),
    .Y(_00479_),
    .A1(net2330),
    .A2(net1759));
 sg13g2_nand2_1 _14135_ (.Y(_05902_),
    .A(net2785),
    .B(net1758));
 sg13g2_o21ai_1 _14136_ (.B1(_05902_),
    .Y(_00480_),
    .A1(_01133_),
    .A2(net1758));
 sg13g2_mux2_1 _14137_ (.A0(net2421),
    .A1(net3391),
    .S(net1760),
    .X(_00481_));
 sg13g2_nand2_1 _14138_ (.Y(_05903_),
    .A(net2792),
    .B(net1759));
 sg13g2_o21ai_1 _14139_ (.B1(_05903_),
    .Y(_00482_),
    .A1(_01125_),
    .A2(net1759));
 sg13g2_nand2_1 _14140_ (.Y(_05904_),
    .A(net2843),
    .B(net1760));
 sg13g2_o21ai_1 _14141_ (.B1(_05904_),
    .Y(_00483_),
    .A1(_01129_),
    .A2(net1760));
 sg13g2_mux2_1 _14142_ (.A0(net2419),
    .A1(net3495),
    .S(net1760),
    .X(_00484_));
 sg13g2_nand2_2 _14143_ (.Y(_05905_),
    .A(net2237),
    .B(_02629_));
 sg13g2_mux2_1 _14144_ (.A0(_02664_),
    .A1(net2479),
    .S(_05905_),
    .X(_00485_));
 sg13g2_nand2_1 _14145_ (.Y(_05906_),
    .A(_01318_),
    .B(_01407_));
 sg13g2_nor2_1 _14146_ (.A(_01328_),
    .B(_01407_),
    .Y(_05907_));
 sg13g2_nor2_1 _14147_ (.A(_05905_),
    .B(_05907_),
    .Y(_05908_));
 sg13g2_a22oi_1 _14148_ (.Y(_00486_),
    .B1(_05906_),
    .B2(_05908_),
    .A2(_05905_),
    .A1(net2334));
 sg13g2_mux2_1 _14149_ (.A0(_01292_),
    .A1(_01282_),
    .S(_01407_),
    .X(_05909_));
 sg13g2_mux2_1 _14150_ (.A0(_05909_),
    .A1(net3862),
    .S(_05905_),
    .X(_00487_));
 sg13g2_or2_1 _14151_ (.X(_05910_),
    .B(_01407_),
    .A(_01254_));
 sg13g2_a21oi_1 _14152_ (.A1(_01223_),
    .A2(_01407_),
    .Y(_05911_),
    .B1(_05905_));
 sg13g2_a22oi_1 _14153_ (.Y(_00488_),
    .B1(_05910_),
    .B2(_05911_),
    .A2(_05905_),
    .A1(_01122_));
 sg13g2_mux2_1 _14154_ (.A0(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A1(net3579),
    .S(net2298),
    .X(_00489_));
 sg13g2_mux2_1 _14155_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(net3765),
    .S(net2297),
    .X(_00490_));
 sg13g2_mux2_1 _14156_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(net3325),
    .S(net2295),
    .X(_00491_));
 sg13g2_mux2_1 _14157_ (.A0(net3397),
    .A1(net3357),
    .S(net2298),
    .X(_00492_));
 sg13g2_mux2_1 _14158_ (.A0(net3579),
    .A1(net3581),
    .S(net2297),
    .X(_00493_));
 sg13g2_mux2_1 _14159_ (.A0(\i_tinyqv.cpu.i_core.mepc[5] ),
    .A1(net3565),
    .S(net2297),
    .X(_00494_));
 sg13g2_mux2_1 _14160_ (.A0(net3325),
    .A1(net3382),
    .S(net2295),
    .X(_00495_));
 sg13g2_mux2_1 _14161_ (.A0(net3357),
    .A1(\i_tinyqv.cpu.i_core.mepc[11] ),
    .S(net2298),
    .X(_00496_));
 sg13g2_mux2_1 _14162_ (.A0(\i_tinyqv.cpu.i_core.mepc[8] ),
    .A1(net3387),
    .S(net2297),
    .X(_00497_));
 sg13g2_mux2_1 _14163_ (.A0(\i_tinyqv.cpu.i_core.mepc[9] ),
    .A1(net3275),
    .S(net2296),
    .X(_00498_));
 sg13g2_mux2_1 _14164_ (.A0(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A1(net3344),
    .S(net2295),
    .X(_00499_));
 sg13g2_mux2_1 _14165_ (.A0(net3513),
    .A1(net3403),
    .S(net2297),
    .X(_00500_));
 sg13g2_mux2_1 _14166_ (.A0(\i_tinyqv.cpu.i_core.mepc[12] ),
    .A1(net3339),
    .S(net2297),
    .X(_00501_));
 sg13g2_mux2_1 _14167_ (.A0(net3275),
    .A1(net3355),
    .S(net2296),
    .X(_00502_));
 sg13g2_mux2_1 _14168_ (.A0(net3344),
    .A1(net3437),
    .S(net2295),
    .X(_00503_));
 sg13g2_mux2_1 _14169_ (.A0(net3403),
    .A1(net3338),
    .S(net2295),
    .X(_00504_));
 sg13g2_mux2_1 _14170_ (.A0(net3339),
    .A1(net2837),
    .S(net2296),
    .X(_00505_));
 sg13g2_mux2_1 _14171_ (.A0(net3355),
    .A1(net2861),
    .S(net2296),
    .X(_00506_));
 sg13g2_mux2_1 _14172_ (.A0(net3437),
    .A1(net2859),
    .S(net2295),
    .X(_00507_));
 sg13g2_mux2_1 _14173_ (.A0(net3338),
    .A1(net2828),
    .S(net2295),
    .X(_00508_));
 sg13g2_o21ai_1 _14174_ (.B1(_01832_),
    .Y(_05912_),
    .A1(net2368),
    .A2(_01718_));
 sg13g2_mux2_1 _14175_ (.A0(net3540),
    .A1(net2466),
    .S(net2154),
    .X(_00509_));
 sg13g2_mux2_1 _14176_ (.A0(net2463),
    .A1(net2465),
    .S(net2154),
    .X(_00510_));
 sg13g2_mux2_1 _14177_ (.A0(net2461),
    .A1(net3993),
    .S(net2154),
    .X(_00511_));
 sg13g2_mux2_1 _14178_ (.A0(net3719),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .S(_05912_),
    .X(_00512_));
 sg13g2_mux2_1 _14179_ (.A0(net2459),
    .A1(net2464),
    .S(net2154),
    .X(_00513_));
 sg13g2_mux2_1 _14180_ (.A0(net2458),
    .A1(net2463),
    .S(net2154),
    .X(_00514_));
 sg13g2_mux2_1 _14181_ (.A0(net2457),
    .A1(net2461),
    .S(net2153),
    .X(_00515_));
 sg13g2_mux2_1 _14182_ (.A0(net2456),
    .A1(net2460),
    .S(net2153),
    .X(_00516_));
 sg13g2_mux2_1 _14183_ (.A0(net2455),
    .A1(net2459),
    .S(net2153),
    .X(_00517_));
 sg13g2_mux2_1 _14184_ (.A0(net2454),
    .A1(net2458),
    .S(net2153),
    .X(_00518_));
 sg13g2_mux2_1 _14185_ (.A0(net2453),
    .A1(net3918),
    .S(net2155),
    .X(_00519_));
 sg13g2_mux2_1 _14186_ (.A0(net3638),
    .A1(net3645),
    .S(net2156),
    .X(_00520_));
 sg13g2_mux2_1 _14187_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .A1(net3538),
    .S(net2156),
    .X(_00521_));
 sg13g2_mux2_1 _14188_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .A1(net3686),
    .S(net2156),
    .X(_00522_));
 sg13g2_mux2_1 _14189_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .A1(net3615),
    .S(net2155),
    .X(_00523_));
 sg13g2_mux2_1 _14190_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .A1(net3638),
    .S(net2156),
    .X(_00524_));
 sg13g2_mux2_1 _14191_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .A1(net3721),
    .S(net2155),
    .X(_00525_));
 sg13g2_mux2_1 _14192_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .A1(net3832),
    .S(net2153),
    .X(_00526_));
 sg13g2_mux2_1 _14193_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .A1(net3848),
    .S(net2155),
    .X(_00527_));
 sg13g2_mux2_1 _14194_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .A1(net3786),
    .S(net2155),
    .X(_00528_));
 sg13g2_mux2_1 _14195_ (.A0(net3398),
    .A1(net3813),
    .S(net2155),
    .X(_00529_));
 sg13g2_mux2_1 _14196_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .A1(net3929),
    .S(net2155),
    .X(_00530_));
 sg13g2_mux2_1 _14197_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .A1(net3950),
    .S(net2156),
    .X(_00531_));
 sg13g2_mux2_1 _14198_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .A1(net3941),
    .S(net2153),
    .X(_00532_));
 sg13g2_nand2_1 _14199_ (.Y(_05913_),
    .A(net3398),
    .B(net2153));
 sg13g2_o21ai_1 _14200_ (.B1(_05913_),
    .Y(_00533_),
    .A1(_01119_),
    .A2(net2153));
 sg13g2_mux2_1 _14201_ (.A0(net3697),
    .A1(net3931),
    .S(net2156),
    .X(_00534_));
 sg13g2_mux2_1 _14202_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A1(net4018),
    .S(net2155),
    .X(_00535_));
 sg13g2_mux2_1 _14203_ (.A0(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .A1(net3980),
    .S(net2156),
    .X(_00536_));
 sg13g2_or2_1 _14204_ (.X(_05914_),
    .B(net2157),
    .A(net2145));
 sg13g2_nor2b_2 _14205_ (.A(_01896_),
    .B_N(_02629_),
    .Y(_05915_));
 sg13g2_o21ai_1 _14206_ (.B1(_02629_),
    .Y(_05916_),
    .A1(net2369),
    .A2(_01193_));
 sg13g2_nand2_2 _14207_ (.Y(_05917_),
    .A(_01195_),
    .B(_01410_));
 sg13g2_a21oi_1 _14208_ (.A1(_02225_),
    .A2(_05915_),
    .Y(_05918_),
    .B1(_05917_));
 sg13g2_o21ai_1 _14209_ (.B1(_05918_),
    .Y(_05919_),
    .A1(_01292_),
    .A2(_05915_));
 sg13g2_o21ai_1 _14210_ (.B1(_05917_),
    .Y(_05920_),
    .A1(_01261_),
    .A2(_01268_));
 sg13g2_a21oi_1 _14211_ (.A1(_05919_),
    .A2(_05920_),
    .Y(_05921_),
    .B1(_05914_));
 sg13g2_a21oi_1 _14212_ (.A1(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A2(net2157),
    .Y(_05922_),
    .B1(_05921_));
 sg13g2_o21ai_1 _14213_ (.B1(_05922_),
    .Y(_00537_),
    .A1(net2999),
    .A2(_02675_));
 sg13g2_nand2_1 _14214_ (.Y(_05923_),
    .A(_01254_),
    .B(_05916_));
 sg13g2_a21oi_1 _14215_ (.A1(_02378_),
    .A2(_05915_),
    .Y(_05924_),
    .B1(_05917_));
 sg13g2_a22oi_1 _14216_ (.Y(_05925_),
    .B1(_05923_),
    .B2(_05924_),
    .A2(_05917_),
    .A1(_01189_));
 sg13g2_nor2_1 _14217_ (.A(_02689_),
    .B(net2157),
    .Y(_05926_));
 sg13g2_a21oi_1 _14218_ (.A1(net4041),
    .A2(net2157),
    .Y(_05927_),
    .B1(_05926_));
 sg13g2_o21ai_1 _14219_ (.B1(_05927_),
    .Y(_00538_),
    .A1(_05914_),
    .A2(_05925_));
 sg13g2_nor2_1 _14220_ (.A(net2346),
    .B(net1755),
    .Y(_05928_));
 sg13g2_a22oi_1 _14221_ (.Y(_00539_),
    .B1(_05928_),
    .B2(_01087_),
    .A2(net1755),
    .A1(_01117_));
 sg13g2_a22oi_1 _14222_ (.Y(_00540_),
    .B1(_05928_),
    .B2(_01091_),
    .A2(net1755),
    .A1(_01123_));
 sg13g2_nor2_1 _14223_ (.A(_05177_),
    .B(_05512_),
    .Y(_05929_));
 sg13g2_a21oi_1 _14224_ (.A1(\data_to_write[0] ),
    .A2(net2012),
    .Y(_05930_),
    .B1(net2246));
 sg13g2_o21ai_1 _14225_ (.B1(_05930_),
    .Y(_00541_),
    .A1(_01019_),
    .A2(net2012));
 sg13g2_o21ai_1 _14226_ (.B1(net2270),
    .Y(_05931_),
    .A1(net3551),
    .A2(net2012));
 sg13g2_a21oi_1 _14227_ (.A1(_00973_),
    .A2(net2012),
    .Y(_00542_),
    .B1(_05931_));
 sg13g2_o21ai_1 _14228_ (.B1(net2271),
    .Y(_05932_),
    .A1(net3776),
    .A2(net2012));
 sg13g2_a21oi_1 _14229_ (.A1(_00972_),
    .A2(net2013),
    .Y(_00543_),
    .B1(_05932_));
 sg13g2_o21ai_1 _14230_ (.B1(net2272),
    .Y(_05933_),
    .A1(net3378),
    .A2(net2013));
 sg13g2_a21oi_1 _14231_ (.A1(_00971_),
    .A2(net2013),
    .Y(_00544_),
    .B1(_05933_));
 sg13g2_o21ai_1 _14232_ (.B1(net2271),
    .Y(_05934_),
    .A1(net3723),
    .A2(net2012));
 sg13g2_a21oi_1 _14233_ (.A1(_00970_),
    .A2(net2013),
    .Y(_00545_),
    .B1(_05934_));
 sg13g2_o21ai_1 _14234_ (.B1(net2272),
    .Y(_05935_),
    .A1(net3499),
    .A2(net2012));
 sg13g2_a21oi_1 _14235_ (.A1(net2352),
    .A2(net2012),
    .Y(_00546_),
    .B1(_05935_));
 sg13g2_nor2_2 _14236_ (.A(_05175_),
    .B(_05512_),
    .Y(_05936_));
 sg13g2_nand2_2 _14237_ (.Y(_05937_),
    .A(_05306_),
    .B(_05936_));
 sg13g2_and4_1 _14238_ (.A(net2385),
    .B(_05173_),
    .C(_05306_),
    .D(_05511_),
    .X(_05938_));
 sg13g2_a21oi_1 _14239_ (.A1(net3497),
    .A2(_05937_),
    .Y(_05939_),
    .B1(net2247));
 sg13g2_o21ai_1 _14240_ (.B1(_05939_),
    .Y(_00547_),
    .A1(net2351),
    .A2(_05937_));
 sg13g2_o21ai_1 _14241_ (.B1(net2266),
    .Y(_05940_),
    .A1(net2397),
    .A2(_05937_));
 sg13g2_a21oi_1 _14242_ (.A1(_01018_),
    .A2(_05937_),
    .Y(_00548_),
    .B1(_05940_));
 sg13g2_o21ai_1 _14243_ (.B1(net2266),
    .Y(_05941_),
    .A1(net2395),
    .A2(_05937_));
 sg13g2_a21oi_1 _14244_ (.A1(_01017_),
    .A2(_05937_),
    .Y(_00549_),
    .B1(_05941_));
 sg13g2_o21ai_1 _14245_ (.B1(net2267),
    .Y(_05942_),
    .A1(net3348),
    .A2(_05938_));
 sg13g2_a21oi_1 _14246_ (.A1(_00971_),
    .A2(_05938_),
    .Y(_00550_),
    .B1(_05942_));
 sg13g2_o21ai_1 _14247_ (.B1(net2266),
    .Y(_05943_),
    .A1(net2391),
    .A2(_05937_));
 sg13g2_a21oi_1 _14248_ (.A1(_01016_),
    .A2(_05937_),
    .Y(_00551_),
    .B1(_05943_));
 sg13g2_o21ai_1 _14249_ (.B1(net2267),
    .Y(_05944_),
    .A1(net3529),
    .A2(_05938_));
 sg13g2_a21oi_1 _14250_ (.A1(net2352),
    .A2(_05938_),
    .Y(_00552_),
    .B1(_05944_));
 sg13g2_nand2_1 _14251_ (.Y(_05945_),
    .A(_05246_),
    .B(_05936_));
 sg13g2_o21ai_1 _14252_ (.B1(net2263),
    .Y(_05946_),
    .A1(net2351),
    .A2(net1977));
 sg13g2_a21o_1 _14253_ (.A2(net1977),
    .A1(net3228),
    .B1(_05946_),
    .X(_00553_));
 sg13g2_o21ai_1 _14254_ (.B1(net2259),
    .Y(_05947_),
    .A1(net2397),
    .A2(net1976));
 sg13g2_a21oi_1 _14255_ (.A1(_01015_),
    .A2(net1976),
    .Y(_00554_),
    .B1(_05947_));
 sg13g2_o21ai_1 _14256_ (.B1(net2260),
    .Y(_05948_),
    .A1(net2395),
    .A2(net1976));
 sg13g2_a21oi_1 _14257_ (.A1(_01014_),
    .A2(net1977),
    .Y(_00555_),
    .B1(_05948_));
 sg13g2_o21ai_1 _14258_ (.B1(net2260),
    .Y(_05949_),
    .A1(net2393),
    .A2(net1976));
 sg13g2_a21oi_1 _14259_ (.A1(_01013_),
    .A2(net1976),
    .Y(_00556_),
    .B1(_05949_));
 sg13g2_o21ai_1 _14260_ (.B1(net2260),
    .Y(_05950_),
    .A1(net2391),
    .A2(net1976));
 sg13g2_a21oi_1 _14261_ (.A1(_01012_),
    .A2(net1977),
    .Y(_00557_),
    .B1(_05950_));
 sg13g2_o21ai_1 _14262_ (.B1(net2260),
    .Y(_05951_),
    .A1(net2389),
    .A2(net1976));
 sg13g2_a21oi_1 _14263_ (.A1(_01011_),
    .A2(net1976),
    .Y(_00558_),
    .B1(_05951_));
 sg13g2_nand2_2 _14264_ (.Y(_05952_),
    .A(_05216_),
    .B(_05936_));
 sg13g2_o21ai_1 _14265_ (.B1(net2262),
    .Y(_05953_),
    .A1(net2351),
    .A2(net1975));
 sg13g2_a21o_1 _14266_ (.A2(net1975),
    .A1(net3268),
    .B1(_05953_),
    .X(_00559_));
 sg13g2_o21ai_1 _14267_ (.B1(net2257),
    .Y(_05954_),
    .A1(net2397),
    .A2(net1974));
 sg13g2_a21oi_1 _14268_ (.A1(_01010_),
    .A2(net1974),
    .Y(_00560_),
    .B1(_05954_));
 sg13g2_o21ai_1 _14269_ (.B1(net2262),
    .Y(_05955_),
    .A1(net2395),
    .A2(net1974));
 sg13g2_a21oi_1 _14270_ (.A1(_01009_),
    .A2(net1975),
    .Y(_00561_),
    .B1(_05955_));
 sg13g2_o21ai_1 _14271_ (.B1(net2258),
    .Y(_05956_),
    .A1(net2393),
    .A2(net1974));
 sg13g2_a21oi_1 _14272_ (.A1(_01008_),
    .A2(net1974),
    .Y(_00562_),
    .B1(_05956_));
 sg13g2_o21ai_1 _14273_ (.B1(net2262),
    .Y(_05957_),
    .A1(net2391),
    .A2(net1974));
 sg13g2_a21oi_1 _14274_ (.A1(_01007_),
    .A2(net1975),
    .Y(_00563_),
    .B1(_05957_));
 sg13g2_o21ai_1 _14275_ (.B1(net2258),
    .Y(_05958_),
    .A1(net2389),
    .A2(net1974));
 sg13g2_a21oi_1 _14276_ (.A1(_01006_),
    .A2(net1974),
    .Y(_00564_),
    .B1(_05958_));
 sg13g2_nand4_1 _14277_ (.B(net2388),
    .C(net2158),
    .A(net2386),
    .Y(_05959_),
    .D(_05522_));
 sg13g2_o21ai_1 _14278_ (.B1(net2262),
    .Y(_05960_),
    .A1(net2351),
    .A2(net2011));
 sg13g2_a21o_1 _14279_ (.A2(net2011),
    .A1(net3215),
    .B1(_05960_),
    .X(_00565_));
 sg13g2_o21ai_1 _14280_ (.B1(net2257),
    .Y(_05961_),
    .A1(net2397),
    .A2(net2010));
 sg13g2_a21oi_1 _14281_ (.A1(_01005_),
    .A2(net2010),
    .Y(_00566_),
    .B1(_05961_));
 sg13g2_o21ai_1 _14282_ (.B1(net2262),
    .Y(_05962_),
    .A1(net2395),
    .A2(net2010));
 sg13g2_a21oi_1 _14283_ (.A1(_01004_),
    .A2(net2011),
    .Y(_00567_),
    .B1(_05962_));
 sg13g2_o21ai_1 _14284_ (.B1(net2258),
    .Y(_05963_),
    .A1(net2393),
    .A2(net2010));
 sg13g2_a21oi_1 _14285_ (.A1(_01003_),
    .A2(net2010),
    .Y(_00568_),
    .B1(_05963_));
 sg13g2_o21ai_1 _14286_ (.B1(net2262),
    .Y(_05964_),
    .A1(net2391),
    .A2(net2010));
 sg13g2_a21oi_1 _14287_ (.A1(_01002_),
    .A2(net2011),
    .Y(_00569_),
    .B1(_05964_));
 sg13g2_o21ai_1 _14288_ (.B1(net2257),
    .Y(_05965_),
    .A1(net2389),
    .A2(net2010));
 sg13g2_a21oi_1 _14289_ (.A1(_01001_),
    .A2(net2010),
    .Y(_00570_),
    .B1(_05965_));
 sg13g2_nand3_1 _14290_ (.B(net2158),
    .C(_05522_),
    .A(_05306_),
    .Y(_05966_));
 sg13g2_nand3_1 _14291_ (.B(net2158),
    .C(_05522_),
    .A(_05306_),
    .Y(_05967_));
 sg13g2_a21oi_1 _14292_ (.A1(net3617),
    .A2(_05967_),
    .Y(_05968_),
    .B1(net2247));
 sg13g2_o21ai_1 _14293_ (.B1(_05968_),
    .Y(_00571_),
    .A1(net2351),
    .A2(_05966_));
 sg13g2_o21ai_1 _14294_ (.B1(net2257),
    .Y(_05969_),
    .A1(net2397),
    .A2(net2009));
 sg13g2_a21oi_1 _14295_ (.A1(_01000_),
    .A2(net2009),
    .Y(_00572_),
    .B1(_05969_));
 sg13g2_o21ai_1 _14296_ (.B1(net2258),
    .Y(_05970_),
    .A1(net2395),
    .A2(net2009));
 sg13g2_a21oi_1 _14297_ (.A1(_00999_),
    .A2(net2009),
    .Y(_00573_),
    .B1(_05970_));
 sg13g2_o21ai_1 _14298_ (.B1(net2257),
    .Y(_05971_),
    .A1(net2393),
    .A2(net2009));
 sg13g2_a21oi_1 _14299_ (.A1(_00998_),
    .A2(net2009),
    .Y(_00574_),
    .B1(_05971_));
 sg13g2_o21ai_1 _14300_ (.B1(net2262),
    .Y(_05972_),
    .A1(net2391),
    .A2(_05967_));
 sg13g2_a21oi_1 _14301_ (.A1(_00997_),
    .A2(_05967_),
    .Y(_00575_),
    .B1(_05972_));
 sg13g2_o21ai_1 _14302_ (.B1(net2257),
    .Y(_05973_),
    .A1(net2389),
    .A2(net2009));
 sg13g2_a21oi_1 _14303_ (.A1(_00996_),
    .A2(net2009),
    .Y(_00576_),
    .B1(_05973_));
 sg13g2_nand3_1 _14304_ (.B(net2158),
    .C(_05522_),
    .A(_05246_),
    .Y(_05974_));
 sg13g2_nand3_1 _14305_ (.B(net2158),
    .C(_05522_),
    .A(_05246_),
    .Y(_05975_));
 sg13g2_o21ai_1 _14306_ (.B1(net2263),
    .Y(_05976_),
    .A1(net2399),
    .A2(net2008));
 sg13g2_a21oi_1 _14307_ (.A1(_00995_),
    .A2(net2008),
    .Y(_00577_),
    .B1(_05976_));
 sg13g2_a21oi_1 _14308_ (.A1(net3277),
    .A2(net2008),
    .Y(_05977_),
    .B1(net2247));
 sg13g2_o21ai_1 _14309_ (.B1(_05977_),
    .Y(_00578_),
    .A1(_00973_),
    .A2(_05974_));
 sg13g2_o21ai_1 _14310_ (.B1(net2263),
    .Y(_05978_),
    .A1(net2395),
    .A2(_05975_));
 sg13g2_a21oi_1 _14311_ (.A1(_00994_),
    .A2(_05975_),
    .Y(_00579_),
    .B1(_05978_));
 sg13g2_o21ai_1 _14312_ (.B1(net2263),
    .Y(_05979_),
    .A1(net2393),
    .A2(net2008));
 sg13g2_a21oi_1 _14313_ (.A1(_00993_),
    .A2(net2008),
    .Y(_00580_),
    .B1(_05979_));
 sg13g2_o21ai_1 _14314_ (.B1(net2263),
    .Y(_05980_),
    .A1(net2391),
    .A2(net2008));
 sg13g2_a21oi_1 _14315_ (.A1(_00992_),
    .A2(_05975_),
    .Y(_00581_),
    .B1(_05980_));
 sg13g2_o21ai_1 _14316_ (.B1(net2263),
    .Y(_05981_),
    .A1(net2389),
    .A2(net2008));
 sg13g2_a21oi_1 _14317_ (.A1(_00991_),
    .A2(net2008),
    .Y(_00582_),
    .B1(_05981_));
 sg13g2_nor3_2 _14318_ (.A(\i_tinyqv.cpu.data_write_n[1] ),
    .B(\i_tinyqv.cpu.data_write_n[0] ),
    .C(_01904_),
    .Y(_05982_));
 sg13g2_or2_1 _14319_ (.X(_05983_),
    .B(_05982_),
    .A(net2082));
 sg13g2_o21ai_1 _14320_ (.B1(net2279),
    .Y(_05984_),
    .A1(\data_to_write[8] ),
    .A2(net2007));
 sg13g2_a21oi_1 _14321_ (.A1(_00990_),
    .A2(net2007),
    .Y(_00583_),
    .B1(_05984_));
 sg13g2_a21oi_1 _14322_ (.A1(net3924),
    .A2(net2007),
    .Y(_05985_),
    .B1(net2252));
 sg13g2_o21ai_1 _14323_ (.B1(_05985_),
    .Y(_00584_),
    .A1(_00966_),
    .A2(net2007));
 sg13g2_o21ai_1 _14324_ (.B1(net2275),
    .Y(_05986_),
    .A1(\data_to_write[10] ),
    .A2(_05983_));
 sg13g2_a21oi_1 _14325_ (.A1(_00988_),
    .A2(net2007),
    .Y(_00585_),
    .B1(_05986_));
 sg13g2_o21ai_1 _14326_ (.B1(net2277),
    .Y(_05987_),
    .A1(\data_to_write[11] ),
    .A2(net2007));
 sg13g2_a21oi_1 _14327_ (.A1(_00987_),
    .A2(_05983_),
    .Y(_00586_),
    .B1(_05987_));
 sg13g2_o21ai_1 _14328_ (.B1(net2275),
    .Y(_05988_),
    .A1(\data_to_write[12] ),
    .A2(net2007));
 sg13g2_a21oi_1 _14329_ (.A1(_00986_),
    .A2(net2007),
    .Y(_00587_),
    .B1(_05988_));
 sg13g2_o21ai_1 _14330_ (.B1(net3937),
    .Y(_05989_),
    .A1(net3702),
    .A2(net3022));
 sg13g2_a21oi_1 _14331_ (.A1(net2039),
    .A2(_05989_),
    .Y(_00588_),
    .B1(net2253));
 sg13g2_nand3_1 _14332_ (.B(net1699),
    .C(_04921_),
    .A(_04712_),
    .Y(_05990_));
 sg13g2_and2_1 _14333_ (.A(net1945),
    .B(_04308_),
    .X(_05991_));
 sg13g2_a221oi_1 _14334_ (.B2(net1762),
    .C1(_05991_),
    .B1(_05155_),
    .A1(net1774),
    .Y(_05992_),
    .A2(_04783_));
 sg13g2_a21oi_1 _14335_ (.A1(_04716_),
    .A2(_05109_),
    .Y(_05993_),
    .B1(_05992_));
 sg13g2_and3_1 _14336_ (.X(_05994_),
    .A(_04853_),
    .B(_05990_),
    .C(_05993_));
 sg13g2_nand2_1 _14337_ (.Y(_05995_),
    .A(_05094_),
    .B(_05164_));
 sg13g2_or4_1 _14338_ (.A(_05110_),
    .B(_05126_),
    .C(_05146_),
    .D(_05995_),
    .X(_05996_));
 sg13g2_or3_1 _14339_ (.A(_05060_),
    .B(_05076_),
    .C(_05996_),
    .X(_05997_));
 sg13g2_o21ai_1 _14340_ (.B1(net1692),
    .Y(_05998_),
    .A1(_04755_),
    .A2(_05992_));
 sg13g2_a21oi_1 _14341_ (.A1(_05994_),
    .A2(_05997_),
    .Y(_05999_),
    .B1(_05998_));
 sg13g2_o21ai_1 _14342_ (.B1(_04795_),
    .Y(_06000_),
    .A1(net1692),
    .A2(_05165_));
 sg13g2_nor2_1 _14343_ (.A(_05999_),
    .B(_06000_),
    .Y(_06001_));
 sg13g2_a21oi_1 _14344_ (.A1(_01145_),
    .A2(net2198),
    .Y(_00589_),
    .B1(_06001_));
 sg13g2_nor2_1 _14345_ (.A(_05994_),
    .B(_05996_),
    .Y(_06002_));
 sg13g2_nand4_1 _14346_ (.B(_05059_),
    .C(_05075_),
    .A(_04755_),
    .Y(_06003_),
    .D(_06002_));
 sg13g2_nand3_1 _14347_ (.B(_04746_),
    .C(_06003_),
    .A(net1696),
    .Y(_06004_));
 sg13g2_a21o_1 _14348_ (.A2(_06003_),
    .A1(net1696),
    .B1(_04746_),
    .X(_06005_));
 sg13g2_a21oi_1 _14349_ (.A1(_06004_),
    .A2(_06005_),
    .Y(_06006_),
    .B1(net2197));
 sg13g2_a21oi_1 _14350_ (.A1(net2329),
    .A2(net2197),
    .Y(_00590_),
    .B1(_06006_));
 sg13g2_nand2_1 _14351_ (.Y(_06007_),
    .A(_04715_),
    .B(_06005_));
 sg13g2_nor2_1 _14352_ (.A(_04715_),
    .B(_06005_),
    .Y(_06008_));
 sg13g2_nand3b_1 _14353_ (.B(_03108_),
    .C(_06007_),
    .Y(_06009_),
    .A_N(_06008_));
 sg13g2_o21ai_1 _14354_ (.B1(_06009_),
    .Y(_00591_),
    .A1(_01142_),
    .A2(_03108_));
 sg13g2_a21oi_2 _14355_ (.B1(_04818_),
    .Y(_06010_),
    .A2(_06003_),
    .A1(net1696));
 sg13g2_xor2_1 _14356_ (.B(_06008_),
    .A(_04716_),
    .X(_06011_));
 sg13g2_nand2_1 _14357_ (.Y(_06012_),
    .A(net3430),
    .B(net2197));
 sg13g2_o21ai_1 _14358_ (.B1(_06012_),
    .Y(_00592_),
    .A1(net2198),
    .A2(_06011_));
 sg13g2_nand2_1 _14359_ (.Y(_06013_),
    .A(_04720_),
    .B(_06010_));
 sg13g2_xnor2_1 _14360_ (.Y(_06014_),
    .A(_04719_),
    .B(_06010_));
 sg13g2_nor2_1 _14361_ (.A(net2197),
    .B(_06014_),
    .Y(_06015_));
 sg13g2_a21oi_1 _14362_ (.A1(_01144_),
    .A2(net2198),
    .Y(_00593_),
    .B1(_06015_));
 sg13g2_nor2_1 _14363_ (.A(net3704),
    .B(_03108_),
    .Y(_06016_));
 sg13g2_nor2_1 _14364_ (.A(_04712_),
    .B(_06013_),
    .Y(_06017_));
 sg13g2_xnor2_1 _14365_ (.Y(_06018_),
    .A(_04712_),
    .B(_06013_));
 sg13g2_a21oi_1 _14366_ (.A1(_03108_),
    .A2(_06018_),
    .Y(_00594_),
    .B1(net3705));
 sg13g2_and4_1 _14367_ (.A(_04711_),
    .B(_04713_),
    .C(_04720_),
    .D(_06010_),
    .X(_06019_));
 sg13g2_xnor2_1 _14368_ (.Y(_06020_),
    .A(_04711_),
    .B(_06017_));
 sg13g2_nand2_1 _14369_ (.Y(_06021_),
    .A(net3059),
    .B(net2198));
 sg13g2_o21ai_1 _14370_ (.B1(_06021_),
    .Y(_00595_),
    .A1(net2198),
    .A2(_06020_));
 sg13g2_a21oi_1 _14371_ (.A1(_04830_),
    .A2(_06010_),
    .Y(_06022_),
    .B1(_04725_));
 sg13g2_or2_1 _14372_ (.X(_06023_),
    .B(_04793_),
    .A(_04710_));
 sg13g2_o21ai_1 _14373_ (.B1(_04788_),
    .Y(_06024_),
    .A1(_06022_),
    .A2(_06023_));
 sg13g2_a21oi_1 _14374_ (.A1(_04830_),
    .A2(_06010_),
    .Y(_06025_),
    .B1(_04790_));
 sg13g2_o21ai_1 _14375_ (.B1(_06025_),
    .Y(_06026_),
    .A1(_04827_),
    .A2(_06019_));
 sg13g2_or2_1 _14376_ (.X(_06027_),
    .B(_06026_),
    .A(_06024_));
 sg13g2_a22oi_1 _14377_ (.Y(_00596_),
    .B1(_04795_),
    .B2(_06027_),
    .A2(net2197),
    .A1(_01148_));
 sg13g2_nor2_1 _14378_ (.A(_04794_),
    .B(_06024_),
    .Y(_06028_));
 sg13g2_nand3_1 _14379_ (.B(_04830_),
    .C(_06010_),
    .A(_04725_),
    .Y(_06029_));
 sg13g2_nor2_1 _14380_ (.A(_04790_),
    .B(_06022_),
    .Y(_06030_));
 sg13g2_nand2_1 _14381_ (.Y(_06031_),
    .A(_06029_),
    .B(_06030_));
 sg13g2_a22oi_1 _14382_ (.Y(_00597_),
    .B1(_06028_),
    .B2(_06031_),
    .A2(net2197),
    .A1(_01147_));
 sg13g2_a21o_1 _14383_ (.A2(_06029_),
    .A1(_04710_),
    .B1(_04790_),
    .X(_06032_));
 sg13g2_a22oi_1 _14384_ (.Y(_00598_),
    .B1(_06028_),
    .B2(_06032_),
    .A2(net2197),
    .A1(_01146_));
 sg13g2_nor2_1 _14385_ (.A(_03156_),
    .B(net1834),
    .Y(_06033_));
 sg13g2_and2_1 _14386_ (.A(_04302_),
    .B(_04788_),
    .X(_06034_));
 sg13g2_o21ai_1 _14387_ (.B1(_06034_),
    .Y(_06035_),
    .A1(_03132_),
    .A2(net1840));
 sg13g2_nor3_1 _14388_ (.A(net1776),
    .B(_06033_),
    .C(_06035_),
    .Y(_06036_));
 sg13g2_o21ai_1 _14389_ (.B1(_03133_),
    .Y(_06037_),
    .A1(_03444_),
    .A2(_03448_));
 sg13g2_a221oi_1 _14390_ (.B2(_03156_),
    .C1(_06036_),
    .B1(_06037_),
    .A1(_03132_),
    .Y(_06038_),
    .A2(_04787_));
 sg13g2_xnor2_1 _14391_ (.Y(_06039_),
    .A(_03133_),
    .B(net1729));
 sg13g2_nand4_1 _14392_ (.B(_04784_),
    .C(_06034_),
    .A(net1776),
    .Y(_06040_),
    .D(_06039_));
 sg13g2_a21oi_1 _14393_ (.A1(_06038_),
    .A2(_06040_),
    .Y(_06041_),
    .B1(_04794_));
 sg13g2_a21o_1 _14394_ (.A2(net2198),
    .A1(net2835),
    .B1(_06041_),
    .X(_00599_));
 sg13g2_o21ai_1 _14395_ (.B1(_02480_),
    .Y(_06042_),
    .A1(_02477_),
    .A2(net1861));
 sg13g2_nor2_2 _14396_ (.A(net1852),
    .B(_02749_),
    .Y(_06043_));
 sg13g2_nand2b_1 _14397_ (.Y(_06044_),
    .B(_02480_),
    .A_N(_02749_));
 sg13g2_nor2_1 _14398_ (.A(net2339),
    .B(net1815),
    .Y(_06045_));
 sg13g2_nand2_1 _14399_ (.Y(_06046_),
    .A(net2492),
    .B(net1816));
 sg13g2_nand3b_1 _14400_ (.B(_02536_),
    .C(net2138),
    .Y(_06047_),
    .A_N(net2137));
 sg13g2_nor2_1 _14401_ (.A(net2132),
    .B(_06047_),
    .Y(_06048_));
 sg13g2_or2_1 _14402_ (.X(_06049_),
    .B(_06047_),
    .A(net2132));
 sg13g2_nor2_2 _14403_ (.A(net2065),
    .B(net1973),
    .Y(_06050_));
 sg13g2_nand2b_1 _14404_ (.Y(_06051_),
    .B(net2134),
    .A_N(net2131));
 sg13g2_and2_1 _14405_ (.A(_02538_),
    .B(net2134),
    .X(_06052_));
 sg13g2_nand2_2 _14406_ (.Y(_06053_),
    .A(_02538_),
    .B(net2134));
 sg13g2_nand2b_1 _14407_ (.Y(_06054_),
    .B(_06052_),
    .A_N(net2132));
 sg13g2_nor2_2 _14408_ (.A(net2180),
    .B(net2214),
    .Y(_06055_));
 sg13g2_nand2_1 _14409_ (.Y(_06056_),
    .A(_02491_),
    .B(net2218));
 sg13g2_nor2_2 _14410_ (.A(_02491_),
    .B(net2218),
    .Y(_06057_));
 sg13g2_nor2_2 _14411_ (.A(_06055_),
    .B(_06057_),
    .Y(_06058_));
 sg13g2_mux4_1 _14412_ (.S0(net2183),
    .A0(\i_tinyqv.cpu.instr_data[1][4] ),
    .A1(\i_tinyqv.cpu.instr_data[3][4] ),
    .A2(\i_tinyqv.cpu.instr_data[2][4] ),
    .A3(\i_tinyqv.cpu.instr_data[0][4] ),
    .S1(net2215),
    .X(_06059_));
 sg13g2_nand3_1 _14413_ (.B(_06053_),
    .C(_06059_),
    .A(_02565_),
    .Y(_06060_));
 sg13g2_o21ai_1 _14414_ (.B1(_06060_),
    .Y(_06061_),
    .A1(_02552_),
    .A2(_06054_));
 sg13g2_nor3_2 _14415_ (.A(net2143),
    .B(_02527_),
    .C(_02529_),
    .Y(_06062_));
 sg13g2_nor2b_1 _14416_ (.A(net2130),
    .B_N(_06062_),
    .Y(_06063_));
 sg13g2_mux4_1 _14417_ (.S0(net2217),
    .A0(\i_tinyqv.cpu.instr_data[1][11] ),
    .A1(\i_tinyqv.cpu.instr_data[0][11] ),
    .A2(\i_tinyqv.cpu.instr_data[3][11] ),
    .A3(\i_tinyqv.cpu.instr_data[2][11] ),
    .S1(net2182),
    .X(_06064_));
 sg13g2_inv_1 _14418_ (.Y(_06065_),
    .A(_06064_));
 sg13g2_and2_1 _14419_ (.A(net2130),
    .B(_06064_),
    .X(_06066_));
 sg13g2_nand2_1 _14420_ (.Y(_06067_),
    .A(net2127),
    .B(_06066_));
 sg13g2_nor2_2 _14421_ (.A(_02772_),
    .B(_06067_),
    .Y(_06068_));
 sg13g2_nor2_1 _14422_ (.A(_02549_),
    .B(_02551_),
    .Y(_06069_));
 sg13g2_nand3b_1 _14423_ (.B(_06065_),
    .C(_06069_),
    .Y(_06070_),
    .A_N(net2129));
 sg13g2_inv_1 _14424_ (.Y(_06071_),
    .A(_06070_));
 sg13g2_a221oi_1 _14425_ (.B2(_02532_),
    .C1(_06068_),
    .B1(_06071_),
    .A1(net2131),
    .Y(_06072_),
    .A2(_06063_));
 sg13g2_a22oi_1 _14426_ (.Y(_06073_),
    .B1(net1955),
    .B2(_06061_),
    .A2(_02777_),
    .A1(_02536_));
 sg13g2_a21oi_1 _14427_ (.A1(_06072_),
    .A2(_06073_),
    .Y(_06074_),
    .B1(net1780));
 sg13g2_a21o_1 _14428_ (.A2(net1782),
    .A1(net3658),
    .B1(_06074_),
    .X(_00600_));
 sg13g2_nand2_2 _14429_ (.Y(_06075_),
    .A(net2139),
    .B(_02770_));
 sg13g2_nand2_1 _14430_ (.Y(_06076_),
    .A(_02562_),
    .B(_06075_));
 sg13g2_or2_1 _14431_ (.X(_06077_),
    .B(_06076_),
    .A(_02777_));
 sg13g2_nor2_2 _14432_ (.A(_02525_),
    .B(_02529_),
    .Y(_06078_));
 sg13g2_nand2b_1 _14433_ (.Y(_06079_),
    .B(net2139),
    .A_N(_02529_));
 sg13g2_nand2_2 _14434_ (.Y(_06080_),
    .A(_02498_),
    .B(net2141));
 sg13g2_nor2_2 _14435_ (.A(_06079_),
    .B(_06080_),
    .Y(_06081_));
 sg13g2_or2_1 _14436_ (.X(_06082_),
    .B(_06080_),
    .A(_06079_));
 sg13g2_and2_1 _14437_ (.A(_02498_),
    .B(_02757_),
    .X(_06083_));
 sg13g2_nor2_1 _14438_ (.A(_06081_),
    .B(_06083_),
    .Y(_06084_));
 sg13g2_nand2_2 _14439_ (.Y(_06085_),
    .A(net2144),
    .B(_06078_));
 sg13g2_nand2_1 _14440_ (.Y(_06086_),
    .A(_06084_),
    .B(_06085_));
 sg13g2_or4_1 _14441_ (.A(_02496_),
    .B(net2143),
    .C(net2142),
    .D(_02525_),
    .X(_06087_));
 sg13g2_nand2b_1 _14442_ (.Y(_06088_),
    .B(_06087_),
    .A_N(_06062_));
 sg13g2_nand3_1 _14443_ (.B(_02756_),
    .C(_02762_),
    .A(_02533_),
    .Y(_06089_));
 sg13g2_nor4_1 _14444_ (.A(_06077_),
    .B(_06086_),
    .C(_06088_),
    .D(_06089_),
    .Y(_06090_));
 sg13g2_a22oi_1 _14445_ (.Y(_06091_),
    .B1(_06077_),
    .B2(net2136),
    .A2(_06062_),
    .A1(net2134));
 sg13g2_nand2b_1 _14446_ (.Y(_06092_),
    .B(_06091_),
    .A_N(_06068_));
 sg13g2_o21ai_1 _14447_ (.B1(net2064),
    .Y(_06093_),
    .A1(_06090_),
    .A2(_06092_));
 sg13g2_nor2_1 _14448_ (.A(net2129),
    .B(_06053_),
    .Y(_06094_));
 sg13g2_mux4_1 _14449_ (.S0(net2183),
    .A0(\i_tinyqv.cpu.instr_data[1][5] ),
    .A1(\i_tinyqv.cpu.instr_data[3][5] ),
    .A2(\i_tinyqv.cpu.instr_data[2][5] ),
    .A3(\i_tinyqv.cpu.instr_data[0][5] ),
    .S1(net2215),
    .X(_06095_));
 sg13g2_o21ai_1 _14450_ (.B1(net1955),
    .Y(_06096_),
    .A1(_06052_),
    .A2(_06095_));
 sg13g2_o21ai_1 _14451_ (.B1(_06093_),
    .Y(_06097_),
    .A1(_06094_),
    .A2(_06096_));
 sg13g2_mux2_1 _14452_ (.A0(net2439),
    .A1(_06097_),
    .S(net1784),
    .X(_00601_));
 sg13g2_o21ai_1 _14453_ (.B1(_06077_),
    .Y(_06098_),
    .A1(net2138),
    .A2(_06068_));
 sg13g2_mux4_1 _14454_ (.S0(net2180),
    .A0(\i_tinyqv.cpu.instr_data[1][6] ),
    .A1(\i_tinyqv.cpu.instr_data[3][6] ),
    .A2(\i_tinyqv.cpu.instr_data[2][6] ),
    .A3(\i_tinyqv.cpu.instr_data[0][6] ),
    .S1(net2214),
    .X(_06099_));
 sg13g2_mux2_1 _14455_ (.A0(_02548_),
    .A1(_06099_),
    .S(_06053_),
    .X(_06100_));
 sg13g2_nor2b_1 _14456_ (.A(_06083_),
    .B_N(_06087_),
    .Y(_06101_));
 sg13g2_inv_1 _14457_ (.Y(_06102_),
    .A(_06101_));
 sg13g2_nand3_1 _14458_ (.B(_02548_),
    .C(_06078_),
    .A(net2143),
    .Y(_06103_));
 sg13g2_o21ai_1 _14459_ (.B1(_06103_),
    .Y(_06104_),
    .A1(_02766_),
    .A2(_02793_));
 sg13g2_a221oi_1 _14460_ (.B2(net2133),
    .C1(_06104_),
    .B1(_06102_),
    .A1(net1955),
    .Y(_06105_),
    .A2(_06100_));
 sg13g2_a21o_1 _14461_ (.A2(_06105_),
    .A1(_06098_),
    .B1(net1780),
    .X(_06106_));
 sg13g2_o21ai_1 _14462_ (.B1(_06106_),
    .Y(_00602_),
    .A1(_01070_),
    .A2(net1784));
 sg13g2_or2_1 _14463_ (.X(_06107_),
    .B(_06083_),
    .A(_02561_));
 sg13g2_nand2b_1 _14464_ (.Y(_06108_),
    .B(_02766_),
    .A_N(_06107_));
 sg13g2_o21ai_1 _14465_ (.B1(net2135),
    .Y(_06109_),
    .A1(_02777_),
    .A2(_06108_));
 sg13g2_mux4_1 _14466_ (.S0(net2182),
    .A0(\i_tinyqv.cpu.instr_data[1][7] ),
    .A1(\i_tinyqv.cpu.instr_data[3][7] ),
    .A2(\i_tinyqv.cpu.instr_data[2][7] ),
    .A3(\i_tinyqv.cpu.instr_data[0][7] ),
    .S1(net2214),
    .X(_06110_));
 sg13g2_mux2_1 _14467_ (.A0(_02547_),
    .A1(_06110_),
    .S(_06053_),
    .X(_06111_));
 sg13g2_nand2_1 _14468_ (.Y(_06112_),
    .A(_06075_),
    .B(_06087_));
 sg13g2_nand3_1 _14469_ (.B(_06085_),
    .C(_06087_),
    .A(_06075_),
    .Y(_06113_));
 sg13g2_a221oi_1 _14470_ (.B2(_02547_),
    .C1(_06068_),
    .B1(_06113_),
    .A1(net1955),
    .Y(_06114_),
    .A2(_06111_));
 sg13g2_a21oi_1 _14471_ (.A1(_06109_),
    .A2(_06114_),
    .Y(_06115_),
    .B1(net1780));
 sg13g2_a21o_1 _14472_ (.A2(net1782),
    .A1(net4007),
    .B1(_06115_),
    .X(_00603_));
 sg13g2_nand2_1 _14473_ (.Y(_06116_),
    .A(_02562_),
    .B(_06084_));
 sg13g2_o21ai_1 _14474_ (.B1(_06064_),
    .Y(_06117_),
    .A1(_06113_),
    .A2(_06116_));
 sg13g2_o21ai_1 _14475_ (.B1(_02780_),
    .Y(_06118_),
    .A1(net2133),
    .A2(_06068_));
 sg13g2_nand2_1 _14476_ (.Y(_06119_),
    .A(net2129),
    .B(_06069_));
 sg13g2_nor2_2 _14477_ (.A(_02762_),
    .B(_06119_),
    .Y(_06120_));
 sg13g2_or2_1 _14478_ (.X(_06121_),
    .B(_06119_),
    .A(_02762_));
 sg13g2_a22oi_1 _14479_ (.Y(_06122_),
    .B1(net2214),
    .B2(\i_tinyqv.cpu.instr_data[2][8] ),
    .A2(net2180),
    .A1(\i_tinyqv.cpu.instr_data[3][8] ));
 sg13g2_a22oi_1 _14480_ (.Y(_06123_),
    .B1(_06058_),
    .B2(_06122_),
    .A2(_06057_),
    .A1(_01096_));
 sg13g2_o21ai_1 _14481_ (.B1(_06123_),
    .Y(_06124_),
    .A1(\i_tinyqv.cpu.instr_data[1][8] ),
    .A2(_06056_));
 sg13g2_nand2_1 _14482_ (.Y(_06125_),
    .A(_06052_),
    .B(_06064_));
 sg13g2_o21ai_1 _14483_ (.B1(_06125_),
    .Y(_06126_),
    .A1(_06052_),
    .A2(_06124_));
 sg13g2_a22oi_1 _14484_ (.Y(_06127_),
    .B1(_06126_),
    .B2(net1955),
    .A2(_06120_),
    .A1(net2133));
 sg13g2_nand3_1 _14485_ (.B(_06118_),
    .C(_06127_),
    .A(_06117_),
    .Y(_06128_));
 sg13g2_mux2_1 _14486_ (.A0(net4009),
    .A1(_06128_),
    .S(net1785),
    .X(_00604_));
 sg13g2_nand2_1 _14487_ (.Y(_06129_),
    .A(_02775_),
    .B(_06121_));
 sg13g2_o21ai_1 _14488_ (.B1(_02536_),
    .Y(_06130_),
    .A1(_06076_),
    .A2(_06129_));
 sg13g2_nand3_1 _14489_ (.B(_06085_),
    .C(_06101_),
    .A(_02766_),
    .Y(_06131_));
 sg13g2_mux4_1 _14490_ (.S0(net2182),
    .A0(\i_tinyqv.cpu.instr_data[1][9] ),
    .A1(\i_tinyqv.cpu.instr_data[3][9] ),
    .A2(\i_tinyqv.cpu.instr_data[2][9] ),
    .A3(\i_tinyqv.cpu.instr_data[0][9] ),
    .S1(net2215),
    .X(_06132_));
 sg13g2_nand2_1 _14491_ (.Y(_06133_),
    .A(net2071),
    .B(_06132_));
 sg13g2_inv_1 _14492_ (.Y(_06134_),
    .A(_06133_));
 sg13g2_a22oi_1 _14493_ (.Y(_06135_),
    .B1(_06134_),
    .B2(_06049_),
    .A2(_06081_),
    .A1(net2130));
 sg13g2_o21ai_1 _14494_ (.B1(net2128),
    .Y(_06136_),
    .A1(_02777_),
    .A2(_06131_));
 sg13g2_nand4_1 _14495_ (.B(_06130_),
    .C(_06135_),
    .A(net1791),
    .Y(_06137_),
    .D(_06136_));
 sg13g2_o21ai_1 _14496_ (.B1(_06137_),
    .Y(_06138_),
    .A1(net4043),
    .A2(net1784));
 sg13g2_inv_1 _14497_ (.Y(_00605_),
    .A(_06138_));
 sg13g2_o21ai_1 _14498_ (.B1(net2135),
    .Y(_06139_),
    .A1(_06112_),
    .A2(_06129_));
 sg13g2_o21ai_1 _14499_ (.B1(_02551_),
    .Y(_06140_),
    .A1(_02561_),
    .A2(_06086_));
 sg13g2_nor2_1 _14500_ (.A(_02537_),
    .B(_02766_),
    .Y(_06141_));
 sg13g2_mux4_1 _14501_ (.S0(net2183),
    .A0(\i_tinyqv.cpu.instr_data[1][10] ),
    .A1(\i_tinyqv.cpu.instr_data[3][10] ),
    .A2(\i_tinyqv.cpu.instr_data[2][10] ),
    .A3(\i_tinyqv.cpu.instr_data[0][10] ),
    .S1(net2215),
    .X(_06142_));
 sg13g2_a221oi_1 _14502_ (.B2(_06142_),
    .C1(_06141_),
    .B1(net1955),
    .A1(net2128),
    .Y(_06143_),
    .A2(_02777_));
 sg13g2_nand3_1 _14503_ (.B(_06140_),
    .C(_06143_),
    .A(_06139_),
    .Y(_06144_));
 sg13g2_mux2_1 _14504_ (.A0(net4048),
    .A1(_06144_),
    .S(net1784),
    .X(_00606_));
 sg13g2_nand2_1 _14505_ (.Y(_06145_),
    .A(_02779_),
    .B(_06121_));
 sg13g2_a22oi_1 _14506_ (.Y(_06146_),
    .B1(_06145_),
    .B2(net2137),
    .A2(_06086_),
    .A1(net2129));
 sg13g2_mux4_1 _14507_ (.S0(net2182),
    .A0(\i_tinyqv.cpu.instr_data[1][11] ),
    .A1(\i_tinyqv.cpu.instr_data[3][11] ),
    .A2(\i_tinyqv.cpu.instr_data[2][11] ),
    .A3(\i_tinyqv.cpu.instr_data[0][11] ),
    .S1(net2215),
    .X(_06147_));
 sg13g2_a22oi_1 _14508_ (.Y(_06148_),
    .B1(_06076_),
    .B2(net2133),
    .A2(_02777_),
    .A1(net2126));
 sg13g2_nand2_1 _14509_ (.Y(_06149_),
    .A(_06146_),
    .B(_06148_));
 sg13g2_a21oi_1 _14510_ (.A1(net1955),
    .A2(_06147_),
    .Y(_06150_),
    .B1(_06149_));
 sg13g2_nor2_1 _14511_ (.A(net3891),
    .B(net1790),
    .Y(_06151_));
 sg13g2_a21oi_1 _14512_ (.A1(net1790),
    .A2(_06150_),
    .Y(_00607_),
    .B1(_06151_));
 sg13g2_nand3_1 _14513_ (.B(net2126),
    .C(_02771_),
    .A(net2136),
    .Y(_06152_));
 sg13g2_nand2_1 _14514_ (.Y(_06153_),
    .A(_02759_),
    .B(net1940));
 sg13g2_a21oi_1 _14515_ (.A1(_06047_),
    .A2(_06066_),
    .Y(_06154_),
    .B1(_02772_));
 sg13g2_o21ai_1 _14516_ (.B1(net2127),
    .Y(_06155_),
    .A1(_06153_),
    .A2(_06154_));
 sg13g2_and2_1 _14517_ (.A(_06152_),
    .B(_06155_),
    .X(_06156_));
 sg13g2_o21ai_1 _14518_ (.B1(net2126),
    .Y(_06157_),
    .A1(_06081_),
    .A2(_06120_));
 sg13g2_nand2_1 _14519_ (.Y(_06158_),
    .A(net2126),
    .B(_02774_));
 sg13g2_nand3_1 _14520_ (.B(_06157_),
    .C(_06158_),
    .A(_06156_),
    .Y(_06159_));
 sg13g2_mux4_1 _14521_ (.S0(net2185),
    .A0(\i_tinyqv.cpu.instr_data[1][14] ),
    .A1(\i_tinyqv.cpu.instr_data[3][14] ),
    .A2(\i_tinyqv.cpu.instr_data[2][14] ),
    .A3(\i_tinyqv.cpu.instr_data[0][14] ),
    .S1(net2216),
    .X(_06160_));
 sg13g2_and2_1 _14522_ (.A(net2067),
    .B(_06160_),
    .X(_06161_));
 sg13g2_a221oi_1 _14523_ (.B2(_06161_),
    .C1(_06159_),
    .B1(net1972),
    .A1(net2129),
    .Y(_06162_),
    .A2(_02561_));
 sg13g2_nor2_1 _14524_ (.A(net3979),
    .B(net1785),
    .Y(_06163_));
 sg13g2_a21oi_1 _14525_ (.A1(net1784),
    .A2(_06162_),
    .Y(_00608_),
    .B1(_06163_));
 sg13g2_o21ai_1 _14526_ (.B1(net2126),
    .Y(_06164_),
    .A1(_02561_),
    .A2(_02774_));
 sg13g2_and2_1 _14527_ (.A(_06156_),
    .B(_06164_),
    .X(_06165_));
 sg13g2_mux4_1 _14528_ (.S0(net2185),
    .A0(\i_tinyqv.cpu.instr_data[1][15] ),
    .A1(\i_tinyqv.cpu.instr_data[3][15] ),
    .A2(\i_tinyqv.cpu.instr_data[2][15] ),
    .A3(\i_tinyqv.cpu.instr_data[0][15] ),
    .S1(net2214),
    .X(_06166_));
 sg13g2_nand2_1 _14529_ (.Y(_06167_),
    .A(_02565_),
    .B(_06166_));
 sg13g2_inv_1 _14530_ (.Y(_06168_),
    .A(_06167_));
 sg13g2_nor2_1 _14531_ (.A(_02539_),
    .B(_02563_),
    .Y(_06169_));
 sg13g2_nand2_2 _14532_ (.Y(_06170_),
    .A(net2132),
    .B(_06052_));
 sg13g2_nand3_1 _14533_ (.B(_02564_),
    .C(_06059_),
    .A(net2136),
    .Y(_06171_));
 sg13g2_nand3_1 _14534_ (.B(_06170_),
    .C(_06171_),
    .A(_06167_),
    .Y(_06172_));
 sg13g2_o21ai_1 _14535_ (.B1(_06050_),
    .Y(_06173_),
    .A1(_02551_),
    .A2(_06170_));
 sg13g2_nand2b_1 _14536_ (.Y(_06174_),
    .B(_06172_),
    .A_N(_06173_));
 sg13g2_nand4_1 _14537_ (.B(_06157_),
    .C(_06165_),
    .A(net1791),
    .Y(_06175_),
    .D(_06174_));
 sg13g2_o21ai_1 _14538_ (.B1(_06175_),
    .Y(_06176_),
    .A1(net4089),
    .A2(net1788));
 sg13g2_inv_1 _14539_ (.Y(_00609_),
    .A(_06176_));
 sg13g2_nor2_1 _14540_ (.A(net3907),
    .B(net1785),
    .Y(_06177_));
 sg13g2_nand2_1 _14541_ (.Y(_06178_),
    .A(net2067),
    .B(_06166_));
 sg13g2_nand2_1 _14542_ (.Y(_06179_),
    .A(_06050_),
    .B(_06168_));
 sg13g2_nand3_1 _14543_ (.B(_06165_),
    .C(_06179_),
    .A(_06157_),
    .Y(_06180_));
 sg13g2_nor2b_2 _14544_ (.A(_02762_),
    .B_N(_06119_),
    .Y(_06181_));
 sg13g2_nand2_2 _14545_ (.Y(_06182_),
    .A(_02565_),
    .B(net1972));
 sg13g2_inv_1 _14546_ (.Y(_06183_),
    .A(_06182_));
 sg13g2_and2_1 _14547_ (.A(net2067),
    .B(net2126),
    .X(_06184_));
 sg13g2_a221oi_1 _14548_ (.B2(_06184_),
    .C1(_06180_),
    .B1(_06182_),
    .A1(_02536_),
    .Y(_06185_),
    .A2(_06181_));
 sg13g2_a21oi_1 _14549_ (.A1(net1785),
    .A2(_06185_),
    .Y(_00610_),
    .B1(_06177_));
 sg13g2_nor2_1 _14550_ (.A(net3904),
    .B(net1791),
    .Y(_06186_));
 sg13g2_and2_1 _14551_ (.A(net2067),
    .B(net2141),
    .X(_06187_));
 sg13g2_a221oi_1 _14552_ (.B2(_06187_),
    .C1(_06180_),
    .B1(_06182_),
    .A1(net2136),
    .Y(_06188_),
    .A2(_06181_));
 sg13g2_a21oi_1 _14553_ (.A1(net1792),
    .A2(_06188_),
    .Y(_00611_),
    .B1(_06186_));
 sg13g2_nand2_1 _14554_ (.Y(_06189_),
    .A(net2140),
    .B(_06182_));
 sg13g2_a21oi_1 _14555_ (.A1(net1972),
    .A2(_06168_),
    .Y(_06190_),
    .B1(net2065));
 sg13g2_nand2_1 _14556_ (.Y(_06191_),
    .A(net2065),
    .B(_06157_));
 sg13g2_a21oi_1 _14557_ (.A1(net2138),
    .A2(_06181_),
    .Y(_06192_),
    .B1(_06191_));
 sg13g2_a221oi_1 _14558_ (.B2(_06165_),
    .C1(net1780),
    .B1(_06192_),
    .A1(_06189_),
    .Y(_06193_),
    .A2(_06190_));
 sg13g2_a21o_1 _14559_ (.A2(net1781),
    .A1(net3998),
    .B1(_06193_),
    .X(_00612_));
 sg13g2_nand2_1 _14560_ (.Y(_06194_),
    .A(_02528_),
    .B(_06182_));
 sg13g2_a21oi_1 _14561_ (.A1(net2134),
    .A2(_06181_),
    .Y(_06195_),
    .B1(_06191_));
 sg13g2_a22oi_1 _14562_ (.Y(_06196_),
    .B1(_06195_),
    .B2(_06165_),
    .A2(_06194_),
    .A1(_06190_));
 sg13g2_nand2_1 _14563_ (.Y(_06197_),
    .A(net1788),
    .B(_06196_));
 sg13g2_o21ai_1 _14564_ (.B1(_06197_),
    .Y(_00613_),
    .A1(_01068_),
    .A2(net1784));
 sg13g2_a22oi_1 _14565_ (.Y(_06198_),
    .B1(net2214),
    .B2(_01090_),
    .A2(net2180),
    .A1(_01089_));
 sg13g2_nor2_1 _14566_ (.A(_01087_),
    .B(_06056_),
    .Y(_06199_));
 sg13g2_a221oi_1 _14567_ (.B2(_06198_),
    .C1(_06199_),
    .B1(_06058_),
    .A1(\i_tinyqv.cpu.instr_data[0][0] ),
    .Y(_06200_),
    .A2(_06057_));
 sg13g2_o21ai_1 _14568_ (.B1(_06190_),
    .Y(_06201_),
    .A1(_06183_),
    .A2(_06200_));
 sg13g2_a21oi_1 _14569_ (.A1(net2132),
    .A2(_06181_),
    .Y(_06202_),
    .B1(_06191_));
 sg13g2_nand3_1 _14570_ (.B(_06164_),
    .C(_06202_),
    .A(_06155_),
    .Y(_06203_));
 sg13g2_nand3_1 _14571_ (.B(_06201_),
    .C(_06203_),
    .A(net1791),
    .Y(_06204_));
 sg13g2_o21ai_1 _14572_ (.B1(_06204_),
    .Y(_00614_),
    .A1(_01074_),
    .A2(net1785));
 sg13g2_o21ai_1 _14573_ (.B1(net2127),
    .Y(_06205_),
    .A1(_02763_),
    .A2(_06081_));
 sg13g2_and3_2 _14574_ (.X(_06206_),
    .A(_06155_),
    .B(_06164_),
    .C(_06205_));
 sg13g2_nand2_1 _14575_ (.Y(_06207_),
    .A(_06179_),
    .B(_06206_));
 sg13g2_a22oi_1 _14576_ (.Y(_06208_),
    .B1(net2214),
    .B2(_01094_),
    .A2(net2180),
    .A1(_01093_));
 sg13g2_nand2_1 _14577_ (.Y(_06209_),
    .A(_06058_),
    .B(_06208_));
 sg13g2_a22oi_1 _14578_ (.Y(_06210_),
    .B1(_06057_),
    .B2(\i_tinyqv.cpu.instr_data[0][1] ),
    .A2(_06055_),
    .A1(\i_tinyqv.cpu.instr_data[1][1] ));
 sg13g2_a21oi_2 _14579_ (.B1(net2065),
    .Y(_06211_),
    .A2(_06210_),
    .A1(_06209_));
 sg13g2_a21oi_1 _14580_ (.A1(_06182_),
    .A2(_06211_),
    .Y(_06212_),
    .B1(_06207_));
 sg13g2_nor2_1 _14581_ (.A(net3911),
    .B(net1784),
    .Y(_06213_));
 sg13g2_a21oi_1 _14582_ (.A1(net1785),
    .A2(_06212_),
    .Y(_00615_),
    .B1(_06213_));
 sg13g2_nor2_1 _14583_ (.A(\i_tinyqv.cpu.instr_data[2][2] ),
    .B(net2180),
    .Y(_06214_));
 sg13g2_o21ai_1 _14584_ (.B1(_06058_),
    .Y(_06215_),
    .A1(\i_tinyqv.cpu.instr_data[3][2] ),
    .A2(_02491_));
 sg13g2_a22oi_1 _14585_ (.Y(_06216_),
    .B1(_06057_),
    .B2(\i_tinyqv.cpu.instr_data[0][2] ),
    .A2(_06055_),
    .A1(\i_tinyqv.cpu.instr_data[1][2] ));
 sg13g2_o21ai_1 _14586_ (.B1(_06216_),
    .Y(_06217_),
    .A1(_06214_),
    .A2(_06215_));
 sg13g2_nand2_1 _14587_ (.Y(_06218_),
    .A(net2071),
    .B(_06217_));
 sg13g2_inv_1 _14588_ (.Y(_06219_),
    .A(_06218_));
 sg13g2_a21oi_1 _14589_ (.A1(_06182_),
    .A2(_06219_),
    .Y(_06220_),
    .B1(_06207_));
 sg13g2_nor2_1 _14590_ (.A(net3919),
    .B(net1791),
    .Y(_06221_));
 sg13g2_a21oi_1 _14591_ (.A1(net1791),
    .A2(_06220_),
    .Y(_00616_),
    .B1(_06221_));
 sg13g2_mux2_1 _14592_ (.A0(\i_tinyqv.cpu.instr_data[3][3] ),
    .A1(\i_tinyqv.cpu.instr_data[2][3] ),
    .S(_02491_),
    .X(_06222_));
 sg13g2_nand2_1 _14593_ (.Y(_06223_),
    .A(_06058_),
    .B(_06222_));
 sg13g2_a22oi_1 _14594_ (.Y(_06224_),
    .B1(_06057_),
    .B2(\i_tinyqv.cpu.instr_data[0][3] ),
    .A2(_06055_),
    .A1(\i_tinyqv.cpu.instr_data[1][3] ));
 sg13g2_a21oi_1 _14595_ (.A1(_06223_),
    .A2(_06224_),
    .Y(_06225_),
    .B1(_02500_));
 sg13g2_a21oi_1 _14596_ (.A1(_06182_),
    .A2(_06225_),
    .Y(_06226_),
    .B1(_06207_));
 sg13g2_nor2_1 _14597_ (.A(net3831),
    .B(net1786),
    .Y(_06227_));
 sg13g2_a21oi_1 _14598_ (.A1(net1786),
    .A2(_06226_),
    .Y(_00617_),
    .B1(_06227_));
 sg13g2_o21ai_1 _14599_ (.B1(_06206_),
    .Y(_06228_),
    .A1(net1973),
    .A2(_06178_));
 sg13g2_and2_1 _14600_ (.A(net2067),
    .B(_06059_),
    .X(_06229_));
 sg13g2_a21oi_1 _14601_ (.A1(net1973),
    .A2(_06229_),
    .Y(_06230_),
    .B1(_06228_));
 sg13g2_nor2_1 _14602_ (.A(net3847),
    .B(net1789),
    .Y(_06231_));
 sg13g2_a21oi_1 _14603_ (.A1(net1789),
    .A2(_06230_),
    .Y(_00618_),
    .B1(_06231_));
 sg13g2_nand2_2 _14604_ (.Y(_06232_),
    .A(net2070),
    .B(_06095_));
 sg13g2_nor2_1 _14605_ (.A(net1972),
    .B(_06232_),
    .Y(_06233_));
 sg13g2_nor3_1 _14606_ (.A(net1780),
    .B(_06228_),
    .C(_06233_),
    .Y(_06234_));
 sg13g2_a21oi_1 _14607_ (.A1(_01072_),
    .A2(net1782),
    .Y(_00619_),
    .B1(_06234_));
 sg13g2_nand2_2 _14608_ (.Y(_06235_),
    .A(net2070),
    .B(_06099_));
 sg13g2_nor2_1 _14609_ (.A(net1972),
    .B(_06235_),
    .Y(_06236_));
 sg13g2_nor3_1 _14610_ (.A(net1780),
    .B(net1899),
    .C(_06236_),
    .Y(_06237_));
 sg13g2_a21oi_1 _14611_ (.A1(_01071_),
    .A2(net1781),
    .Y(_00620_),
    .B1(_06237_));
 sg13g2_nand2_2 _14612_ (.Y(_06238_),
    .A(net2071),
    .B(_06110_));
 sg13g2_nor2_1 _14613_ (.A(net1972),
    .B(_06238_),
    .Y(_06239_));
 sg13g2_nor3_1 _14614_ (.A(net1780),
    .B(_06228_),
    .C(_06239_),
    .Y(_06240_));
 sg13g2_a21oi_1 _14615_ (.A1(_01069_),
    .A2(net1781),
    .Y(_00621_),
    .B1(_06240_));
 sg13g2_nor3_1 _14616_ (.A(net2065),
    .B(net1972),
    .C(_06124_),
    .Y(_06241_));
 sg13g2_nor3_1 _14617_ (.A(net1781),
    .B(net1899),
    .C(_06241_),
    .Y(_06242_));
 sg13g2_a21oi_1 _14618_ (.A1(_01075_),
    .A2(net1782),
    .Y(_00622_),
    .B1(_06242_));
 sg13g2_a21oi_1 _14619_ (.A1(net1973),
    .A2(_06134_),
    .Y(_06243_),
    .B1(net1899));
 sg13g2_nor2_1 _14620_ (.A(net3071),
    .B(net1789),
    .Y(_06244_));
 sg13g2_a21oi_1 _14621_ (.A1(net1789),
    .A2(_06243_),
    .Y(_00623_),
    .B1(_06244_));
 sg13g2_nand3_1 _14622_ (.B(net1973),
    .C(_06142_),
    .A(net2067),
    .Y(_06245_));
 sg13g2_nor2b_1 _14623_ (.A(net1899),
    .B_N(_06245_),
    .Y(_06246_));
 sg13g2_nor2_1 _14624_ (.A(net3053),
    .B(net1789),
    .Y(_06247_));
 sg13g2_a21oi_1 _14625_ (.A1(net1786),
    .A2(_06246_),
    .Y(_00624_),
    .B1(_06247_));
 sg13g2_nand3_1 _14626_ (.B(net1973),
    .C(_06147_),
    .A(net2067),
    .Y(_06248_));
 sg13g2_nor2b_1 _14627_ (.A(net1899),
    .B_N(_06248_),
    .Y(_06249_));
 sg13g2_nor2_1 _14628_ (.A(net3042),
    .B(net1787),
    .Y(_06250_));
 sg13g2_a21oi_1 _14629_ (.A1(net1787),
    .A2(_06249_),
    .Y(_00625_),
    .B1(_06250_));
 sg13g2_mux4_1 _14630_ (.S0(net2181),
    .A0(\i_tinyqv.cpu.instr_data[1][12] ),
    .A1(\i_tinyqv.cpu.instr_data[3][12] ),
    .A2(\i_tinyqv.cpu.instr_data[2][12] ),
    .A3(\i_tinyqv.cpu.instr_data[0][12] ),
    .S1(net2214),
    .X(_06251_));
 sg13g2_nand3_1 _14631_ (.B(net1973),
    .C(_06251_),
    .A(net2067),
    .Y(_06252_));
 sg13g2_nor2b_1 _14632_ (.A(net1899),
    .B_N(_06252_),
    .Y(_06253_));
 sg13g2_nor2_1 _14633_ (.A(net2834),
    .B(net1786),
    .Y(_06254_));
 sg13g2_a21oi_1 _14634_ (.A1(net1786),
    .A2(_06253_),
    .Y(_00626_),
    .B1(_06254_));
 sg13g2_mux4_1 _14635_ (.S0(net2183),
    .A0(\i_tinyqv.cpu.instr_data[1][13] ),
    .A1(\i_tinyqv.cpu.instr_data[3][13] ),
    .A2(\i_tinyqv.cpu.instr_data[2][13] ),
    .A3(\i_tinyqv.cpu.instr_data[0][13] ),
    .S1(net2215),
    .X(_06255_));
 sg13g2_nand3_1 _14636_ (.B(_06048_),
    .C(_06255_),
    .A(net2068),
    .Y(_06256_));
 sg13g2_nor2b_1 _14637_ (.A(net1899),
    .B_N(_06256_),
    .Y(_06257_));
 sg13g2_nor2_1 _14638_ (.A(net3133),
    .B(net1787),
    .Y(_06258_));
 sg13g2_a21oi_1 _14639_ (.A1(net1787),
    .A2(_06257_),
    .Y(_00627_),
    .B1(_06258_));
 sg13g2_a21oi_1 _14640_ (.A1(net1973),
    .A2(_06161_),
    .Y(_06259_),
    .B1(net1899));
 sg13g2_nor2_1 _14641_ (.A(net3039),
    .B(net1786),
    .Y(_06260_));
 sg13g2_a21oi_1 _14642_ (.A1(net1786),
    .A2(_06259_),
    .Y(_00628_),
    .B1(_06260_));
 sg13g2_nand3_1 _14643_ (.B(_06178_),
    .C(_06206_),
    .A(net1791),
    .Y(_06261_));
 sg13g2_o21ai_1 _14644_ (.B1(_06261_),
    .Y(_06262_),
    .A1(net3631),
    .A2(net1786));
 sg13g2_inv_1 _14645_ (.Y(_00629_),
    .A(_06262_));
 sg13g2_a22oi_1 _14646_ (.Y(_06263_),
    .B1(_06129_),
    .B2(net2138),
    .A2(_06116_),
    .A1(_02548_));
 sg13g2_nand2_1 _14647_ (.Y(_06264_),
    .A(_06156_),
    .B(_06263_));
 sg13g2_a21oi_2 _14648_ (.B1(_06264_),
    .Y(_06265_),
    .A2(_06251_),
    .A1(_06050_));
 sg13g2_o21ai_1 _14649_ (.B1(net2490),
    .Y(_06266_),
    .A1(net4097),
    .A2(net1818));
 sg13g2_a21oi_1 _14650_ (.A1(net1818),
    .A2(_06265_),
    .Y(_00630_),
    .B1(_06266_));
 sg13g2_and2_1 _14651_ (.A(net2064),
    .B(net2130),
    .X(_06267_));
 sg13g2_a221oi_1 _14652_ (.B2(_06107_),
    .C1(_06159_),
    .B1(_06267_),
    .A1(net1955),
    .Y(_06268_),
    .A2(_06255_));
 sg13g2_o21ai_1 _14653_ (.B1(net2493),
    .Y(_06269_),
    .A1(net4118),
    .A2(net1816));
 sg13g2_a21oi_1 _14654_ (.A1(net1816),
    .A2(_06268_),
    .Y(_00631_),
    .B1(_06269_));
 sg13g2_and2_1 _14655_ (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .B(net1855),
    .X(_06270_));
 sg13g2_mux2_1 _14656_ (.A0(\i_tinyqv.cpu.i_core.mepc[1] ),
    .A1(net2463),
    .S(net2222),
    .X(_06271_));
 sg13g2_nor2_1 _14657_ (.A(net2240),
    .B(_06271_),
    .Y(_06272_));
 sg13g2_a21oi_1 _14658_ (.A1(net2240),
    .A2(_05287_),
    .Y(_06273_),
    .B1(_06272_));
 sg13g2_a22oi_1 _14659_ (.Y(_06274_),
    .B1(_06273_),
    .B2(net1862),
    .A2(_06270_),
    .A1(net1812));
 sg13g2_o21ai_1 _14660_ (.B1(_06274_),
    .Y(_06275_),
    .A1(_02581_),
    .A2(_02639_));
 sg13g2_and2_1 _14661_ (.A(net2494),
    .B(_06275_),
    .X(_00632_));
 sg13g2_mux2_1 _14662_ (.A0(\i_tinyqv.cpu.i_core.mepc[2] ),
    .A1(net2462),
    .S(net2223),
    .X(_06276_));
 sg13g2_nor2_1 _14663_ (.A(net2306),
    .B(_05294_),
    .Y(_06277_));
 sg13g2_a21oi_1 _14664_ (.A1(net2306),
    .A2(_06276_),
    .Y(_06278_),
    .B1(_06277_));
 sg13g2_a21oi_1 _14665_ (.A1(net1862),
    .A2(_06278_),
    .Y(_06279_),
    .B1(net2342));
 sg13g2_o21ai_1 _14666_ (.B1(_06279_),
    .Y(_06280_),
    .A1(net2746),
    .A2(net1862));
 sg13g2_nand2b_1 _14667_ (.Y(_06281_),
    .B(_02639_),
    .A_N(_06280_));
 sg13g2_o21ai_1 _14668_ (.B1(_06281_),
    .Y(_00633_),
    .A1(net4153),
    .A2(_02640_));
 sg13g2_nand2_1 _14669_ (.Y(_06282_),
    .A(net2417),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ));
 sg13g2_nor2_1 _14670_ (.A(net2417),
    .B(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .Y(_06283_));
 sg13g2_xor2_1 _14671_ (.B(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .A(\i_tinyqv.cpu.instr_data_start[4] ),
    .X(_06284_));
 sg13g2_a21oi_1 _14672_ (.A1(net2418),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .Y(_06285_),
    .B1(_05300_));
 sg13g2_xnor2_1 _14673_ (.Y(_06286_),
    .A(_06284_),
    .B(_06285_));
 sg13g2_and3_1 _14674_ (.X(_06287_),
    .A(net2417),
    .B(net2418),
    .C(\i_tinyqv.cpu.instr_write_offset[3] ));
 sg13g2_a21oi_1 _14675_ (.A1(net2418),
    .A2(\i_tinyqv.cpu.instr_write_offset[3] ),
    .Y(_06288_),
    .B1(net2417));
 sg13g2_nor3_1 _14676_ (.A(net2407),
    .B(_06287_),
    .C(_06288_),
    .Y(_06289_));
 sg13g2_a21oi_1 _14677_ (.A1(net2407),
    .A2(_06286_),
    .Y(_06290_),
    .B1(_06289_));
 sg13g2_a22oi_1 _14678_ (.Y(_06291_),
    .B1(net2063),
    .B2(net2385),
    .A2(_02807_),
    .A1(net2781));
 sg13g2_o21ai_1 _14679_ (.B1(_06291_),
    .Y(_06292_),
    .A1(_05285_),
    .A2(_06290_));
 sg13g2_mux2_1 _14680_ (.A0(_06292_),
    .A1(net3149),
    .S(net1743),
    .X(_00634_));
 sg13g2_xnor2_1 _14681_ (.Y(_06293_),
    .A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[5] ));
 sg13g2_o21ai_1 _14682_ (.B1(_06282_),
    .Y(_06294_),
    .A1(_06283_),
    .A2(_06285_));
 sg13g2_nor2b_1 _14683_ (.A(_06293_),
    .B_N(_06294_),
    .Y(_06295_));
 sg13g2_xnor2_1 _14684_ (.Y(_06296_),
    .A(_06293_),
    .B(_06294_));
 sg13g2_and2_1 _14685_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(_06287_),
    .X(_06297_));
 sg13g2_nor2_1 _14686_ (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .B(_06287_),
    .Y(_06298_));
 sg13g2_nor3_1 _14687_ (.A(net2407),
    .B(_06297_),
    .C(_06298_),
    .Y(_06299_));
 sg13g2_a21oi_1 _14688_ (.A1(net2407),
    .A2(_06296_),
    .Y(_06300_),
    .B1(_06299_));
 sg13g2_a22oi_1 _14689_ (.Y(_06301_),
    .B1(net2062),
    .B2(\addr[5] ),
    .A2(net1752),
    .A1(\i_tinyqv.mem.q_ctrl.addr[1] ));
 sg13g2_o21ai_1 _14690_ (.B1(_06301_),
    .Y(_06302_),
    .A1(_05285_),
    .A2(_06300_));
 sg13g2_mux2_1 _14691_ (.A0(_06302_),
    .A1(net3164),
    .S(net1746),
    .X(_00635_));
 sg13g2_and2_1 _14692_ (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(_06297_),
    .X(_06303_));
 sg13g2_xnor2_1 _14693_ (.Y(_06304_),
    .A(_00981_),
    .B(_06297_));
 sg13g2_a21oi_1 _14694_ (.A1(\i_tinyqv.cpu.instr_data_start[5] ),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .Y(_06305_),
    .B1(_06295_));
 sg13g2_nand2_1 _14695_ (.Y(_06306_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_nor2_1 _14696_ (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .Y(_06307_));
 sg13g2_xnor2_1 _14697_ (.Y(_06308_),
    .A(\i_tinyqv.cpu.instr_data_start[6] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[6] ));
 sg13g2_xnor2_1 _14698_ (.Y(_06309_),
    .A(_06305_),
    .B(_06308_));
 sg13g2_nor2_1 _14699_ (.A(net2407),
    .B(_06304_),
    .Y(_06310_));
 sg13g2_a21oi_1 _14700_ (.A1(net2407),
    .A2(_06309_),
    .Y(_06311_),
    .B1(_06310_));
 sg13g2_a22oi_1 _14701_ (.Y(_06312_),
    .B1(net2062),
    .B2(\addr[6] ),
    .A2(net1752),
    .A1(net3291));
 sg13g2_a22oi_1 _14702_ (.Y(_06313_),
    .B1(_06311_),
    .B2(net1733),
    .A2(net1747),
    .A1(net3561));
 sg13g2_o21ai_1 _14703_ (.B1(_06313_),
    .Y(_00636_),
    .A1(net1747),
    .A2(_06312_));
 sg13g2_xnor2_1 _14704_ (.Y(_06314_),
    .A(net2416),
    .B(_06303_));
 sg13g2_and2_1 _14705_ (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(_06315_));
 sg13g2_xor2_1 _14706_ (.B(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .A(\i_tinyqv.cpu.instr_data_start[7] ),
    .X(_06316_));
 sg13g2_o21ai_1 _14707_ (.B1(_06306_),
    .Y(_06317_),
    .A1(_06305_),
    .A2(_06307_));
 sg13g2_and2_1 _14708_ (.A(_06316_),
    .B(_06317_),
    .X(_06318_));
 sg13g2_xor2_1 _14709_ (.B(_06317_),
    .A(_06316_),
    .X(_06319_));
 sg13g2_nand2_1 _14710_ (.Y(_06320_),
    .A(net2407),
    .B(_06319_));
 sg13g2_o21ai_1 _14711_ (.B1(_06320_),
    .Y(_06321_),
    .A1(net2404),
    .A2(_06314_));
 sg13g2_nand2_1 _14712_ (.Y(_06322_),
    .A(net1733),
    .B(_06321_));
 sg13g2_a221oi_1 _14713_ (.B2(\addr[7] ),
    .C1(net1746),
    .B1(net2063),
    .A1(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .Y(_06323_),
    .A2(net1752));
 sg13g2_a22oi_1 _14714_ (.Y(_00637_),
    .B1(_06322_),
    .B2(_06323_),
    .A2(net1747),
    .A1(_01153_));
 sg13g2_a22oi_1 _14715_ (.Y(_06324_),
    .B1(net2060),
    .B2(\addr[8] ),
    .A2(net1750),
    .A1(net3149));
 sg13g2_a21oi_1 _14716_ (.A1(net2416),
    .A2(_06303_),
    .Y(_06325_),
    .B1(\i_tinyqv.cpu.instr_data_start[8] ));
 sg13g2_nand3_1 _14717_ (.B(net2416),
    .C(_06303_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .Y(_06326_));
 sg13g2_nand2b_1 _14718_ (.Y(_06327_),
    .B(_06326_),
    .A_N(_06325_));
 sg13g2_nand2_1 _14719_ (.Y(_06328_),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[8] ));
 sg13g2_xor2_1 _14720_ (.B(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .A(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(_06329_));
 sg13g2_o21ai_1 _14721_ (.B1(_06329_),
    .Y(_06330_),
    .A1(_06315_),
    .A2(_06318_));
 sg13g2_or3_1 _14722_ (.A(_06315_),
    .B(_06318_),
    .C(_06329_),
    .X(_06331_));
 sg13g2_and2_1 _14723_ (.A(_06330_),
    .B(_06331_),
    .X(_06332_));
 sg13g2_nand2_1 _14724_ (.Y(_06333_),
    .A(net2404),
    .B(_06332_));
 sg13g2_o21ai_1 _14725_ (.B1(_06333_),
    .Y(_06334_),
    .A1(net2404),
    .A2(_06327_));
 sg13g2_a22oi_1 _14726_ (.Y(_06335_),
    .B1(_06334_),
    .B2(net1732),
    .A2(net1742),
    .A1(net3599));
 sg13g2_o21ai_1 _14727_ (.B1(_06335_),
    .Y(_00638_),
    .A1(net1743),
    .A2(_06324_));
 sg13g2_and2_1 _14728_ (.A(_00980_),
    .B(_06326_),
    .X(_06336_));
 sg13g2_nor2_2 _14729_ (.A(_00980_),
    .B(_06326_),
    .Y(_06337_));
 sg13g2_xnor2_1 _14730_ (.Y(_06338_),
    .A(\i_tinyqv.cpu.instr_data_start[9] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[9] ));
 sg13g2_a21oi_1 _14731_ (.A1(_06328_),
    .A2(_06330_),
    .Y(_06339_),
    .B1(_06338_));
 sg13g2_nand3_1 _14732_ (.B(_06330_),
    .C(_06338_),
    .A(_06328_),
    .Y(_06340_));
 sg13g2_nor2b_1 _14733_ (.A(_06339_),
    .B_N(_06340_),
    .Y(_06341_));
 sg13g2_nor3_1 _14734_ (.A(net2404),
    .B(_06336_),
    .C(_06337_),
    .Y(_06342_));
 sg13g2_a21oi_1 _14735_ (.A1(net2404),
    .A2(_06341_),
    .Y(_06343_),
    .B1(_06342_));
 sg13g2_a22oi_1 _14736_ (.Y(_06344_),
    .B1(net2062),
    .B2(\addr[9] ),
    .A2(net1752),
    .A1(net3164));
 sg13g2_o21ai_1 _14737_ (.B1(_06344_),
    .Y(_06345_),
    .A1(_05285_),
    .A2(_06343_));
 sg13g2_mux2_1 _14738_ (.A0(_06345_),
    .A1(net3208),
    .S(net1742),
    .X(_00639_));
 sg13g2_a22oi_1 _14739_ (.Y(_06346_),
    .B1(net2062),
    .B2(net3376),
    .A2(net1752),
    .A1(net3561));
 sg13g2_xnor2_1 _14740_ (.Y(_06347_),
    .A(net2415),
    .B(_06337_));
 sg13g2_a21o_1 _14741_ (.A2(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .A1(\i_tinyqv.cpu.instr_data_start[9] ),
    .B1(_06339_),
    .X(_06348_));
 sg13g2_xnor2_1 _14742_ (.Y(_06349_),
    .A(\i_tinyqv.cpu.instr_data_start[10] ),
    .B(\i_tinyqv.cpu.i_core.imm_lo[10] ));
 sg13g2_xnor2_1 _14743_ (.Y(_06350_),
    .A(_06348_),
    .B(_06349_));
 sg13g2_nand2_1 _14744_ (.Y(_06351_),
    .A(net2400),
    .B(_06350_));
 sg13g2_o21ai_1 _14745_ (.B1(_06351_),
    .Y(_06352_),
    .A1(net2401),
    .A2(_06347_));
 sg13g2_a22oi_1 _14746_ (.Y(_06353_),
    .B1(_06352_),
    .B2(net1732),
    .A2(net1744),
    .A1(net3604));
 sg13g2_o21ai_1 _14747_ (.B1(_06353_),
    .Y(_00640_),
    .A1(net1744),
    .A2(_06346_));
 sg13g2_a22oi_1 _14748_ (.Y(_06354_),
    .B1(net2061),
    .B2(\addr[11] ),
    .A2(net1750),
    .A1(net3174));
 sg13g2_a21oi_1 _14749_ (.A1(net2415),
    .A2(_06337_),
    .Y(_06355_),
    .B1(\i_tinyqv.cpu.instr_data_start[11] ));
 sg13g2_nand3_1 _14750_ (.B(net2415),
    .C(_06337_),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .Y(_06356_));
 sg13g2_nand2b_1 _14751_ (.Y(_06357_),
    .B(_06356_),
    .A_N(_06355_));
 sg13g2_xor2_1 _14752_ (.B(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .A(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(_06358_));
 sg13g2_a21o_1 _14753_ (.A2(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .A1(\i_tinyqv.cpu.instr_data_start[10] ),
    .B1(_06348_),
    .X(_06359_));
 sg13g2_o21ai_1 _14754_ (.B1(_06359_),
    .Y(_06360_),
    .A1(\i_tinyqv.cpu.instr_data_start[10] ),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[10] ));
 sg13g2_nor2b_1 _14755_ (.A(_06360_),
    .B_N(_06358_),
    .Y(_06361_));
 sg13g2_xnor2_1 _14756_ (.Y(_06362_),
    .A(_06358_),
    .B(_06360_));
 sg13g2_nand2_1 _14757_ (.Y(_06363_),
    .A(net2400),
    .B(_06362_));
 sg13g2_o21ai_1 _14758_ (.B1(_06363_),
    .Y(_06364_),
    .A1(net2400),
    .A2(_06357_));
 sg13g2_a22oi_1 _14759_ (.Y(_06365_),
    .B1(_06364_),
    .B2(net1732),
    .A2(net1744),
    .A1(net3656));
 sg13g2_o21ai_1 _14760_ (.B1(_06365_),
    .Y(_00641_),
    .A1(net1742),
    .A2(_06354_));
 sg13g2_a22oi_1 _14761_ (.Y(_06366_),
    .B1(net2060),
    .B2(net2991),
    .A2(net1749),
    .A1(net3599));
 sg13g2_nor2_1 _14762_ (.A(_00979_),
    .B(_06356_),
    .Y(_06367_));
 sg13g2_xnor2_1 _14763_ (.Y(_06368_),
    .A(_00979_),
    .B(_06356_));
 sg13g2_a21oi_1 _14764_ (.A1(\i_tinyqv.cpu.instr_data_start[11] ),
    .A2(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .Y(_06369_),
    .B1(_06361_));
 sg13g2_xor2_1 _14765_ (.B(\i_tinyqv.cpu.imm[12] ),
    .A(\i_tinyqv.cpu.instr_data_start[12] ),
    .X(_06370_));
 sg13g2_xnor2_1 _14766_ (.Y(_06371_),
    .A(_06369_),
    .B(_06370_));
 sg13g2_nand2_1 _14767_ (.Y(_06372_),
    .A(net2400),
    .B(_06371_));
 sg13g2_o21ai_1 _14768_ (.B1(_06372_),
    .Y(_06373_),
    .A1(net2400),
    .A2(_06368_));
 sg13g2_a22oi_1 _14769_ (.Y(_06374_),
    .B1(_06373_),
    .B2(net1732),
    .A2(net1742),
    .A1(net3603));
 sg13g2_o21ai_1 _14770_ (.B1(_06374_),
    .Y(_00642_),
    .A1(net1742),
    .A2(_06366_));
 sg13g2_xnor2_1 _14771_ (.Y(_06375_),
    .A(net2414),
    .B(_06367_));
 sg13g2_xor2_1 _14772_ (.B(\i_tinyqv.cpu.imm[13] ),
    .A(\i_tinyqv.cpu.instr_data_start[13] ),
    .X(_06376_));
 sg13g2_o21ai_1 _14773_ (.B1(_06369_),
    .Y(_06377_),
    .A1(_00979_),
    .A2(_01073_));
 sg13g2_o21ai_1 _14774_ (.B1(_06377_),
    .Y(_06378_),
    .A1(\i_tinyqv.cpu.instr_data_start[12] ),
    .A2(\i_tinyqv.cpu.imm[12] ));
 sg13g2_nor2b_1 _14775_ (.A(_06378_),
    .B_N(_06376_),
    .Y(_06379_));
 sg13g2_xnor2_1 _14776_ (.Y(_06380_),
    .A(_06376_),
    .B(_06378_));
 sg13g2_nand2_1 _14777_ (.Y(_06381_),
    .A(net2400),
    .B(_06380_));
 sg13g2_o21ai_1 _14778_ (.B1(_06381_),
    .Y(_06382_),
    .A1(net2400),
    .A2(_06375_));
 sg13g2_nand2_1 _14779_ (.Y(_06383_),
    .A(net1732),
    .B(_06382_));
 sg13g2_a221oi_1 _14780_ (.B2(\addr[13] ),
    .C1(net1743),
    .B1(net2060),
    .A1(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .Y(_06384_),
    .A2(net1749));
 sg13g2_a22oi_1 _14781_ (.Y(_00643_),
    .B1(_06383_),
    .B2(_06384_),
    .A2(net1742),
    .A1(_01154_));
 sg13g2_a22oi_1 _14782_ (.Y(_06385_),
    .B1(net2060),
    .B2(net3172),
    .A2(net1749),
    .A1(\i_tinyqv.mem.q_ctrl.addr[10] ));
 sg13g2_a21oi_1 _14783_ (.A1(net2414),
    .A2(_06367_),
    .Y(_06386_),
    .B1(net2413));
 sg13g2_nand3_1 _14784_ (.B(net2414),
    .C(_06367_),
    .A(net2413),
    .Y(_06387_));
 sg13g2_nand2b_1 _14785_ (.Y(_06388_),
    .B(_06387_),
    .A_N(_06386_));
 sg13g2_a21oi_1 _14786_ (.A1(net2414),
    .A2(\i_tinyqv.cpu.imm[13] ),
    .Y(_06389_),
    .B1(_06379_));
 sg13g2_nor2_1 _14787_ (.A(net2413),
    .B(\i_tinyqv.cpu.imm[14] ),
    .Y(_06390_));
 sg13g2_xor2_1 _14788_ (.B(\i_tinyqv.cpu.imm[14] ),
    .A(net2413),
    .X(_06391_));
 sg13g2_xnor2_1 _14789_ (.Y(_06392_),
    .A(_06389_),
    .B(_06391_));
 sg13g2_nand2_1 _14790_ (.Y(_06393_),
    .A(net2401),
    .B(_06392_));
 sg13g2_o21ai_1 _14791_ (.B1(_06393_),
    .Y(_06394_),
    .A1(net2401),
    .A2(_06388_));
 sg13g2_a22oi_1 _14792_ (.Y(_06395_),
    .B1(_06394_),
    .B2(net1732),
    .A2(net1744),
    .A1(net3523));
 sg13g2_o21ai_1 _14793_ (.B1(_06395_),
    .Y(_00644_),
    .A1(net1742),
    .A2(_06385_));
 sg13g2_nor2_2 _14794_ (.A(_00978_),
    .B(_06387_),
    .Y(_06396_));
 sg13g2_xnor2_1 _14795_ (.Y(_06397_),
    .A(_00978_),
    .B(_06387_));
 sg13g2_xor2_1 _14796_ (.B(\i_tinyqv.cpu.imm[15] ),
    .A(\i_tinyqv.cpu.instr_data_start[15] ),
    .X(_06398_));
 sg13g2_nor2_1 _14797_ (.A(_06389_),
    .B(_06390_),
    .Y(_06399_));
 sg13g2_a21oi_1 _14798_ (.A1(net2413),
    .A2(\i_tinyqv.cpu.imm[14] ),
    .Y(_06400_),
    .B1(_06399_));
 sg13g2_nand2b_1 _14799_ (.Y(_06401_),
    .B(_06398_),
    .A_N(_06400_));
 sg13g2_xnor2_1 _14800_ (.Y(_06402_),
    .A(_06398_),
    .B(_06400_));
 sg13g2_nand2_1 _14801_ (.Y(_06403_),
    .A(net2400),
    .B(_06402_));
 sg13g2_o21ai_1 _14802_ (.B1(_06403_),
    .Y(_06404_),
    .A1(net2401),
    .A2(_06397_));
 sg13g2_a22oi_1 _14803_ (.Y(_06405_),
    .B1(net2060),
    .B2(net3237),
    .A2(net1749),
    .A1(net3656));
 sg13g2_a22oi_1 _14804_ (.Y(_06406_),
    .B1(_06404_),
    .B2(net1732),
    .A2(net1744),
    .A1(net3778));
 sg13g2_o21ai_1 _14805_ (.B1(_06406_),
    .Y(_00645_),
    .A1(net1742),
    .A2(_06405_));
 sg13g2_a22oi_1 _14806_ (.Y(_06407_),
    .B1(net2060),
    .B2(net3095),
    .A2(net1749),
    .A1(\i_tinyqv.mem.q_ctrl.addr[12] ));
 sg13g2_xor2_1 _14807_ (.B(_06396_),
    .A(net2412),
    .X(_06408_));
 sg13g2_nor2_1 _14808_ (.A(net2402),
    .B(_06408_),
    .Y(_06409_));
 sg13g2_o21ai_1 _14809_ (.B1(_06401_),
    .Y(_06410_),
    .A1(_00978_),
    .A2(_01068_));
 sg13g2_xor2_1 _14810_ (.B(\i_tinyqv.cpu.imm[16] ),
    .A(\i_tinyqv.cpu.instr_data_start[16] ),
    .X(_06411_));
 sg13g2_xnor2_1 _14811_ (.Y(_06412_),
    .A(_06410_),
    .B(_06411_));
 sg13g2_a21oi_1 _14812_ (.A1(net2402),
    .A2(_06412_),
    .Y(_06413_),
    .B1(_06409_));
 sg13g2_a22oi_1 _14813_ (.Y(_06414_),
    .B1(_06413_),
    .B2(net1732),
    .A2(net1745),
    .A1(net3536));
 sg13g2_o21ai_1 _14814_ (.B1(_06414_),
    .Y(_00646_),
    .A1(net1744),
    .A2(_06407_));
 sg13g2_a21o_1 _14815_ (.A2(_06396_),
    .A1(net2412),
    .B1(net2411),
    .X(_06415_));
 sg13g2_nand3_1 _14816_ (.B(net2412),
    .C(_06396_),
    .A(net2411),
    .Y(_06416_));
 sg13g2_a21oi_1 _14817_ (.A1(_06415_),
    .A2(_06416_),
    .Y(_06417_),
    .B1(net2403));
 sg13g2_nand2_1 _14818_ (.Y(_06418_),
    .A(net2411),
    .B(\i_tinyqv.cpu.imm[17] ));
 sg13g2_nor2_1 _14819_ (.A(net2411),
    .B(\i_tinyqv.cpu.imm[17] ),
    .Y(_06419_));
 sg13g2_xor2_1 _14820_ (.B(\i_tinyqv.cpu.imm[17] ),
    .A(\i_tinyqv.cpu.instr_data_start[17] ),
    .X(_06420_));
 sg13g2_a21o_1 _14821_ (.A2(\i_tinyqv.cpu.imm[16] ),
    .A1(\i_tinyqv.cpu.instr_data_start[16] ),
    .B1(_06410_),
    .X(_06421_));
 sg13g2_o21ai_1 _14822_ (.B1(_06421_),
    .Y(_06422_),
    .A1(net2412),
    .A2(\i_tinyqv.cpu.imm[16] ));
 sg13g2_xnor2_1 _14823_ (.Y(_06423_),
    .A(_06420_),
    .B(_06422_));
 sg13g2_nor2b_1 _14824_ (.A(_06423_),
    .B_N(net2403),
    .Y(_06424_));
 sg13g2_or3_1 _14825_ (.A(_05285_),
    .B(_06417_),
    .C(_06424_),
    .X(_06425_));
 sg13g2_a221oi_1 _14826_ (.B2(\addr[17] ),
    .C1(net1743),
    .B1(net2060),
    .A1(net2809),
    .Y(_06426_),
    .A2(net1749));
 sg13g2_a22oi_1 _14827_ (.Y(_00647_),
    .B1(_06425_),
    .B2(_06426_),
    .A2(net1743),
    .A1(_01155_));
 sg13g2_nor2_1 _14828_ (.A(_00977_),
    .B(_06416_),
    .Y(_06427_));
 sg13g2_xnor2_1 _14829_ (.Y(_06428_),
    .A(\i_tinyqv.cpu.instr_data_start[18] ),
    .B(_06416_));
 sg13g2_nor2_1 _14830_ (.A(net2403),
    .B(_06428_),
    .Y(_06429_));
 sg13g2_o21ai_1 _14831_ (.B1(_06418_),
    .Y(_06430_),
    .A1(_06419_),
    .A2(_06422_));
 sg13g2_xor2_1 _14832_ (.B(\i_tinyqv.cpu.imm[18] ),
    .A(\i_tinyqv.cpu.instr_data_start[18] ),
    .X(_06431_));
 sg13g2_xnor2_1 _14833_ (.Y(_06432_),
    .A(_06430_),
    .B(_06431_));
 sg13g2_a21oi_1 _14834_ (.A1(net2403),
    .A2(_06432_),
    .Y(_06433_),
    .B1(_06429_));
 sg13g2_a22oi_1 _14835_ (.Y(_06434_),
    .B1(net2060),
    .B2(net3168),
    .A2(net1749),
    .A1(net3523));
 sg13g2_a22oi_1 _14836_ (.Y(_06435_),
    .B1(_06433_),
    .B2(net1733),
    .A2(net1745),
    .A1(net3655));
 sg13g2_o21ai_1 _14837_ (.B1(_06435_),
    .Y(_00648_),
    .A1(net1748),
    .A2(_06434_));
 sg13g2_xor2_1 _14838_ (.B(_06427_),
    .A(net2410),
    .X(_06436_));
 sg13g2_nor2_1 _14839_ (.A(net2403),
    .B(_06436_),
    .Y(_06437_));
 sg13g2_nand2_1 _14840_ (.Y(_06438_),
    .A(net2410),
    .B(\i_tinyqv.cpu.imm[19] ));
 sg13g2_xnor2_1 _14841_ (.Y(_06439_),
    .A(net2410),
    .B(\i_tinyqv.cpu.imm[19] ));
 sg13g2_a21o_1 _14842_ (.A2(\i_tinyqv.cpu.imm[18] ),
    .A1(\i_tinyqv.cpu.instr_data_start[18] ),
    .B1(_06430_),
    .X(_06440_));
 sg13g2_o21ai_1 _14843_ (.B1(_06440_),
    .Y(_06441_),
    .A1(\i_tinyqv.cpu.instr_data_start[18] ),
    .A2(\i_tinyqv.cpu.imm[18] ));
 sg13g2_xnor2_1 _14844_ (.Y(_06442_),
    .A(_06439_),
    .B(_06441_));
 sg13g2_a21oi_1 _14845_ (.A1(net2403),
    .A2(_06442_),
    .Y(_06443_),
    .B1(_06437_));
 sg13g2_a22oi_1 _14846_ (.Y(_06444_),
    .B1(net2061),
    .B2(net3197),
    .A2(net1750),
    .A1(\i_tinyqv.mem.q_ctrl.addr[15] ));
 sg13g2_a22oi_1 _14847_ (.Y(_06445_),
    .B1(_06443_),
    .B2(net1733),
    .A2(net1746),
    .A1(net3543));
 sg13g2_o21ai_1 _14848_ (.B1(_06445_),
    .Y(_00649_),
    .A1(net1745),
    .A2(_06444_));
 sg13g2_o21ai_1 _14849_ (.B1(_06438_),
    .Y(_06446_),
    .A1(_06439_),
    .A2(_06441_));
 sg13g2_nor2_1 _14850_ (.A(net2409),
    .B(\i_tinyqv.cpu.imm[20] ),
    .Y(_06447_));
 sg13g2_xor2_1 _14851_ (.B(\i_tinyqv.cpu.imm[20] ),
    .A(net2409),
    .X(_06448_));
 sg13g2_xnor2_1 _14852_ (.Y(_06449_),
    .A(_06446_),
    .B(_06448_));
 sg13g2_nand3_1 _14853_ (.B(\i_tinyqv.cpu.instr_data_start[19] ),
    .C(_06427_),
    .A(net2409),
    .Y(_06450_));
 sg13g2_a21o_1 _14854_ (.A2(_06427_),
    .A1(\i_tinyqv.cpu.instr_data_start[19] ),
    .B1(net2409),
    .X(_06451_));
 sg13g2_a21oi_1 _14855_ (.A1(_06450_),
    .A2(_06451_),
    .Y(_06452_),
    .B1(net2405));
 sg13g2_a21oi_1 _14856_ (.A1(net2405),
    .A2(_06449_),
    .Y(_06453_),
    .B1(_06452_));
 sg13g2_a22oi_1 _14857_ (.Y(_06454_),
    .B1(net2061),
    .B2(net3309),
    .A2(net1751),
    .A1(net3536));
 sg13g2_a22oi_1 _14858_ (.Y(_06455_),
    .B1(_06453_),
    .B2(net1733),
    .A2(net1746),
    .A1(net3742));
 sg13g2_o21ai_1 _14859_ (.B1(_06455_),
    .Y(_00650_),
    .A1(net1745),
    .A2(_06454_));
 sg13g2_xnor2_1 _14860_ (.Y(_06456_),
    .A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(\i_tinyqv.cpu.imm[21] ));
 sg13g2_a21oi_1 _14861_ (.A1(\i_tinyqv.cpu.instr_data_start[20] ),
    .A2(\i_tinyqv.cpu.imm[20] ),
    .Y(_06457_),
    .B1(_06446_));
 sg13g2_or3_1 _14862_ (.A(_06447_),
    .B(_06456_),
    .C(_06457_),
    .X(_06458_));
 sg13g2_o21ai_1 _14863_ (.B1(_06456_),
    .Y(_06459_),
    .A1(_06447_),
    .A2(_06457_));
 sg13g2_nand2_1 _14864_ (.Y(_06460_),
    .A(_06458_),
    .B(_06459_));
 sg13g2_nor2_1 _14865_ (.A(_00976_),
    .B(_06450_),
    .Y(_06461_));
 sg13g2_xnor2_1 _14866_ (.Y(_06462_),
    .A(\i_tinyqv.cpu.instr_data_start[21] ),
    .B(_06450_));
 sg13g2_nor2_1 _14867_ (.A(net2405),
    .B(_06462_),
    .Y(_06463_));
 sg13g2_a21oi_1 _14868_ (.A1(net2404),
    .A2(_06460_),
    .Y(_06464_),
    .B1(_06463_));
 sg13g2_a22oi_1 _14869_ (.Y(_06465_),
    .B1(_06464_),
    .B2(net1733),
    .A2(net1745),
    .A1(net3685));
 sg13g2_a22oi_1 _14870_ (.Y(_06466_),
    .B1(net2061),
    .B2(net3154),
    .A2(net1749),
    .A1(net2916));
 sg13g2_o21ai_1 _14871_ (.B1(_06465_),
    .Y(_00651_),
    .A1(net1745),
    .A2(_06466_));
 sg13g2_a221oi_1 _14872_ (.B2(net3043),
    .C1(net1745),
    .B1(net2061),
    .A1(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .Y(_06467_),
    .A2(net1751));
 sg13g2_nor2b_1 _14873_ (.A(net3303),
    .B_N(net1746),
    .Y(_06468_));
 sg13g2_o21ai_1 _14874_ (.B1(_06458_),
    .Y(_06469_),
    .A1(_00976_),
    .A2(_01072_));
 sg13g2_xor2_1 _14875_ (.B(\i_tinyqv.cpu.imm[22] ),
    .A(\i_tinyqv.cpu.instr_data_start[22] ),
    .X(_06470_));
 sg13g2_xnor2_1 _14876_ (.Y(_06471_),
    .A(_06469_),
    .B(_06470_));
 sg13g2_nand2_1 _14877_ (.Y(_06472_),
    .A(\i_tinyqv.cpu.instr_data_start[22] ),
    .B(_06461_));
 sg13g2_xnor2_1 _14878_ (.Y(_06473_),
    .A(_00975_),
    .B(_06461_));
 sg13g2_a21oi_1 _14879_ (.A1(net2405),
    .A2(_06471_),
    .Y(_06474_),
    .B1(_05285_));
 sg13g2_o21ai_1 _14880_ (.B1(_06474_),
    .Y(_06475_),
    .A1(net2404),
    .A2(_06473_));
 sg13g2_o21ai_1 _14881_ (.B1(_06475_),
    .Y(_00652_),
    .A1(_06467_),
    .A2(_06468_));
 sg13g2_a21o_1 _14882_ (.A2(\i_tinyqv.cpu.imm[22] ),
    .A1(\i_tinyqv.cpu.instr_data_start[22] ),
    .B1(_06469_),
    .X(_06476_));
 sg13g2_o21ai_1 _14883_ (.B1(_06476_),
    .Y(_06477_),
    .A1(\i_tinyqv.cpu.instr_data_start[22] ),
    .A2(\i_tinyqv.cpu.imm[22] ));
 sg13g2_xnor2_1 _14884_ (.Y(_06478_),
    .A(\i_tinyqv.cpu.instr_data_start[23] ),
    .B(\i_tinyqv.cpu.imm[23] ));
 sg13g2_xnor2_1 _14885_ (.Y(_06479_),
    .A(_06477_),
    .B(_06478_));
 sg13g2_a21oi_1 _14886_ (.A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(_06472_),
    .Y(_06480_),
    .B1(net2405));
 sg13g2_o21ai_1 _14887_ (.B1(_06480_),
    .Y(_06481_),
    .A1(\i_tinyqv.cpu.instr_data_start[23] ),
    .A2(_06472_));
 sg13g2_a21oi_1 _14888_ (.A1(net2404),
    .A2(_06479_),
    .Y(_06482_),
    .B1(net1753));
 sg13g2_a22oi_1 _14889_ (.Y(_06483_),
    .B1(_06481_),
    .B2(_06482_),
    .A2(net1753),
    .A1(\addr[23] ));
 sg13g2_a22oi_1 _14890_ (.Y(_06484_),
    .B1(net1746),
    .B2(net3318),
    .A2(_02810_),
    .A1(\i_tinyqv.mem.q_ctrl.addr[19] ));
 sg13g2_o21ai_1 _14891_ (.B1(net3319),
    .Y(_00653_),
    .A1(net1751),
    .A2(_06483_));
 sg13g2_nor2_1 _14892_ (.A(net2346),
    .B(net1739),
    .Y(_06485_));
 sg13g2_a22oi_1 _14893_ (.Y(_00654_),
    .B1(_06485_),
    .B2(_01088_),
    .A2(net1739),
    .A1(_01117_));
 sg13g2_a22oi_1 _14894_ (.Y(_00655_),
    .B1(_06485_),
    .B2(_01092_),
    .A2(net1739),
    .A1(_01123_));
 sg13g2_nor3_1 _14895_ (.A(_01076_),
    .B(\i_tinyqv.cpu.instr_write_offset[1] ),
    .C(_02641_),
    .Y(_06486_));
 sg13g2_nand2b_1 _14896_ (.Y(_06487_),
    .B(net2497),
    .A_N(net1735));
 sg13g2_nor2_1 _14897_ (.A(net3223),
    .B(_06487_),
    .Y(_06488_));
 sg13g2_a21oi_1 _14898_ (.A1(_01117_),
    .A2(net1735),
    .Y(_00656_),
    .B1(_06488_));
 sg13g2_nor2_1 _14899_ (.A(net3113),
    .B(_06487_),
    .Y(_06489_));
 sg13g2_a21oi_1 _14900_ (.A1(_01123_),
    .A2(net1735),
    .Y(_00657_),
    .B1(_06489_));
 sg13g2_xnor2_1 _14901_ (.Y(_06490_),
    .A(net3948),
    .B(_02837_));
 sg13g2_o21ai_1 _14902_ (.B1(net2495),
    .Y(_06491_),
    .A1(_02816_),
    .A2(net1992));
 sg13g2_a21oi_1 _14903_ (.A1(net1992),
    .A2(net3949),
    .Y(_00658_),
    .B1(_06491_));
 sg13g2_xnor2_1 _14904_ (.Y(_06492_),
    .A(net3760),
    .B(_02838_));
 sg13g2_o21ai_1 _14905_ (.B1(net2495),
    .Y(_06493_),
    .A1(_02817_),
    .A2(net1992));
 sg13g2_a21oi_1 _14906_ (.A1(net1992),
    .A2(_06492_),
    .Y(_00659_),
    .B1(_06493_));
 sg13g2_nand3_1 _14907_ (.B(net3760),
    .C(_02838_),
    .A(net4142),
    .Y(_06494_));
 sg13g2_xor2_1 _14908_ (.B(_02839_),
    .A(net4142),
    .X(_06495_));
 sg13g2_o21ai_1 _14909_ (.B1(net2495),
    .Y(_06496_),
    .A1(_02821_),
    .A2(net1992));
 sg13g2_a21oi_1 _14910_ (.A1(net1992),
    .A2(_06495_),
    .Y(_00660_),
    .B1(_06496_));
 sg13g2_xor2_1 _14911_ (.B(_06494_),
    .A(net4038),
    .X(_06497_));
 sg13g2_o21ai_1 _14912_ (.B1(net2495),
    .Y(_06498_),
    .A1(_02823_),
    .A2(net1992));
 sg13g2_a21oi_2 _14913_ (.B1(_06498_),
    .Y(_00661_),
    .A2(_06497_),
    .A1(net1992));
 sg13g2_nand2_1 _14914_ (.Y(_06499_),
    .A(_01434_),
    .B(_01435_));
 sg13g2_nand2_1 _14915_ (.Y(_06500_),
    .A(\i_tinyqv.mem.q_ctrl.data_req ),
    .B(_06499_));
 sg13g2_o21ai_1 _14916_ (.B1(_01906_),
    .Y(_06501_),
    .A1(_01436_),
    .A2(_06500_));
 sg13g2_a21oi_1 _14917_ (.A1(net2273),
    .A2(_06501_),
    .Y(_06502_),
    .B1(net2957));
 sg13g2_nand3b_1 _14918_ (.B(_01916_),
    .C(net2957),
    .Y(_06503_),
    .A_N(_02589_));
 sg13g2_o21ai_1 _14919_ (.B1(net3646),
    .Y(_06504_),
    .A1(_06501_),
    .A2(_06503_));
 sg13g2_a21oi_1 _14920_ (.A1(net2273),
    .A2(_06504_),
    .Y(_00662_),
    .B1(net2958));
 sg13g2_nor2_1 _14921_ (.A(net3945),
    .B(_02803_),
    .Y(_06505_));
 sg13g2_a21oi_1 _14922_ (.A1(net3800),
    .A2(\i_tinyqv.cpu.data_write_n[1] ),
    .Y(_06506_),
    .B1(_02804_));
 sg13g2_a221oi_1 _14923_ (.B2(net3798),
    .C1(_02804_),
    .B1(\i_tinyqv.cpu.data_write_n[0] ),
    .A1(net3800),
    .Y(_06507_),
    .A2(\i_tinyqv.cpu.data_write_n[1] ));
 sg13g2_o21ai_1 _14924_ (.B1(net2273),
    .Y(_00663_),
    .A1(net3946),
    .A2(_06507_));
 sg13g2_nor2_1 _14925_ (.A(net3882),
    .B(_02803_),
    .Y(_06508_));
 sg13g2_o21ai_1 _14926_ (.B1(net2273),
    .Y(_00664_),
    .A1(_06506_),
    .A2(net3883));
 sg13g2_o21ai_1 _14927_ (.B1(debug_data_continue),
    .Y(_06509_),
    .A1(net3646),
    .A2(_02803_));
 sg13g2_a21oi_1 _14928_ (.A1(_06504_),
    .A2(_06509_),
    .Y(_00665_),
    .B1(net2246));
 sg13g2_a21oi_1 _14929_ (.A1(_01437_),
    .A2(net1753),
    .Y(_06510_),
    .B1(_02592_));
 sg13g2_nor2_1 _14930_ (.A(net4028),
    .B(_06510_),
    .Y(_06511_));
 sg13g2_nand2_1 _14931_ (.Y(_06512_),
    .A(net2273),
    .B(net1752));
 sg13g2_nor2_1 _14932_ (.A(_00985_),
    .B(_02592_),
    .Y(_06513_));
 sg13g2_nor3_1 _14933_ (.A(_06511_),
    .B(_06512_),
    .C(_06513_),
    .Y(_00666_));
 sg13g2_nand2_1 _14934_ (.Y(_06514_),
    .A(net4030),
    .B(_00985_));
 sg13g2_nand3_1 _14935_ (.B(_02572_),
    .C(_02806_),
    .A(_02045_),
    .Y(_06515_));
 sg13g2_nand2_1 _14936_ (.Y(_06516_),
    .A(_06514_),
    .B(_06515_));
 sg13g2_a22oi_1 _14937_ (.Y(_06517_),
    .B1(_06510_),
    .B2(_06516_),
    .A2(_02592_),
    .A1(net4030));
 sg13g2_nor2_1 _14938_ (.A(_06512_),
    .B(net4031),
    .Y(_00667_));
 sg13g2_a21oi_1 _14939_ (.A1(\i_tinyqv.mem.data_stall ),
    .A2(_01909_),
    .Y(_06518_),
    .B1(net2435));
 sg13g2_nor2b_2 _14940_ (.A(_01915_),
    .B_N(_06518_),
    .Y(_06519_));
 sg13g2_nor2_1 _14941_ (.A(net2335),
    .B(_01916_),
    .Y(_06520_));
 sg13g2_or2_1 _14942_ (.X(_06521_),
    .B(_06520_),
    .A(net2006));
 sg13g2_nand2b_1 _14943_ (.Y(_06522_),
    .B(net2429),
    .A_N(net2423));
 sg13g2_o21ai_1 _14944_ (.B1(_06522_),
    .Y(_06523_),
    .A1(\data_to_write[0] ),
    .A2(net2429));
 sg13g2_nand2_1 _14945_ (.Y(_06524_),
    .A(net3245),
    .B(net1970));
 sg13g2_o21ai_1 _14946_ (.B1(_06524_),
    .Y(_00668_),
    .A1(net1970),
    .A2(_06523_));
 sg13g2_nand2_1 _14947_ (.Y(_06525_),
    .A(net2430),
    .B(_01124_));
 sg13g2_o21ai_1 _14948_ (.B1(_06525_),
    .Y(_06526_),
    .A1(net2398),
    .A2(net2433));
 sg13g2_nand2_1 _14949_ (.Y(_06527_),
    .A(net3554),
    .B(net1971));
 sg13g2_o21ai_1 _14950_ (.B1(_06527_),
    .Y(_00669_),
    .A1(net1971),
    .A2(_06526_));
 sg13g2_nand2_1 _14951_ (.Y(_06528_),
    .A(net2430),
    .B(net2330));
 sg13g2_o21ai_1 _14952_ (.B1(_06528_),
    .Y(_06529_),
    .A1(net2396),
    .A2(net2430));
 sg13g2_nand2_1 _14953_ (.Y(_06530_),
    .A(net3844),
    .B(net1971));
 sg13g2_o21ai_1 _14954_ (.B1(_06530_),
    .Y(_00670_),
    .A1(net1971),
    .A2(_06529_));
 sg13g2_nand2_1 _14955_ (.Y(_06531_),
    .A(net2435),
    .B(_01133_));
 sg13g2_o21ai_1 _14956_ (.B1(_06531_),
    .Y(_06532_),
    .A1(net2394),
    .A2(net2435));
 sg13g2_nand2_1 _14957_ (.Y(_06533_),
    .A(net3636),
    .B(net1970));
 sg13g2_o21ai_1 _14958_ (.B1(_06533_),
    .Y(_00671_),
    .A1(net1970),
    .A2(_06532_));
 sg13g2_nand2b_1 _14959_ (.Y(_06534_),
    .B(net2431),
    .A_N(net2420));
 sg13g2_o21ai_1 _14960_ (.B1(_06534_),
    .Y(_06535_),
    .A1(net2392),
    .A2(net2431));
 sg13g2_nand2_1 _14961_ (.Y(_06536_),
    .A(net3045),
    .B(net1971));
 sg13g2_o21ai_1 _14962_ (.B1(_06536_),
    .Y(_00672_),
    .A1(net1970),
    .A2(_06535_));
 sg13g2_nand2_2 _14963_ (.Y(_06537_),
    .A(net2434),
    .B(\i_tinyqv.cpu.instr_data_in[13] ));
 sg13g2_o21ai_1 _14964_ (.B1(_06537_),
    .Y(_06538_),
    .A1(_00969_),
    .A2(net2431));
 sg13g2_mux2_1 _14965_ (.A0(_06538_),
    .A1(net4086),
    .S(net1971),
    .X(_00673_));
 sg13g2_nand2_2 _14966_ (.Y(_06539_),
    .A(net2429),
    .B(net3996));
 sg13g2_o21ai_1 _14967_ (.B1(_06539_),
    .Y(_06540_),
    .A1(_00968_),
    .A2(net2430));
 sg13g2_mux2_1 _14968_ (.A0(_06540_),
    .A1(net4055),
    .S(net1970),
    .X(_00674_));
 sg13g2_nand2_2 _14969_ (.Y(_06541_),
    .A(net2434),
    .B(net2419));
 sg13g2_a21oi_1 _14970_ (.A1(\data_to_write[7] ),
    .A2(net2335),
    .Y(_06542_),
    .B1(net1970));
 sg13g2_a22oi_1 _14971_ (.Y(_00675_),
    .B1(_06541_),
    .B2(_06542_),
    .A2(net1970),
    .A1(_01134_));
 sg13g2_nor2_1 _14972_ (.A(net2335),
    .B(_02572_),
    .Y(_06543_));
 sg13g2_or2_1 _14973_ (.X(_06544_),
    .B(_06543_),
    .A(net2006));
 sg13g2_nand2_1 _14974_ (.Y(_06545_),
    .A(net2949),
    .B(net1969));
 sg13g2_a22oi_1 _14975_ (.Y(_06546_),
    .B1(net2423),
    .B2(_02573_),
    .A2(net2335),
    .A1(\data_to_write[8] ));
 sg13g2_o21ai_1 _14976_ (.B1(_06545_),
    .Y(_00676_),
    .A1(net2006),
    .A2(_06546_));
 sg13g2_nand2_1 _14977_ (.Y(_06547_),
    .A(net3018),
    .B(net1969));
 sg13g2_a22oi_1 _14978_ (.Y(_06548_),
    .B1(\i_tinyqv.cpu.instr_data_in[9] ),
    .B2(_02573_),
    .A2(net2335),
    .A1(\data_to_write[9] ));
 sg13g2_o21ai_1 _14979_ (.B1(_06547_),
    .Y(_00677_),
    .A1(net2006),
    .A2(_06548_));
 sg13g2_nand2_1 _14980_ (.Y(_06549_),
    .A(net2931),
    .B(net1969));
 sg13g2_a22oi_1 _14981_ (.Y(_06550_),
    .B1(\i_tinyqv.cpu.instr_data_in[10] ),
    .B2(_02573_),
    .A2(_01078_),
    .A1(\data_to_write[10] ));
 sg13g2_o21ai_1 _14982_ (.B1(_06549_),
    .Y(_00678_),
    .A1(net2006),
    .A2(_06550_));
 sg13g2_nand2_1 _14983_ (.Y(_06551_),
    .A(net2787),
    .B(net1969));
 sg13g2_a22oi_1 _14984_ (.Y(_06552_),
    .B1(\i_tinyqv.cpu.instr_data_in[11] ),
    .B2(_02573_),
    .A2(_01078_),
    .A1(\data_to_write[11] ));
 sg13g2_o21ai_1 _14985_ (.B1(_06551_),
    .Y(_00679_),
    .A1(net2006),
    .A2(_06552_));
 sg13g2_nand2_1 _14986_ (.Y(_06553_),
    .A(net2882),
    .B(net1969));
 sg13g2_a22oi_1 _14987_ (.Y(_06554_),
    .B1(net2420),
    .B2(_02573_),
    .A2(_01078_),
    .A1(\data_to_write[12] ));
 sg13g2_o21ai_1 _14988_ (.B1(_06553_),
    .Y(_00680_),
    .A1(_06519_),
    .A2(_06554_));
 sg13g2_o21ai_1 _14989_ (.B1(_06537_),
    .Y(_06555_),
    .A1(_00965_),
    .A2(net2434));
 sg13g2_nor2_1 _14990_ (.A(net1969),
    .B(_06555_),
    .Y(_06556_));
 sg13g2_a21oi_1 _14991_ (.A1(_01127_),
    .A2(net1969),
    .Y(_00681_),
    .B1(_06556_));
 sg13g2_o21ai_1 _14992_ (.B1(_06539_),
    .Y(_06557_),
    .A1(_00964_),
    .A2(net2430));
 sg13g2_mux2_1 _14993_ (.A0(_06557_),
    .A1(net3629),
    .S(net1969),
    .X(_00682_));
 sg13g2_o21ai_1 _14994_ (.B1(_06541_),
    .Y(_06558_),
    .A1(_00963_),
    .A2(net2429));
 sg13g2_mux2_1 _14995_ (.A0(_06558_),
    .A1(net3664),
    .S(_06544_),
    .X(_00683_));
 sg13g2_a21o_1 _14996_ (.A2(_06514_),
    .A1(net2435),
    .B1(net2006),
    .X(_06559_));
 sg13g2_o21ai_1 _14997_ (.B1(_06522_),
    .Y(_06560_),
    .A1(\data_to_write[16] ),
    .A2(net2429));
 sg13g2_nand2_1 _14998_ (.Y(_06561_),
    .A(net2851),
    .B(net1968));
 sg13g2_o21ai_1 _14999_ (.B1(_06561_),
    .Y(_00684_),
    .A1(net1968),
    .A2(_06560_));
 sg13g2_o21ai_1 _15000_ (.B1(_06525_),
    .Y(_06562_),
    .A1(\data_to_write[17] ),
    .A2(net2430));
 sg13g2_nand2_1 _15001_ (.Y(_06563_),
    .A(net2839),
    .B(net1967));
 sg13g2_o21ai_1 _15002_ (.B1(_06563_),
    .Y(_00685_),
    .A1(net1967),
    .A2(_06562_));
 sg13g2_o21ai_1 _15003_ (.B1(_06528_),
    .Y(_06564_),
    .A1(\data_to_write[18] ),
    .A2(net2430));
 sg13g2_nand2_1 _15004_ (.Y(_06565_),
    .A(net2867),
    .B(net1967));
 sg13g2_o21ai_1 _15005_ (.B1(_06565_),
    .Y(_00686_),
    .A1(net1967),
    .A2(_06564_));
 sg13g2_o21ai_1 _15006_ (.B1(_06531_),
    .Y(_06566_),
    .A1(\data_to_write[19] ),
    .A2(net2435));
 sg13g2_nand2_1 _15007_ (.Y(_06567_),
    .A(net2832),
    .B(net1968));
 sg13g2_o21ai_1 _15008_ (.B1(_06567_),
    .Y(_00687_),
    .A1(net1968),
    .A2(_06566_));
 sg13g2_o21ai_1 _15009_ (.B1(_06534_),
    .Y(_06568_),
    .A1(\data_to_write[20] ),
    .A2(net2431));
 sg13g2_nand2_1 _15010_ (.Y(_06569_),
    .A(net3009),
    .B(net1967));
 sg13g2_o21ai_1 _15011_ (.B1(_06569_),
    .Y(_00688_),
    .A1(net1968),
    .A2(_06568_));
 sg13g2_o21ai_1 _15012_ (.B1(_06537_),
    .Y(_06570_),
    .A1(_00958_),
    .A2(net2431));
 sg13g2_mux2_1 _15013_ (.A0(_06570_),
    .A1(net3613),
    .S(net1967),
    .X(_00689_));
 sg13g2_o21ai_1 _15014_ (.B1(_06539_),
    .Y(_06571_),
    .A1(_00957_),
    .A2(net2429));
 sg13g2_mux2_1 _15015_ (.A0(_06571_),
    .A1(net3593),
    .S(net1967),
    .X(_00690_));
 sg13g2_o21ai_1 _15016_ (.B1(_06541_),
    .Y(_06572_),
    .A1(_00956_),
    .A2(net2429));
 sg13g2_mux2_1 _15017_ (.A0(_06572_),
    .A1(net3493),
    .S(net1967),
    .X(_00691_));
 sg13g2_a21oi_1 _15018_ (.A1(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .A2(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .Y(_06573_),
    .B1(net2335));
 sg13g2_nor2_1 _15019_ (.A(net2006),
    .B(_06573_),
    .Y(_06574_));
 sg13g2_nor2_1 _15020_ (.A(_00955_),
    .B(net2431),
    .Y(_06575_));
 sg13g2_a21oi_1 _15021_ (.A1(net2432),
    .A2(net2422),
    .Y(_06576_),
    .B1(_06575_));
 sg13g2_nor2_1 _15022_ (.A(net3342),
    .B(net1965),
    .Y(_06577_));
 sg13g2_a21oi_1 _15023_ (.A1(net1965),
    .A2(_06576_),
    .Y(_00692_),
    .B1(_06577_));
 sg13g2_mux2_1 _15024_ (.A0(_00954_),
    .A1(_01124_),
    .S(net2432),
    .X(_06578_));
 sg13g2_nor2_1 _15025_ (.A(net3433),
    .B(net1965),
    .Y(_06579_));
 sg13g2_a21oi_1 _15026_ (.A1(net1965),
    .A2(_06578_),
    .Y(_00693_),
    .B1(_06579_));
 sg13g2_mux2_1 _15027_ (.A0(_00953_),
    .A1(net2330),
    .S(net2432),
    .X(_06580_));
 sg13g2_nor2_1 _15028_ (.A(net3425),
    .B(net1965),
    .Y(_06581_));
 sg13g2_a21oi_1 _15029_ (.A1(net1965),
    .A2(_06580_),
    .Y(_00694_),
    .B1(_06581_));
 sg13g2_mux2_1 _15030_ (.A0(_00952_),
    .A1(_01133_),
    .S(net2432),
    .X(_06582_));
 sg13g2_nor2_1 _15031_ (.A(net3454),
    .B(net1965),
    .Y(_06583_));
 sg13g2_a21oi_1 _15032_ (.A1(net1965),
    .A2(_06582_),
    .Y(_00695_),
    .B1(_06583_));
 sg13g2_nor2_1 _15033_ (.A(_00951_),
    .B(net2431),
    .Y(_06584_));
 sg13g2_a21oi_1 _15034_ (.A1(net2432),
    .A2(net2420),
    .Y(_06585_),
    .B1(_06584_));
 sg13g2_nor2_1 _15035_ (.A(net3321),
    .B(net1966),
    .Y(_06586_));
 sg13g2_a21oi_1 _15036_ (.A1(net1966),
    .A2(_06585_),
    .Y(_00696_),
    .B1(_06586_));
 sg13g2_o21ai_1 _15037_ (.B1(_06537_),
    .Y(_06587_),
    .A1(_00950_),
    .A2(net2431));
 sg13g2_mux2_1 _15038_ (.A0(net3611),
    .A1(_06587_),
    .S(net1966),
    .X(_00697_));
 sg13g2_o21ai_1 _15039_ (.B1(_06539_),
    .Y(_06588_),
    .A1(_00949_),
    .A2(net2430));
 sg13g2_mux2_1 _15040_ (.A0(net3659),
    .A1(_06588_),
    .S(net1966),
    .X(_00698_));
 sg13g2_o21ai_1 _15041_ (.B1(_06541_),
    .Y(_06589_),
    .A1(_00948_),
    .A2(net2429));
 sg13g2_mux2_1 _15042_ (.A0(net3385),
    .A1(_06589_),
    .S(net1966),
    .X(_00699_));
 sg13g2_and2_1 _15043_ (.A(net2273),
    .B(_02805_),
    .X(_00700_));
 sg13g2_nor2_1 _15044_ (.A(net2438),
    .B(_01911_),
    .Y(_06590_));
 sg13g2_o21ai_1 _15045_ (.B1(net2273),
    .Y(_06591_),
    .A1(_01912_),
    .A2(_02805_));
 sg13g2_nor3_1 _15046_ (.A(_02595_),
    .B(net4115),
    .C(_06591_),
    .Y(_00701_));
 sg13g2_nor2_1 _15047_ (.A(net2267),
    .B(net10),
    .Y(_06592_));
 sg13g2_a21oi_1 _15048_ (.A1(net2267),
    .A2(_01152_),
    .Y(_00702_),
    .B1(_06592_));
 sg13g2_mux2_1 _15049_ (.A0(net11),
    .A1(net3479),
    .S(net2266),
    .X(_00703_));
 sg13g2_nand2_2 _15050_ (.Y(_06593_),
    .A(net2425),
    .B(net2426));
 sg13g2_nand3_1 _15051_ (.B(net2426),
    .C(net2428),
    .A(net2425),
    .Y(_06594_));
 sg13g2_nand2_2 _15052_ (.Y(_06595_),
    .A(net2425),
    .B(net2428));
 sg13g2_a21oi_1 _15053_ (.A1(net2436),
    .A2(_06594_),
    .Y(_06596_),
    .B1(_06595_));
 sg13g2_nor2_1 _15054_ (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .Y(_06597_));
 sg13g2_mux2_1 _15055_ (.A0(net3753),
    .A1(_06597_),
    .S(_06596_),
    .X(_06598_));
 sg13g2_nor2_1 _15056_ (.A(net3814),
    .B(net3482),
    .Y(_06599_));
 sg13g2_nor3_2 _15057_ (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .B(net3814),
    .C(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .Y(_06600_));
 sg13g2_nand2b_1 _15058_ (.Y(_06601_),
    .B(_06599_),
    .A_N(net3239));
 sg13g2_nand2_1 _15059_ (.Y(_06602_),
    .A(net2436),
    .B(_02416_));
 sg13g2_nor4_1 _15060_ (.A(net1731),
    .B(_06598_),
    .C(_06601_),
    .D(_06602_),
    .Y(_00704_));
 sg13g2_nor2_2 _15061_ (.A(net2428),
    .B(_06593_),
    .Y(_06603_));
 sg13g2_or2_1 _15062_ (.X(_06604_),
    .B(_06593_),
    .A(net2428));
 sg13g2_and2_1 _15063_ (.A(_06598_),
    .B(_06600_),
    .X(_06605_));
 sg13g2_nand2_1 _15064_ (.Y(_06606_),
    .A(_06598_),
    .B(_06600_));
 sg13g2_nand2_1 _15065_ (.Y(_06607_),
    .A(_06595_),
    .B(_06605_));
 sg13g2_and2_1 _15066_ (.A(net2425),
    .B(_01910_),
    .X(_06608_));
 sg13g2_nand2_1 _15067_ (.Y(_06609_),
    .A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .B(_06608_));
 sg13g2_o21ai_1 _15068_ (.B1(_06609_),
    .Y(_06610_),
    .A1(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .A2(_06608_));
 sg13g2_o21ai_1 _15069_ (.B1(_06604_),
    .Y(_06611_),
    .A1(_06607_),
    .A2(_06610_));
 sg13g2_nand2b_2 _15070_ (.Y(_06612_),
    .B(_02586_),
    .A_N(\i_tinyqv.mem.data_stall ));
 sg13g2_nand2b_1 _15071_ (.Y(_06613_),
    .B(_00984_),
    .A_N(_06612_));
 sg13g2_and2_1 _15072_ (.A(_06603_),
    .B(_06613_),
    .X(_06614_));
 sg13g2_inv_1 _15073_ (.Y(_06615_),
    .A(_06614_));
 sg13g2_a21oi_1 _15074_ (.A1(_06611_),
    .A2(_06615_),
    .Y(_06616_),
    .B1(net3792));
 sg13g2_nor4_1 _15075_ (.A(net2436),
    .B(_01152_),
    .C(_06604_),
    .D(_06613_),
    .Y(_06617_));
 sg13g2_nor2_2 _15076_ (.A(_06595_),
    .B(_06612_),
    .Y(_06618_));
 sg13g2_nor3_1 _15077_ (.A(_06606_),
    .B(_06611_),
    .C(_06618_),
    .Y(_06619_));
 sg13g2_nor4_1 _15078_ (.A(net2299),
    .B(_06616_),
    .C(_06617_),
    .D(_06619_),
    .Y(_06620_));
 sg13g2_nor2_1 _15079_ (.A(net3792),
    .B(_01912_),
    .Y(_06621_));
 sg13g2_nor3_1 _15080_ (.A(net1731),
    .B(_06620_),
    .C(_06621_),
    .Y(_00705_));
 sg13g2_and2_1 _15081_ (.A(net3707),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .X(_06622_));
 sg13g2_nor2b_1 _15082_ (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .B_N(_06612_),
    .Y(_06623_));
 sg13g2_nor3_1 _15083_ (.A(_06595_),
    .B(_06606_),
    .C(_06623_),
    .Y(_06624_));
 sg13g2_o21ai_1 _15084_ (.B1(_06624_),
    .Y(_06625_),
    .A1(_06612_),
    .A2(_06622_));
 sg13g2_mux2_1 _15085_ (.A0(_06622_),
    .A1(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .S(_06608_),
    .X(_06626_));
 sg13g2_nand3_1 _15086_ (.B(_06605_),
    .C(_06626_),
    .A(_06595_),
    .Y(_06627_));
 sg13g2_a21oi_1 _15087_ (.A1(_06606_),
    .A2(_06622_),
    .Y(_06628_),
    .B1(_06603_));
 sg13g2_nand3_1 _15088_ (.B(_06627_),
    .C(_06628_),
    .A(_06625_),
    .Y(_06629_));
 sg13g2_nor2_1 _15089_ (.A(_06604_),
    .B(_06622_),
    .Y(_06630_));
 sg13g2_nor2_1 _15090_ (.A(net2299),
    .B(_06630_),
    .Y(_06631_));
 sg13g2_a22oi_1 _15091_ (.Y(_06632_),
    .B1(_06629_),
    .B2(_06631_),
    .A2(_01911_),
    .A1(net3707));
 sg13g2_nor2_1 _15092_ (.A(_05884_),
    .B(net3708),
    .Y(_00706_));
 sg13g2_nand2_1 _15093_ (.Y(_06633_),
    .A(net3789),
    .B(net1753));
 sg13g2_nand3_1 _15094_ (.B(_00928_),
    .C(net1753),
    .A(\addr[24] ),
    .Y(_06634_));
 sg13g2_nand3_1 _15095_ (.B(net3444),
    .C(net1753),
    .A(net3789),
    .Y(_06635_));
 sg13g2_inv_1 _15096_ (.Y(_06636_),
    .A(_06635_));
 sg13g2_a21oi_1 _15097_ (.A1(_01097_),
    .A2(_06636_),
    .Y(_06637_),
    .B1(net1750));
 sg13g2_o21ai_1 _15098_ (.B1(_06637_),
    .Y(_06638_),
    .A1(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .A2(_06634_));
 sg13g2_nor2_1 _15099_ (.A(net3753),
    .B(_06603_),
    .Y(_06639_));
 sg13g2_a21oi_1 _15100_ (.A1(_01911_),
    .A2(_06638_),
    .Y(_06640_),
    .B1(_06639_));
 sg13g2_nor2_1 _15101_ (.A(net3753),
    .B(_01912_),
    .Y(_06641_));
 sg13g2_nor3_1 _15102_ (.A(net1731),
    .B(_06640_),
    .C(_06641_),
    .Y(_00707_));
 sg13g2_nor2_1 _15103_ (.A(net2299),
    .B(_06598_),
    .Y(_06642_));
 sg13g2_a22oi_1 _15104_ (.Y(_06643_),
    .B1(_06642_),
    .B2(_06604_),
    .A2(_06638_),
    .A1(net2299));
 sg13g2_nand2_1 _15105_ (.Y(_06644_),
    .A(_06604_),
    .B(_06643_));
 sg13g2_a21o_1 _15106_ (.A2(_01912_),
    .A1(net3482),
    .B1(_06644_),
    .X(_06645_));
 sg13g2_nand2_1 _15107_ (.Y(_06646_),
    .A(net3482),
    .B(_06644_));
 sg13g2_a21oi_1 _15108_ (.A1(_06645_),
    .A2(_06646_),
    .Y(_00708_),
    .B1(net1730));
 sg13g2_nor2b_1 _15109_ (.A(net2436),
    .B_N(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .Y(_06647_));
 sg13g2_o21ai_1 _15110_ (.B1(_02417_),
    .Y(_06648_),
    .A1(net2427),
    .A2(_06647_));
 sg13g2_nor2b_1 _15111_ (.A(net3239),
    .B_N(_06648_),
    .Y(_06649_));
 sg13g2_nor3_1 _15112_ (.A(net2299),
    .B(_06644_),
    .C(_06649_),
    .Y(_06650_));
 sg13g2_a22oi_1 _15113_ (.Y(_06651_),
    .B1(_06650_),
    .B2(_06599_),
    .A2(_06645_),
    .A1(net3814));
 sg13g2_nor2_1 _15114_ (.A(net1730),
    .B(_06651_),
    .Y(_00709_));
 sg13g2_a21oi_1 _15115_ (.A1(_06604_),
    .A2(_06643_),
    .Y(_06652_),
    .B1(net3239));
 sg13g2_a21oi_1 _15116_ (.A1(net3789),
    .A2(net1753),
    .Y(_06653_),
    .B1(_01912_));
 sg13g2_o21ai_1 _15117_ (.B1(net3239),
    .Y(_06654_),
    .A1(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .A2(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ));
 sg13g2_nand3b_1 _15118_ (.B(_02412_),
    .C(_06600_),
    .Y(_06655_),
    .A_N(net2424));
 sg13g2_a21oi_1 _15119_ (.A1(_06654_),
    .A2(_06655_),
    .Y(_06656_),
    .B1(net2299));
 sg13g2_nor3_1 _15120_ (.A(_06644_),
    .B(_06653_),
    .C(_06656_),
    .Y(_06657_));
 sg13g2_nor3_1 _15121_ (.A(net1730),
    .B(_06652_),
    .C(_06657_),
    .Y(_00710_));
 sg13g2_nor2_1 _15122_ (.A(_06633_),
    .B(_06638_),
    .Y(_06658_));
 sg13g2_a22oi_1 _15123_ (.Y(_06659_),
    .B1(_06658_),
    .B2(_02802_),
    .A2(_06638_),
    .A1(net2436));
 sg13g2_nor2_1 _15124_ (.A(net1730),
    .B(_06659_),
    .Y(_00711_));
 sg13g2_nand2_1 _15125_ (.Y(_06660_),
    .A(_06600_),
    .B(_06604_));
 sg13g2_a21oi_1 _15126_ (.A1(_06605_),
    .A2(_06618_),
    .Y(_06661_),
    .B1(_06603_));
 sg13g2_nor4_1 _15127_ (.A(net2437),
    .B(_05884_),
    .C(_06614_),
    .D(_06661_),
    .Y(_00712_));
 sg13g2_nand3_1 _15128_ (.B(_06598_),
    .C(_06601_),
    .A(_06593_),
    .Y(_06662_));
 sg13g2_o21ai_1 _15129_ (.B1(_06643_),
    .Y(_06663_),
    .A1(net2299),
    .A2(_06662_));
 sg13g2_nand2b_2 _15130_ (.Y(_06664_),
    .B(_06615_),
    .A_N(_06663_));
 sg13g2_a21oi_1 _15131_ (.A1(_02417_),
    .A2(_06647_),
    .Y(_06665_),
    .B1(net2427));
 sg13g2_nor4_1 _15132_ (.A(net2299),
    .B(_06618_),
    .C(_06660_),
    .D(_06665_),
    .Y(_06666_));
 sg13g2_nor3_1 _15133_ (.A(_06653_),
    .B(_06664_),
    .C(_06666_),
    .Y(_06667_));
 sg13g2_a21oi_1 _15134_ (.A1(net2427),
    .A2(_06664_),
    .Y(_06668_),
    .B1(_06667_));
 sg13g2_nor2_1 _15135_ (.A(net1731),
    .B(_06668_),
    .Y(_00713_));
 sg13g2_nor2b_1 _15136_ (.A(net3279),
    .B_N(_06663_),
    .Y(_06669_));
 sg13g2_and3_1 _15137_ (.X(_06670_),
    .A(net2350),
    .B(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .C(_06603_));
 sg13g2_nor3_1 _15138_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .B(net2427),
    .C(net2436),
    .Y(_06671_));
 sg13g2_a21o_1 _15139_ (.A2(_06671_),
    .A1(net2426),
    .B1(_02412_),
    .X(_06672_));
 sg13g2_nor2b_1 _15140_ (.A(_06672_),
    .B_N(_06593_),
    .Y(_06673_));
 sg13g2_nor3_1 _15141_ (.A(_06618_),
    .B(_06660_),
    .C(_06673_),
    .Y(_06674_));
 sg13g2_nor4_1 _15142_ (.A(_06653_),
    .B(_06664_),
    .C(_06670_),
    .D(_06674_),
    .Y(_06675_));
 sg13g2_nor3_1 _15143_ (.A(net1731),
    .B(_06669_),
    .C(_06675_),
    .Y(_00714_));
 sg13g2_nor2b_1 _15144_ (.A(net2424),
    .B_N(_06663_),
    .Y(_06676_));
 sg13g2_nand3b_1 _15145_ (.B(_06600_),
    .C(_06672_),
    .Y(_06677_),
    .A_N(net2424));
 sg13g2_a21oi_1 _15146_ (.A1(_01912_),
    .A2(_06677_),
    .Y(_06678_),
    .B1(_06664_));
 sg13g2_nor3_1 _15147_ (.A(net1731),
    .B(_06676_),
    .C(_06678_),
    .Y(_00715_));
 sg13g2_a21oi_1 _15148_ (.A1(net2800),
    .A2(_06638_),
    .Y(_06679_),
    .B1(net1730));
 sg13g2_o21ai_1 _15149_ (.B1(_06679_),
    .Y(_00716_),
    .A1(_06636_),
    .A2(_06638_));
 sg13g2_a22oi_1 _15150_ (.Y(_06680_),
    .B1(_06638_),
    .B2(net2789),
    .A2(_06637_),
    .A1(_06634_));
 sg13g2_nand2b_1 _15151_ (.Y(_00717_),
    .B(net3517),
    .A_N(net1730));
 sg13g2_a21oi_1 _15152_ (.A1(net3857),
    .A2(_06638_),
    .Y(_06681_),
    .B1(net1730));
 sg13g2_nand2b_1 _15153_ (.Y(_00718_),
    .B(_06681_),
    .A_N(_06658_));
 sg13g2_nand2b_1 _15154_ (.Y(_06682_),
    .B(_02810_),
    .A_N(_06647_));
 sg13g2_o21ai_1 _15155_ (.B1(_02413_),
    .Y(_06683_),
    .A1(_06660_),
    .A2(_06682_));
 sg13g2_nor3_1 _15156_ (.A(net2424),
    .B(_06663_),
    .C(_06683_),
    .Y(_06684_));
 sg13g2_nor2_1 _15157_ (.A(net3508),
    .B(_06684_),
    .Y(_06685_));
 sg13g2_nor2b_1 _15158_ (.A(_01910_),
    .B_N(_06684_),
    .Y(_06686_));
 sg13g2_nor3_1 _15159_ (.A(net1730),
    .B(net3509),
    .C(_06686_),
    .Y(_00719_));
 sg13g2_nor2_1 _15160_ (.A(_01894_),
    .B(_05916_),
    .Y(_06687_));
 sg13g2_nor2_1 _15161_ (.A(_01360_),
    .B(_05915_),
    .Y(_06688_));
 sg13g2_nor3_1 _15162_ (.A(_05917_),
    .B(_06687_),
    .C(_06688_),
    .Y(_06689_));
 sg13g2_a21oi_1 _15163_ (.A1(_01341_),
    .A2(_05917_),
    .Y(_06690_),
    .B1(_06689_));
 sg13g2_nand2_1 _15164_ (.Y(_06691_),
    .A(net3651),
    .B(net2157));
 sg13g2_o21ai_1 _15165_ (.B1(_06691_),
    .Y(_00720_),
    .A1(_05914_),
    .A2(_06690_));
 sg13g2_nand2_1 _15166_ (.Y(_06692_),
    .A(net3697),
    .B(_05912_));
 sg13g2_nand2b_1 _15167_ (.Y(_06693_),
    .B(_05915_),
    .A_N(_02102_));
 sg13g2_a21oi_1 _15168_ (.A1(_01328_),
    .A2(_05916_),
    .Y(_06694_),
    .B1(_05917_));
 sg13g2_a22oi_1 _15169_ (.Y(_06695_),
    .B1(_06693_),
    .B2(_06694_),
    .A2(_05917_),
    .A1(_01305_));
 sg13g2_o21ai_1 _15170_ (.B1(_06692_),
    .Y(_00721_),
    .A1(_05914_),
    .A2(_06695_));
 sg13g2_nor4_2 _15171_ (.A(net2437),
    .B(_00984_),
    .C(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .Y(_06696_),
    .D(_06604_));
 sg13g2_mux2_1 _15172_ (.A0(net3155),
    .A1(net10),
    .S(_06696_),
    .X(_00722_));
 sg13g2_mux2_1 _15173_ (.A0(net3131),
    .A1(net11),
    .S(_06696_),
    .X(_00723_));
 sg13g2_mux2_1 _15174_ (.A0(net3138),
    .A1(net12),
    .S(_06696_),
    .X(_00724_));
 sg13g2_mux2_1 _15175_ (.A0(net3170),
    .A1(net13),
    .S(_06696_),
    .X(_00725_));
 sg13g2_nand2_1 _15176_ (.Y(_06697_),
    .A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .B(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_xor2_1 _15177_ (.B(\i_tinyqv.mem.q_ctrl.data_req ),
    .A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .X(_06698_));
 sg13g2_xnor2_1 _15178_ (.Y(_06699_),
    .A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .B(\i_tinyqv.mem.q_ctrl.data_req ));
 sg13g2_xnor2_1 _15179_ (.Y(_06700_),
    .A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .B(_06697_));
 sg13g2_nor2_2 _15180_ (.A(_06600_),
    .B(_06603_),
    .Y(_06701_));
 sg13g2_o21ai_1 _15181_ (.B1(net2436),
    .Y(_06702_),
    .A1(_06600_),
    .A2(_06603_));
 sg13g2_a21oi_1 _15182_ (.A1(_06602_),
    .A2(net2152),
    .Y(_06703_),
    .B1(_06639_));
 sg13g2_nor4_1 _15183_ (.A(net2437),
    .B(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .C(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .D(_06595_),
    .Y(_06704_));
 sg13g2_nor2_2 _15184_ (.A(_06703_),
    .B(_06704_),
    .Y(_06705_));
 sg13g2_or2_1 _15185_ (.X(_06706_),
    .B(_06704_),
    .A(_06703_));
 sg13g2_and2_1 _15186_ (.A(_02416_),
    .B(_06597_),
    .X(_06707_));
 sg13g2_nand2_1 _15187_ (.Y(_06708_),
    .A(net2422),
    .B(net2005));
 sg13g2_nand2_1 _15188_ (.Y(_06709_),
    .A(net3342),
    .B(net2294));
 sg13g2_nand2_1 _15189_ (.Y(_06710_),
    .A(net2851),
    .B(net2290));
 sg13g2_nand3_1 _15190_ (.B(_06709_),
    .C(_06710_),
    .A(net2188),
    .Y(_06711_));
 sg13g2_nand2_1 _15191_ (.Y(_06712_),
    .A(net2949),
    .B(net2293));
 sg13g2_a21oi_1 _15192_ (.A1(\i_tinyqv.cpu.instr_data_in[0] ),
    .A2(net2291),
    .Y(_06713_),
    .B1(net2187));
 sg13g2_a21oi_1 _15193_ (.A1(_06712_),
    .A2(_06713_),
    .Y(_06714_),
    .B1(_06701_));
 sg13g2_a221oi_1 _15194_ (.B2(_06714_),
    .C1(net2350),
    .B1(_06711_),
    .A1(net10),
    .Y(_06715_),
    .A2(_06701_));
 sg13g2_mux2_1 _15195_ (.A0(net3155),
    .A1(net10),
    .S(_06707_),
    .X(_06716_));
 sg13g2_o21ai_1 _15196_ (.B1(_06706_),
    .Y(_06717_),
    .A1(net2437),
    .A2(_06716_));
 sg13g2_o21ai_1 _15197_ (.B1(_06708_),
    .Y(_00726_),
    .A1(_06715_),
    .A2(_06717_));
 sg13g2_nand2_1 _15198_ (.Y(_06718_),
    .A(net3990),
    .B(_06705_));
 sg13g2_nand2_1 _15199_ (.Y(_06719_),
    .A(\i_tinyqv.mem.qspi_data_buf[25] ),
    .B(net2294));
 sg13g2_nand2_1 _15200_ (.Y(_06720_),
    .A(net2839),
    .B(net2290));
 sg13g2_nand3_1 _15201_ (.B(_06719_),
    .C(_06720_),
    .A(net2188),
    .Y(_06721_));
 sg13g2_nand2_1 _15202_ (.Y(_06722_),
    .A(net3018),
    .B(net2293));
 sg13g2_a21oi_1 _15203_ (.A1(\i_tinyqv.cpu.instr_data_in[1] ),
    .A2(net2292),
    .Y(_06723_),
    .B1(net2188));
 sg13g2_a21oi_1 _15204_ (.A1(_06722_),
    .A2(_06723_),
    .Y(_06724_),
    .B1(_06701_));
 sg13g2_a221oi_1 _15205_ (.B2(_06724_),
    .C1(net2350),
    .B1(_06721_),
    .A1(net11),
    .Y(_06725_),
    .A2(_06701_));
 sg13g2_mux2_1 _15206_ (.A0(net3131),
    .A1(net11),
    .S(_06707_),
    .X(_06726_));
 sg13g2_o21ai_1 _15207_ (.B1(_06706_),
    .Y(_06727_),
    .A1(net2437),
    .A2(_06726_));
 sg13g2_o21ai_1 _15208_ (.B1(net3991),
    .Y(_00727_),
    .A1(_06725_),
    .A2(_06727_));
 sg13g2_nand2b_1 _15209_ (.Y(_06728_),
    .B(net2293),
    .A_N(net2931));
 sg13g2_o21ai_1 _15210_ (.B1(_06728_),
    .Y(_06729_),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .A2(net2293));
 sg13g2_o21ai_1 _15211_ (.B1(net2187),
    .Y(_06730_),
    .A1(\i_tinyqv.mem.qspi_data_buf[26] ),
    .A2(net2290));
 sg13g2_a21oi_1 _15212_ (.A1(_01131_),
    .A2(net2290),
    .Y(_06731_),
    .B1(_06730_));
 sg13g2_nor2_1 _15213_ (.A(_06701_),
    .B(_06731_),
    .Y(_06732_));
 sg13g2_o21ai_1 _15214_ (.B1(_06732_),
    .Y(_06733_),
    .A1(net2188),
    .A2(_06729_));
 sg13g2_nand2b_1 _15215_ (.Y(_06734_),
    .B(_06701_),
    .A_N(net12));
 sg13g2_nand3_1 _15216_ (.B(_06733_),
    .C(_06734_),
    .A(net2437),
    .Y(_06735_));
 sg13g2_mux2_1 _15217_ (.A0(net3138),
    .A1(net12),
    .S(_06707_),
    .X(_06736_));
 sg13g2_a21oi_1 _15218_ (.A1(_00983_),
    .A2(_06736_),
    .Y(_06737_),
    .B1(net2005));
 sg13g2_a22oi_1 _15219_ (.Y(_00728_),
    .B1(_06735_),
    .B2(_06737_),
    .A2(net2005),
    .A1(net2330));
 sg13g2_nand2_1 _15220_ (.Y(_06738_),
    .A(net3954),
    .B(net2005));
 sg13g2_a21oi_1 _15221_ (.A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .A2(net2292),
    .Y(_06739_),
    .B1(net2188));
 sg13g2_o21ai_1 _15222_ (.B1(_06739_),
    .Y(_06740_),
    .A1(_01135_),
    .A2(net2292));
 sg13g2_and2_1 _15223_ (.A(\i_tinyqv.mem.qspi_data_buf[27] ),
    .B(net2293),
    .X(_06741_));
 sg13g2_a21oi_1 _15224_ (.A1(\i_tinyqv.mem.data_from_read[19] ),
    .A2(net2291),
    .Y(_06742_),
    .B1(_06741_));
 sg13g2_a21oi_1 _15225_ (.A1(net2188),
    .A2(_06742_),
    .Y(_06743_),
    .B1(_06701_));
 sg13g2_a221oi_1 _15226_ (.B2(_06743_),
    .C1(_00983_),
    .B1(_06740_),
    .A1(net13),
    .Y(_06744_),
    .A2(_06701_));
 sg13g2_mux2_1 _15227_ (.A0(net3170),
    .A1(net13),
    .S(_06707_),
    .X(_06745_));
 sg13g2_o21ai_1 _15228_ (.B1(_06706_),
    .Y(_06746_),
    .A1(\i_tinyqv.mem.q_ctrl.is_writing ),
    .A2(_06745_));
 sg13g2_o21ai_1 _15229_ (.B1(_06738_),
    .Y(_00729_),
    .A1(_06744_),
    .A2(_06746_));
 sg13g2_nor2_1 _15230_ (.A(net2421),
    .B(_06706_),
    .Y(_06747_));
 sg13g2_a21oi_1 _15231_ (.A1(net2882),
    .A2(net2293),
    .Y(_06748_),
    .B1(net2188));
 sg13g2_o21ai_1 _15232_ (.B1(_06748_),
    .Y(_06749_),
    .A1(_01118_),
    .A2(net2293));
 sg13g2_and2_1 _15233_ (.A(\i_tinyqv.mem.data_from_read[20] ),
    .B(net2291),
    .X(_06750_));
 sg13g2_a21oi_1 _15234_ (.A1(net3321),
    .A2(net2294),
    .Y(_06751_),
    .B1(_06750_));
 sg13g2_a21oi_1 _15235_ (.A1(net2187),
    .A2(_06751_),
    .Y(_06752_),
    .B1(net2152));
 sg13g2_a22oi_1 _15236_ (.Y(_06753_),
    .B1(_06749_),
    .B2(_06752_),
    .A2(net2152),
    .A1(net2422));
 sg13g2_a21oi_1 _15237_ (.A1(_06706_),
    .A2(_06753_),
    .Y(_00730_),
    .B1(_06747_));
 sg13g2_nand2_1 _15238_ (.Y(_06754_),
    .A(net3611),
    .B(net2294));
 sg13g2_nand2_1 _15239_ (.Y(_06755_),
    .A(net3613),
    .B(net2290));
 sg13g2_nand3_1 _15240_ (.B(_06754_),
    .C(_06755_),
    .A(net2187),
    .Y(_06756_));
 sg13g2_nand2_1 _15241_ (.Y(_06757_),
    .A(net4086),
    .B(net2290));
 sg13g2_a21oi_1 _15242_ (.A1(net3087),
    .A2(net2294),
    .Y(_06758_),
    .B1(net2187));
 sg13g2_a21oi_1 _15243_ (.A1(_06757_),
    .A2(_06758_),
    .Y(_06759_),
    .B1(net2152));
 sg13g2_a221oi_1 _15244_ (.B2(_06759_),
    .C1(net2005),
    .B1(_06756_),
    .A1(net3990),
    .Y(_06760_),
    .A2(net2152));
 sg13g2_a21oi_1 _15245_ (.A1(_01125_),
    .A2(net2005),
    .Y(_00731_),
    .B1(_06760_));
 sg13g2_mux2_1 _15246_ (.A0(\i_tinyqv.cpu.instr_data_in[6] ),
    .A1(net3629),
    .S(net2294),
    .X(_06761_));
 sg13g2_and2_1 _15247_ (.A(net3593),
    .B(net2290),
    .X(_06762_));
 sg13g2_a21oi_1 _15248_ (.A1(net3659),
    .A2(net2294),
    .Y(_06763_),
    .B1(_06762_));
 sg13g2_a21oi_1 _15249_ (.A1(_06700_),
    .A2(_06763_),
    .Y(_06764_),
    .B1(net2152));
 sg13g2_o21ai_1 _15250_ (.B1(_06764_),
    .Y(_06765_),
    .A1(net2187),
    .A2(_06761_));
 sg13g2_a21oi_1 _15251_ (.A1(\i_tinyqv.cpu.instr_data_in[10] ),
    .A2(net2152),
    .Y(_06766_),
    .B1(net2005));
 sg13g2_a22oi_1 _15252_ (.Y(_00732_),
    .B1(_06765_),
    .B2(_06766_),
    .A2(net2005),
    .A1(_01129_));
 sg13g2_nor2_1 _15253_ (.A(net2419),
    .B(_06706_),
    .Y(_06767_));
 sg13g2_and2_1 _15254_ (.A(\i_tinyqv.mem.qspi_data_buf[31] ),
    .B(net2294),
    .X(_06768_));
 sg13g2_a21oi_1 _15255_ (.A1(net3493),
    .A2(net2290),
    .Y(_06769_),
    .B1(_06768_));
 sg13g2_nand2_1 _15256_ (.Y(_06770_),
    .A(net3932),
    .B(net2291));
 sg13g2_a21oi_1 _15257_ (.A1(net3664),
    .A2(net2293),
    .Y(_06771_),
    .B1(net2187));
 sg13g2_a221oi_1 _15258_ (.B2(_06771_),
    .C1(net2152),
    .B1(_06770_),
    .A1(net2187),
    .Y(_06772_),
    .A2(_06769_));
 sg13g2_a21oi_1 _15259_ (.A1(net3954),
    .A2(_06702_),
    .Y(_06773_),
    .B1(_06772_));
 sg13g2_a21oi_1 _15260_ (.A1(_06706_),
    .A2(_06773_),
    .Y(_00733_),
    .B1(_06767_));
 sg13g2_nand2b_1 _15261_ (.Y(_00734_),
    .B(net2256),
    .A_N(net2800));
 sg13g2_nand2b_1 _15262_ (.Y(_00735_),
    .B(net2256),
    .A_N(net2789));
 sg13g2_nor2_1 _15263_ (.A(net2246),
    .B(_02596_),
    .Y(_00736_));
 sg13g2_mux2_1 _15264_ (.A0(net12),
    .A1(net3380),
    .S(net2265),
    .X(_00737_));
 sg13g2_mux2_1 _15265_ (.A0(net3452),
    .A1(\i_tinyqv.cpu.instr_data_in[2] ),
    .S(net1737),
    .X(_00738_));
 sg13g2_mux2_1 _15266_ (.A0(net3440),
    .A1(\i_tinyqv.cpu.instr_data_in[3] ),
    .S(net1737),
    .X(_00739_));
 sg13g2_nor2_1 _15267_ (.A(net3157),
    .B(net1735),
    .Y(_06774_));
 sg13g2_a21oi_1 _15268_ (.A1(_01118_),
    .A2(net1735),
    .Y(_00740_),
    .B1(_06774_));
 sg13g2_mux2_1 _15269_ (.A0(net3521),
    .A1(\i_tinyqv.cpu.instr_data_in[5] ),
    .S(net1736),
    .X(_00741_));
 sg13g2_mux2_1 _15270_ (.A0(net3421),
    .A1(\i_tinyqv.cpu.instr_data_in[6] ),
    .S(net1734),
    .X(_00742_));
 sg13g2_nor2_1 _15271_ (.A(net3115),
    .B(net1734),
    .Y(_06775_));
 sg13g2_a21oi_1 _15272_ (.A1(_01134_),
    .A2(net1734),
    .Y(_00743_),
    .B1(_06775_));
 sg13g2_mux2_1 _15273_ (.A0(net3438),
    .A1(net2422),
    .S(net1734),
    .X(_00744_));
 sg13g2_nor2_1 _15274_ (.A(net3210),
    .B(net1734),
    .Y(_06776_));
 sg13g2_a21oi_1 _15275_ (.A1(_01124_),
    .A2(net1734),
    .Y(_00745_),
    .B1(_06776_));
 sg13g2_nor2_1 _15276_ (.A(net3230),
    .B(net1735),
    .Y(_06777_));
 sg13g2_a21oi_1 _15277_ (.A1(net2330),
    .A2(net1735),
    .Y(_00746_),
    .B1(_06777_));
 sg13g2_nor2_1 _15278_ (.A(net3079),
    .B(net1734),
    .Y(_06778_));
 sg13g2_a21oi_1 _15279_ (.A1(_01133_),
    .A2(net1734),
    .Y(_00747_),
    .B1(_06778_));
 sg13g2_mux2_1 _15280_ (.A0(net3428),
    .A1(net2421),
    .S(net1735),
    .X(_00748_));
 sg13g2_nor2_1 _15281_ (.A(net3106),
    .B(net1736),
    .Y(_06779_));
 sg13g2_a21oi_1 _15282_ (.A1(_01125_),
    .A2(net1736),
    .Y(_00749_),
    .B1(_06779_));
 sg13g2_nor2_1 _15283_ (.A(net3076),
    .B(net1737),
    .Y(_06780_));
 sg13g2_a21oi_1 _15284_ (.A1(_01129_),
    .A2(net1737),
    .Y(_00750_),
    .B1(net3077));
 sg13g2_mux2_1 _15285_ (.A0(net3711),
    .A1(\i_tinyqv.cpu.instr_data_in[15] ),
    .S(net1737),
    .X(_00751_));
 sg13g2_nor2_1 _15286_ (.A(_00946_),
    .B(_01346_),
    .Y(_06781_));
 sg13g2_nor3_1 _15287_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .C(_06781_),
    .Y(_06782_));
 sg13g2_o21ai_1 _15288_ (.B1(_06782_),
    .Y(_06783_),
    .A1(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .A2(_01343_));
 sg13g2_nor2_1 _15289_ (.A(_01960_),
    .B(_06783_),
    .Y(_06784_));
 sg13g2_nand2_1 _15290_ (.Y(_06785_),
    .A(_02334_),
    .B(_06784_));
 sg13g2_nand2_1 _15291_ (.Y(_06786_),
    .A(net3007),
    .B(net2235));
 sg13g2_o21ai_1 _15292_ (.B1(_06785_),
    .Y(_00752_),
    .A1(_06784_),
    .A2(_06786_));
 sg13g2_nor2_1 _15293_ (.A(_02475_),
    .B(_02639_),
    .Y(_06787_));
 sg13g2_nand2_1 _15294_ (.Y(_06788_),
    .A(_02476_),
    .B(_02638_));
 sg13g2_o21ai_1 _15295_ (.B1(_06274_),
    .Y(_06789_),
    .A1(_02167_),
    .A2(_02639_));
 sg13g2_inv_1 _15296_ (.Y(_06790_),
    .A(_06789_));
 sg13g2_o21ai_1 _15297_ (.B1(net2490),
    .Y(_06791_),
    .A1(net4078),
    .A2(net1768));
 sg13g2_a21oi_1 _15298_ (.A1(net1768),
    .A2(_06790_),
    .Y(_00753_),
    .B1(_06791_));
 sg13g2_a21o_1 _15299_ (.A2(_02475_),
    .A1(_02241_),
    .B1(_02640_),
    .X(_06792_));
 sg13g2_a22oi_1 _15300_ (.Y(_00754_),
    .B1(_06792_),
    .B2(_06281_),
    .A2(net1772),
    .A1(_00982_));
 sg13g2_nand2_2 _15301_ (.Y(_06793_),
    .A(_05171_),
    .B(net2189));
 sg13g2_nand2_1 _15302_ (.Y(_06794_),
    .A(net3111),
    .B(net2078));
 sg13g2_o21ai_1 _15303_ (.B1(_06794_),
    .Y(_00755_),
    .A1(_00974_),
    .A2(net2080));
 sg13g2_nand2_1 _15304_ (.Y(_06795_),
    .A(net2985),
    .B(net2078));
 sg13g2_o21ai_1 _15305_ (.B1(_06795_),
    .Y(_00756_),
    .A1(_00973_),
    .A2(net2080));
 sg13g2_nand2_1 _15306_ (.Y(_06796_),
    .A(net3180),
    .B(net2078));
 sg13g2_o21ai_1 _15307_ (.B1(_06796_),
    .Y(_00757_),
    .A1(_00972_),
    .A2(net2079));
 sg13g2_nand2_1 _15308_ (.Y(_06797_),
    .A(net3262),
    .B(net2078));
 sg13g2_o21ai_1 _15309_ (.B1(_06797_),
    .Y(_00758_),
    .A1(_00971_),
    .A2(net2079));
 sg13g2_nand2_1 _15310_ (.Y(_06798_),
    .A(net3158),
    .B(net2074));
 sg13g2_o21ai_1 _15311_ (.B1(_06798_),
    .Y(_00759_),
    .A1(_00970_),
    .A2(net2075));
 sg13g2_nand2_1 _15312_ (.Y(_06799_),
    .A(net3032),
    .B(net2078));
 sg13g2_o21ai_1 _15313_ (.B1(_06799_),
    .Y(_00760_),
    .A1(net2352),
    .A2(net2078));
 sg13g2_nand2_1 _15314_ (.Y(_06800_),
    .A(net3100),
    .B(net2079));
 sg13g2_o21ai_1 _15315_ (.B1(_06800_),
    .Y(_00761_),
    .A1(_00968_),
    .A2(net2079));
 sg13g2_nand2_1 _15316_ (.Y(_06801_),
    .A(net3241),
    .B(net2074));
 sg13g2_o21ai_1 _15317_ (.B1(_06801_),
    .Y(_00762_),
    .A1(_00967_),
    .A2(net2074));
 sg13g2_mux2_1 _15318_ (.A0(\data_to_write[8] ),
    .A1(net3530),
    .S(net2079),
    .X(_00763_));
 sg13g2_mux2_1 _15319_ (.A0(\data_to_write[9] ),
    .A1(net3582),
    .S(net2074),
    .X(_00764_));
 sg13g2_mux2_1 _15320_ (.A0(\data_to_write[10] ),
    .A1(net3672),
    .S(net2079),
    .X(_00765_));
 sg13g2_mux2_1 _15321_ (.A0(\data_to_write[11] ),
    .A1(net3500),
    .S(net2078),
    .X(_00766_));
 sg13g2_mux2_1 _15322_ (.A0(\data_to_write[12] ),
    .A1(net3488),
    .S(net2079),
    .X(_00767_));
 sg13g2_nand2_1 _15323_ (.Y(_06802_),
    .A(net3020),
    .B(net2076));
 sg13g2_o21ai_1 _15324_ (.B1(_06802_),
    .Y(_00768_),
    .A1(_00965_),
    .A2(net2076));
 sg13g2_nand2_1 _15325_ (.Y(_06803_),
    .A(net2935),
    .B(net2077));
 sg13g2_o21ai_1 _15326_ (.B1(_06803_),
    .Y(_00769_),
    .A1(_00964_),
    .A2(net2077));
 sg13g2_nand2_1 _15327_ (.Y(_06804_),
    .A(net2878),
    .B(net2075));
 sg13g2_o21ai_1 _15328_ (.B1(_06804_),
    .Y(_00770_),
    .A1(_00963_),
    .A2(net2073));
 sg13g2_nand2_1 _15329_ (.Y(_06805_),
    .A(net2902),
    .B(net2076));
 sg13g2_o21ai_1 _15330_ (.B1(_06805_),
    .Y(_00771_),
    .A1(_00962_),
    .A2(net2076));
 sg13g2_nand2_1 _15331_ (.Y(_06806_),
    .A(net2847),
    .B(net2072));
 sg13g2_o21ai_1 _15332_ (.B1(_06806_),
    .Y(_00772_),
    .A1(_00961_),
    .A2(net2072));
 sg13g2_nand2_1 _15333_ (.Y(_06807_),
    .A(net2953),
    .B(net2076));
 sg13g2_o21ai_1 _15334_ (.B1(_06807_),
    .Y(_00773_),
    .A1(_00960_),
    .A2(net2076));
 sg13g2_nand2_1 _15335_ (.Y(_06808_),
    .A(net2880),
    .B(net2073));
 sg13g2_o21ai_1 _15336_ (.B1(_06808_),
    .Y(_00774_),
    .A1(_00959_),
    .A2(net2073));
 sg13g2_mux2_1 _15337_ (.A0(\data_to_write[20] ),
    .A1(net3514),
    .S(net2073),
    .X(_00775_));
 sg13g2_nand2_1 _15338_ (.Y(_06809_),
    .A(net2841),
    .B(net2072));
 sg13g2_o21ai_1 _15339_ (.B1(_06809_),
    .Y(_00776_),
    .A1(_00958_),
    .A2(net2072));
 sg13g2_nand2_1 _15340_ (.Y(_06810_),
    .A(net2913),
    .B(net2072));
 sg13g2_o21ai_1 _15341_ (.B1(_06810_),
    .Y(_00777_),
    .A1(_00957_),
    .A2(net2072));
 sg13g2_nand2_1 _15342_ (.Y(_06811_),
    .A(net3049),
    .B(net2074));
 sg13g2_o21ai_1 _15343_ (.B1(_06811_),
    .Y(_00778_),
    .A1(_00956_),
    .A2(net2074));
 sg13g2_nand2_1 _15344_ (.Y(_06812_),
    .A(net2876),
    .B(net2074));
 sg13g2_o21ai_1 _15345_ (.B1(_06812_),
    .Y(_00779_),
    .A1(_00955_),
    .A2(net2074));
 sg13g2_nand2_1 _15346_ (.Y(_06813_),
    .A(net2807),
    .B(net2075));
 sg13g2_o21ai_1 _15347_ (.B1(_06813_),
    .Y(_00780_),
    .A1(_00954_),
    .A2(net2075));
 sg13g2_nand2_1 _15348_ (.Y(_06814_),
    .A(net2826),
    .B(net2072));
 sg13g2_o21ai_1 _15349_ (.B1(_06814_),
    .Y(_00781_),
    .A1(_00953_),
    .A2(net2072));
 sg13g2_nand2_1 _15350_ (.Y(_06815_),
    .A(net2811),
    .B(net2076));
 sg13g2_o21ai_1 _15351_ (.B1(_06815_),
    .Y(_00782_),
    .A1(_00952_),
    .A2(net2077));
 sg13g2_nand2_1 _15352_ (.Y(_06816_),
    .A(net2874),
    .B(net2073));
 sg13g2_o21ai_1 _15353_ (.B1(_06816_),
    .Y(_00783_),
    .A1(_00951_),
    .A2(net2073));
 sg13g2_nand2_1 _15354_ (.Y(_06817_),
    .A(net2819),
    .B(net2078));
 sg13g2_o21ai_1 _15355_ (.B1(_06817_),
    .Y(_00784_),
    .A1(_00950_),
    .A2(net2077));
 sg13g2_nand2_1 _15356_ (.Y(_06818_),
    .A(net3134),
    .B(net2077));
 sg13g2_o21ai_1 _15357_ (.B1(_06818_),
    .Y(_00785_),
    .A1(_00949_),
    .A2(net2077));
 sg13g2_nand2_1 _15358_ (.Y(_06819_),
    .A(net3005),
    .B(net2076));
 sg13g2_o21ai_1 _15359_ (.B1(_06819_),
    .Y(_00786_),
    .A1(_00948_),
    .A2(net2073));
 sg13g2_nand2_1 _15360_ (.Y(_06820_),
    .A(_02341_),
    .B(net1809));
 sg13g2_a21oi_1 _15361_ (.A1(net2747),
    .A2(net1812),
    .Y(_06821_),
    .B1(net1862));
 sg13g2_mux2_1 _15362_ (.A0(\i_tinyqv.cpu.i_core.mepc[3] ),
    .A1(net2460),
    .S(net2222),
    .X(_06822_));
 sg13g2_nand2_1 _15363_ (.Y(_06823_),
    .A(net2240),
    .B(_05301_));
 sg13g2_a21oi_1 _15364_ (.A1(_01216_),
    .A2(_06822_),
    .Y(_06824_),
    .B1(net1855));
 sg13g2_a221oi_1 _15365_ (.B2(_06824_),
    .C1(net1771),
    .B1(_06823_),
    .A1(_06820_),
    .Y(_06825_),
    .A2(_06821_));
 sg13g2_a21oi_1 _15366_ (.A1(net2418),
    .A2(net1771),
    .Y(_06826_),
    .B1(_06825_));
 sg13g2_nor2_1 _15367_ (.A(net2342),
    .B(_06826_),
    .Y(_00787_));
 sg13g2_nand2_1 _15368_ (.Y(_06827_),
    .A(_01984_),
    .B(net1809));
 sg13g2_and2_1 _15369_ (.A(net2459),
    .B(net2222),
    .X(_06828_));
 sg13g2_a21oi_2 _15370_ (.B1(_06828_),
    .Y(_06829_),
    .A2(net2186),
    .A1(net3579));
 sg13g2_nand2_1 _15371_ (.Y(_06830_),
    .A(net2306),
    .B(_06829_));
 sg13g2_o21ai_1 _15372_ (.B1(_06830_),
    .Y(_06831_),
    .A1(net2306),
    .A2(_06286_));
 sg13g2_a21oi_1 _15373_ (.A1(net2740),
    .A2(net1812),
    .Y(_06832_),
    .B1(net1861));
 sg13g2_a221oi_1 _15374_ (.B2(_06827_),
    .C1(net1771),
    .B1(_06832_),
    .A1(net1861),
    .Y(_06833_),
    .A2(_06831_));
 sg13g2_a21oi_1 _15375_ (.A1(net2417),
    .A2(net1771),
    .Y(_06834_),
    .B1(_06833_));
 sg13g2_nor2_1 _15376_ (.A(net2340),
    .B(_06834_),
    .Y(_00788_));
 sg13g2_a21oi_1 _15377_ (.A1(net2734),
    .A2(net1812),
    .Y(_06835_),
    .B1(net1862));
 sg13g2_o21ai_1 _15378_ (.B1(_06835_),
    .Y(_06836_),
    .A1(_02166_),
    .A2(net1813));
 sg13g2_and2_1 _15379_ (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .B(net2222),
    .X(_06837_));
 sg13g2_a21oi_2 _15380_ (.B1(_06837_),
    .Y(_06838_),
    .A2(net2186),
    .A1(net3765));
 sg13g2_o21ai_1 _15381_ (.B1(net1861),
    .Y(_06839_),
    .A1(net2240),
    .A2(_06838_));
 sg13g2_a21oi_1 _15382_ (.A1(net2240),
    .A2(_06296_),
    .Y(_06840_),
    .B1(_06839_));
 sg13g2_nor2_1 _15383_ (.A(net1772),
    .B(_06840_),
    .Y(_06841_));
 sg13g2_a22oi_1 _15384_ (.Y(_06842_),
    .B1(_06836_),
    .B2(_06841_),
    .A2(net1771),
    .A1(net4011));
 sg13g2_nor2_1 _15385_ (.A(net2342),
    .B(_06842_),
    .Y(_00789_));
 sg13g2_nand2_1 _15386_ (.Y(_06843_),
    .A(net2729),
    .B(net1812));
 sg13g2_o21ai_1 _15387_ (.B1(_06843_),
    .Y(_06844_),
    .A1(_02240_),
    .A2(net1812));
 sg13g2_mux2_1 _15388_ (.A0(net3325),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .S(net2219),
    .X(_06845_));
 sg13g2_nand2_1 _15389_ (.Y(_06846_),
    .A(net2306),
    .B(_06845_));
 sg13g2_o21ai_1 _15390_ (.B1(_06846_),
    .Y(_06847_),
    .A1(net2306),
    .A2(_06309_));
 sg13g2_nand2_1 _15391_ (.Y(_06848_),
    .A(net1855),
    .B(_06844_));
 sg13g2_a21oi_1 _15392_ (.A1(net1861),
    .A2(_06847_),
    .Y(_06849_),
    .B1(net1771));
 sg13g2_a221oi_1 _15393_ (.B2(_06849_),
    .C1(net2342),
    .B1(_06848_),
    .A1(_00981_),
    .Y(_00790_),
    .A2(net1771));
 sg13g2_nand2_1 _15394_ (.Y(_06850_),
    .A(net2707),
    .B(net1811));
 sg13g2_o21ai_1 _15395_ (.B1(_06850_),
    .Y(_06851_),
    .A1(_02340_),
    .A2(net1812));
 sg13g2_nand2_1 _15396_ (.Y(_06852_),
    .A(net1855),
    .B(_06851_));
 sg13g2_mux2_1 _15397_ (.A0(\i_tinyqv.cpu.i_core.mepc[7] ),
    .A1(net2456),
    .S(net2221),
    .X(_06853_));
 sg13g2_mux2_1 _15398_ (.A0(_06319_),
    .A1(_06853_),
    .S(net2306),
    .X(_06854_));
 sg13g2_a21oi_1 _15399_ (.A1(net1861),
    .A2(_06854_),
    .Y(_06855_),
    .B1(net1771));
 sg13g2_o21ai_1 _15400_ (.B1(net2491),
    .Y(_06856_),
    .A1(net2416),
    .A2(net1768));
 sg13g2_a21oi_1 _15401_ (.A1(_06852_),
    .A2(_06855_),
    .Y(_00791_),
    .B1(_06856_));
 sg13g2_nand2_1 _15402_ (.Y(_06857_),
    .A(net2699),
    .B(net1811));
 sg13g2_a21oi_1 _15403_ (.A1(_01982_),
    .A2(net1808),
    .Y(_06858_),
    .B1(net1860));
 sg13g2_and2_1 _15404_ (.A(net3538),
    .B(net2221),
    .X(_06859_));
 sg13g2_a21oi_2 _15405_ (.B1(_06859_),
    .Y(_06860_),
    .A2(net2186),
    .A1(net3581));
 sg13g2_nand2_1 _15406_ (.Y(_06861_),
    .A(net2304),
    .B(_06860_));
 sg13g2_o21ai_1 _15407_ (.B1(_06861_),
    .Y(_06862_),
    .A1(net2305),
    .A2(_06332_));
 sg13g2_a221oi_1 _15408_ (.B2(net1860),
    .C1(net1770),
    .B1(_06862_),
    .A1(_06857_),
    .Y(_06863_),
    .A2(_06858_));
 sg13g2_a21oi_1 _15409_ (.A1(net3896),
    .A2(net1770),
    .Y(_06864_),
    .B1(_06863_));
 sg13g2_nor2_1 _15410_ (.A(net2340),
    .B(_06864_),
    .Y(_00792_));
 sg13g2_a21oi_1 _15411_ (.A1(net2673),
    .A2(net1811),
    .Y(_06865_),
    .B1(net1860));
 sg13g2_o21ai_1 _15412_ (.B1(_06865_),
    .Y(_06866_),
    .A1(_02165_),
    .A2(net1813));
 sg13g2_and2_1 _15413_ (.A(net2454),
    .B(net2221),
    .X(_06867_));
 sg13g2_a21oi_2 _15414_ (.B1(_06867_),
    .Y(_06868_),
    .A2(net2186),
    .A1(net3565));
 sg13g2_nand2_1 _15415_ (.Y(_06869_),
    .A(net2305),
    .B(_06868_));
 sg13g2_o21ai_1 _15416_ (.B1(_06869_),
    .Y(_06870_),
    .A1(net2305),
    .A2(_06341_));
 sg13g2_a21oi_1 _15417_ (.A1(net1860),
    .A2(_06870_),
    .Y(_06871_),
    .B1(net1772));
 sg13g2_a22oi_1 _15418_ (.Y(_06872_),
    .B1(_06866_),
    .B2(_06871_),
    .A2(net1770),
    .A1(net3873));
 sg13g2_nor2_1 _15419_ (.A(net2340),
    .B(_06872_),
    .Y(_00793_));
 sg13g2_nand2_1 _15420_ (.Y(_06873_),
    .A(_02239_),
    .B(net1807));
 sg13g2_a21oi_1 _15421_ (.A1(net2694),
    .A2(net1811),
    .Y(_06874_),
    .B1(net1857));
 sg13g2_nand2_1 _15422_ (.Y(_06875_),
    .A(net2238),
    .B(_06350_));
 sg13g2_mux2_1 _15423_ (.A0(\i_tinyqv.cpu.i_core.mepc[10] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .S(net2220),
    .X(_06876_));
 sg13g2_a21oi_1 _15424_ (.A1(net2304),
    .A2(_06876_),
    .Y(_06877_),
    .B1(net1856));
 sg13g2_a221oi_1 _15425_ (.B2(_06877_),
    .C1(net1769),
    .B1(_06875_),
    .A1(_06873_),
    .Y(_06878_),
    .A2(_06874_));
 sg13g2_a21oi_1 _15426_ (.A1(net2415),
    .A2(net1769),
    .Y(_06879_),
    .B1(_06878_));
 sg13g2_nor2_1 _15427_ (.A(net2341),
    .B(_06879_),
    .Y(_00794_));
 sg13g2_and2_1 _15428_ (.A(net2452),
    .B(net2221),
    .X(_06880_));
 sg13g2_a21oi_2 _15429_ (.B1(_06880_),
    .Y(_06881_),
    .A2(net2186),
    .A1(net3513));
 sg13g2_nor2_1 _15430_ (.A(net2304),
    .B(_06362_),
    .Y(_06882_));
 sg13g2_a21oi_1 _15431_ (.A1(net2304),
    .A2(_06881_),
    .Y(_06883_),
    .B1(_06882_));
 sg13g2_a21oi_1 _15432_ (.A1(net2696),
    .A2(net1810),
    .Y(_06884_),
    .B1(net1859));
 sg13g2_o21ai_1 _15433_ (.B1(_06884_),
    .Y(_06885_),
    .A1(_02345_),
    .A2(net1810));
 sg13g2_o21ai_1 _15434_ (.B1(_06885_),
    .Y(_06886_),
    .A1(net1856),
    .A2(_06883_));
 sg13g2_o21ai_1 _15435_ (.B1(net2484),
    .Y(_06887_),
    .A1(net4054),
    .A2(net1766));
 sg13g2_a21oi_1 _15436_ (.A1(net1766),
    .A2(_06886_),
    .Y(_00795_),
    .B1(_06887_));
 sg13g2_mux2_1 _15437_ (.A0(net2681),
    .A1(_01980_),
    .S(net1807),
    .X(_06888_));
 sg13g2_nand2_1 _15438_ (.Y(_06889_),
    .A(net2238),
    .B(_06371_));
 sg13g2_mux2_1 _15439_ (.A0(\i_tinyqv.cpu.i_core.mepc[12] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .S(net2221),
    .X(_06890_));
 sg13g2_nand2_1 _15440_ (.Y(_06891_),
    .A(net2304),
    .B(_06890_));
 sg13g2_nand3_1 _15441_ (.B(_06889_),
    .C(_06891_),
    .A(net1859),
    .Y(_06892_));
 sg13g2_o21ai_1 _15442_ (.B1(_06892_),
    .Y(_06893_),
    .A1(net1859),
    .A2(_06888_));
 sg13g2_o21ai_1 _15443_ (.B1(net2484),
    .Y(_06894_),
    .A1(net4074),
    .A2(net1766));
 sg13g2_a21oi_1 _15444_ (.A1(net1766),
    .A2(_06893_),
    .Y(_00796_),
    .B1(_06894_));
 sg13g2_mux2_1 _15445_ (.A0(\i_tinyqv.cpu.i_core.mepc[13] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .S(net2219),
    .X(_06895_));
 sg13g2_mux2_1 _15446_ (.A0(_06380_),
    .A1(_06895_),
    .S(net2304),
    .X(_06896_));
 sg13g2_a21oi_1 _15447_ (.A1(net2683),
    .A2(net1810),
    .Y(_06897_),
    .B1(net1859));
 sg13g2_o21ai_1 _15448_ (.B1(_06897_),
    .Y(_06898_),
    .A1(_02164_),
    .A2(net1810));
 sg13g2_o21ai_1 _15449_ (.B1(_06898_),
    .Y(_06899_),
    .A1(net1856),
    .A2(_06896_));
 sg13g2_o21ai_1 _15450_ (.B1(net2484),
    .Y(_06900_),
    .A1(net2414),
    .A2(net1766));
 sg13g2_a21oi_1 _15451_ (.A1(net1766),
    .A2(_06899_),
    .Y(_00797_),
    .B1(_06900_));
 sg13g2_a21oi_1 _15452_ (.A1(net2711),
    .A2(net1811),
    .Y(_06901_),
    .B1(net1857));
 sg13g2_o21ai_1 _15453_ (.B1(_06901_),
    .Y(_06902_),
    .A1(_02238_),
    .A2(net1810));
 sg13g2_nand2_1 _15454_ (.Y(_06903_),
    .A(net2239),
    .B(_06392_));
 sg13g2_mux2_1 _15455_ (.A0(\i_tinyqv.cpu.i_core.mepc[14] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .S(net2219),
    .X(_06904_));
 sg13g2_nand2_1 _15456_ (.Y(_06905_),
    .A(net2304),
    .B(_06904_));
 sg13g2_nand3_1 _15457_ (.B(_06903_),
    .C(_06905_),
    .A(net1857),
    .Y(_06906_));
 sg13g2_a21oi_1 _15458_ (.A1(_06902_),
    .A2(_06906_),
    .Y(_06907_),
    .B1(net1770));
 sg13g2_o21ai_1 _15459_ (.B1(net2484),
    .Y(_06908_),
    .A1(net2413),
    .A2(net1767));
 sg13g2_nor2_1 _15460_ (.A(_06907_),
    .B(_06908_),
    .Y(_00798_));
 sg13g2_a21oi_1 _15461_ (.A1(_02338_),
    .A2(net1807),
    .Y(_06909_),
    .B1(net1859));
 sg13g2_o21ai_1 _15462_ (.B1(_06909_),
    .Y(_06910_),
    .A1(net2690),
    .A2(net1807));
 sg13g2_mux2_1 _15463_ (.A0(\i_tinyqv.cpu.i_core.mepc[15] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .S(net2219),
    .X(_06911_));
 sg13g2_mux2_1 _15464_ (.A0(_06402_),
    .A1(_06911_),
    .S(net2304),
    .X(_06912_));
 sg13g2_a21oi_1 _15465_ (.A1(net1859),
    .A2(_06912_),
    .Y(_06913_),
    .B1(net1769));
 sg13g2_a221oi_1 _15466_ (.B2(_06913_),
    .C1(net2340),
    .B1(_06910_),
    .A1(_00978_),
    .Y(_00799_),
    .A2(net1769));
 sg13g2_a21oi_1 _15467_ (.A1(_01156_),
    .A2(net1810),
    .Y(_06914_),
    .B1(net1859));
 sg13g2_o21ai_1 _15468_ (.B1(_06914_),
    .Y(_06915_),
    .A1(_01979_),
    .A2(net1810));
 sg13g2_mux2_1 _15469_ (.A0(\i_tinyqv.cpu.i_core.mepc[16] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .S(net2221),
    .X(_06916_));
 sg13g2_o21ai_1 _15470_ (.B1(net1857),
    .Y(_06917_),
    .A1(net2238),
    .A2(_06916_));
 sg13g2_a21oi_1 _15471_ (.A1(net2238),
    .A2(_06412_),
    .Y(_06918_),
    .B1(_06917_));
 sg13g2_nor2_1 _15472_ (.A(net1769),
    .B(_06918_),
    .Y(_06919_));
 sg13g2_o21ai_1 _15473_ (.B1(net2484),
    .Y(_06920_),
    .A1(net2412),
    .A2(net1766));
 sg13g2_a21oi_1 _15474_ (.A1(_06915_),
    .A2(_06919_),
    .Y(_00800_),
    .B1(_06920_));
 sg13g2_o21ai_1 _15475_ (.B1(net1856),
    .Y(_06921_),
    .A1(net2710),
    .A2(net1807));
 sg13g2_a21o_1 _15476_ (.A2(net1807),
    .A1(_02162_),
    .B1(_06921_),
    .X(_06922_));
 sg13g2_mux2_1 _15477_ (.A0(\i_tinyqv.cpu.i_core.mepc[17] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .S(net2219),
    .X(_06923_));
 sg13g2_mux2_1 _15478_ (.A0(_06423_),
    .A1(_06923_),
    .S(net2305),
    .X(_06924_));
 sg13g2_a21oi_1 _15479_ (.A1(net1857),
    .A2(_06924_),
    .Y(_06925_),
    .B1(net1770));
 sg13g2_o21ai_1 _15480_ (.B1(net2484),
    .Y(_06926_),
    .A1(net2411),
    .A2(net1767));
 sg13g2_a21oi_1 _15481_ (.A1(_06922_),
    .A2(_06925_),
    .Y(_00801_),
    .B1(_06926_));
 sg13g2_mux2_1 _15482_ (.A0(\i_tinyqv.cpu.i_core.mepc[18] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .S(net2219),
    .X(_06927_));
 sg13g2_nor2_1 _15483_ (.A(_02236_),
    .B(net1810),
    .Y(_06928_));
 sg13g2_o21ai_1 _15484_ (.B1(net1856),
    .Y(_06929_),
    .A1(net2706),
    .A2(net1807));
 sg13g2_o21ai_1 _15485_ (.B1(net1858),
    .Y(_06930_),
    .A1(net2238),
    .A2(_06927_));
 sg13g2_a21oi_1 _15486_ (.A1(net2239),
    .A2(_06432_),
    .Y(_06931_),
    .B1(_06930_));
 sg13g2_o21ai_1 _15487_ (.B1(net1766),
    .Y(_06932_),
    .A1(_06928_),
    .A2(_06929_));
 sg13g2_o21ai_1 _15488_ (.B1(net2484),
    .Y(_06933_),
    .A1(_06931_),
    .A2(_06932_));
 sg13g2_a21oi_1 _15489_ (.A1(_00977_),
    .A2(net1769),
    .Y(_00802_),
    .B1(_06933_));
 sg13g2_mux2_1 _15490_ (.A0(\i_tinyqv.cpu.i_core.mepc[19] ),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .S(net2219),
    .X(_06934_));
 sg13g2_a21oi_1 _15491_ (.A1(net2305),
    .A2(_06934_),
    .Y(_06935_),
    .B1(net1856));
 sg13g2_o21ai_1 _15492_ (.B1(_06935_),
    .Y(_06936_),
    .A1(net2305),
    .A2(_06442_));
 sg13g2_nand2_1 _15493_ (.Y(_06937_),
    .A(_02337_),
    .B(net1807));
 sg13g2_a21oi_1 _15494_ (.A1(net2701),
    .A2(net1811),
    .Y(_06938_),
    .B1(net1857));
 sg13g2_a21oi_1 _15495_ (.A1(_06937_),
    .A2(_06938_),
    .Y(_06939_),
    .B1(net1769));
 sg13g2_a22oi_1 _15496_ (.Y(_06940_),
    .B1(_06936_),
    .B2(_06939_),
    .A2(net1769),
    .A1(net2410));
 sg13g2_nor2_1 _15497_ (.A(net2341),
    .B(_06940_),
    .Y(_00803_));
 sg13g2_mux2_1 _15498_ (.A0(net2837),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .S(net2219),
    .X(_06941_));
 sg13g2_o21ai_1 _15499_ (.B1(net1857),
    .Y(_06942_),
    .A1(net2238),
    .A2(_06941_));
 sg13g2_a21o_1 _15500_ (.A2(_06449_),
    .A1(net2239),
    .B1(_06942_),
    .X(_06943_));
 sg13g2_a21oi_1 _15501_ (.A1(_01978_),
    .A2(net1808),
    .Y(_06944_),
    .B1(net1860));
 sg13g2_o21ai_1 _15502_ (.B1(_06944_),
    .Y(_06945_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .A2(net1808));
 sg13g2_nand3_1 _15503_ (.B(_06943_),
    .C(_06945_),
    .A(net1767),
    .Y(_06946_));
 sg13g2_o21ai_1 _15504_ (.B1(_06946_),
    .Y(_06947_),
    .A1(net2409),
    .A2(net1767));
 sg13g2_nor2_1 _15505_ (.A(net2341),
    .B(net4146),
    .Y(_00804_));
 sg13g2_mux2_1 _15506_ (.A0(net2861),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .S(net2220),
    .X(_06948_));
 sg13g2_o21ai_1 _15507_ (.B1(net1857),
    .Y(_06949_),
    .A1(net2238),
    .A2(_06948_));
 sg13g2_a21oi_1 _15508_ (.A1(net2239),
    .A2(_06460_),
    .Y(_06950_),
    .B1(_06949_));
 sg13g2_nor2_1 _15509_ (.A(_02160_),
    .B(net1811),
    .Y(_06951_));
 sg13g2_o21ai_1 _15510_ (.B1(net1856),
    .Y(_06952_),
    .A1(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .A2(net1808));
 sg13g2_o21ai_1 _15511_ (.B1(net1767),
    .Y(_06953_),
    .A1(_06951_),
    .A2(_06952_));
 sg13g2_o21ai_1 _15512_ (.B1(net2489),
    .Y(_06954_),
    .A1(_06950_),
    .A2(_06953_));
 sg13g2_a21oi_1 _15513_ (.A1(_00976_),
    .A2(net1770),
    .Y(_00805_),
    .B1(_06954_));
 sg13g2_mux2_1 _15514_ (.A0(net2859),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .S(net2220),
    .X(_06955_));
 sg13g2_o21ai_1 _15515_ (.B1(net1858),
    .Y(_06956_),
    .A1(net2239),
    .A2(_06955_));
 sg13g2_a21oi_1 _15516_ (.A1(net2239),
    .A2(_06471_),
    .Y(_06957_),
    .B1(_06956_));
 sg13g2_a21oi_1 _15517_ (.A1(_02235_),
    .A2(net1809),
    .Y(_06958_),
    .B1(net1861));
 sg13g2_o21ai_1 _15518_ (.B1(_06958_),
    .Y(_06959_),
    .A1(net2741),
    .A2(net1808));
 sg13g2_nand2_1 _15519_ (.Y(_06960_),
    .A(net1768),
    .B(_06959_));
 sg13g2_o21ai_1 _15520_ (.B1(net2489),
    .Y(_06961_),
    .A1(_06957_),
    .A2(_06960_));
 sg13g2_a21oi_1 _15521_ (.A1(_00975_),
    .A2(net1770),
    .Y(_00806_),
    .B1(_06961_));
 sg13g2_mux2_1 _15522_ (.A0(net2828),
    .A1(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .S(net2220),
    .X(_06962_));
 sg13g2_o21ai_1 _15523_ (.B1(net1858),
    .Y(_06963_),
    .A1(net2238),
    .A2(_06962_));
 sg13g2_a21oi_1 _15524_ (.A1(net2239),
    .A2(_06479_),
    .Y(_06964_),
    .B1(_06963_));
 sg13g2_o21ai_1 _15525_ (.B1(net1856),
    .Y(_06965_),
    .A1(net2742),
    .A2(net1808));
 sg13g2_a21oi_1 _15526_ (.A1(_02336_),
    .A2(net1808),
    .Y(_06966_),
    .B1(_06965_));
 sg13g2_nor3_1 _15527_ (.A(net1772),
    .B(_06964_),
    .C(_06966_),
    .Y(_06967_));
 sg13g2_o21ai_1 _15528_ (.B1(net2489),
    .Y(_06968_),
    .A1(net4036),
    .A2(net1767));
 sg13g2_nor2_1 _15529_ (.A(_06967_),
    .B(_06968_),
    .Y(_00807_));
 sg13g2_a21oi_1 _15530_ (.A1(\i_tinyqv.cpu.instr_fetch_running ),
    .A2(_01110_),
    .Y(_06969_),
    .B1(net4057));
 sg13g2_o21ai_1 _15531_ (.B1(net1855),
    .Y(_06970_),
    .A1(_02568_),
    .A2(net4058));
 sg13g2_nand2_1 _15532_ (.Y(_06971_),
    .A(net2491),
    .B(_06970_));
 sg13g2_nor2_1 _15533_ (.A(_02569_),
    .B(_06971_),
    .Y(_00808_));
 sg13g2_nand3_1 _15534_ (.B(net2490),
    .C(net2229),
    .A(net2406),
    .Y(_06972_));
 sg13g2_nand2_1 _15535_ (.Y(_00809_),
    .A(_02567_),
    .B(_06972_));
 sg13g2_nor2_2 _15536_ (.A(net2235),
    .B(net3443),
    .Y(_06973_));
 sg13g2_o21ai_1 _15537_ (.B1(net2497),
    .Y(_06974_),
    .A1(net2399),
    .A2(_06973_));
 sg13g2_a21oi_1 _15538_ (.A1(_02815_),
    .A2(_06973_),
    .Y(_00810_),
    .B1(_06974_));
 sg13g2_o21ai_1 _15539_ (.B1(net2497),
    .Y(_06975_),
    .A1(net2398),
    .A2(_06973_));
 sg13g2_a21oi_1 _15540_ (.A1(_02818_),
    .A2(_06973_),
    .Y(_00811_),
    .B1(_06975_));
 sg13g2_o21ai_1 _15541_ (.B1(net2497),
    .Y(_06976_),
    .A1(net2396),
    .A2(_06973_));
 sg13g2_a21oi_1 _15542_ (.A1(_02820_),
    .A2(_06973_),
    .Y(_00812_),
    .B1(_06976_));
 sg13g2_o21ai_1 _15543_ (.B1(net2497),
    .Y(_06977_),
    .A1(net2394),
    .A2(_06973_));
 sg13g2_a21oi_1 _15544_ (.A1(_02824_),
    .A2(_06973_),
    .Y(_00813_),
    .B1(_06977_));
 sg13g2_nand2_2 _15545_ (.Y(_06978_),
    .A(_01343_),
    .B(net2303));
 sg13g2_nor2_1 _15546_ (.A(net2317),
    .B(_02815_),
    .Y(_06979_));
 sg13g2_and3_2 _15547_ (.X(_06980_),
    .A(net2235),
    .B(net2303),
    .C(_02001_));
 sg13g2_a22oi_1 _15548_ (.Y(_06981_),
    .B1(_06979_),
    .B2(net2150),
    .A2(_06978_),
    .A1(net2392));
 sg13g2_nor2_1 _15549_ (.A(net2345),
    .B(_06981_),
    .Y(_00814_));
 sg13g2_nor2_1 _15550_ (.A(net2317),
    .B(_02818_),
    .Y(_06982_));
 sg13g2_a22oi_1 _15551_ (.Y(_06983_),
    .B1(net2150),
    .B2(_06982_),
    .A2(_06978_),
    .A1(net2390));
 sg13g2_nor2_1 _15552_ (.A(net2345),
    .B(_06983_),
    .Y(_00815_));
 sg13g2_nor2_1 _15553_ (.A(net2317),
    .B(_02820_),
    .Y(_06984_));
 sg13g2_a22oi_1 _15554_ (.Y(_06985_),
    .B1(net2150),
    .B2(_06984_),
    .A2(_06978_),
    .A1(net4082));
 sg13g2_nor2_1 _15555_ (.A(net2347),
    .B(_06985_),
    .Y(_00816_));
 sg13g2_nor2_1 _15556_ (.A(_01197_),
    .B(_02824_),
    .Y(_06986_));
 sg13g2_a22oi_1 _15557_ (.Y(_06987_),
    .B1(net2150),
    .B2(_06986_),
    .A2(_06978_),
    .A1(net4150));
 sg13g2_nor2_1 _15558_ (.A(net2345),
    .B(_06987_),
    .Y(_00817_));
 sg13g2_nand2_2 _15559_ (.Y(_06988_),
    .A(_01265_),
    .B(net2303));
 sg13g2_nor2_1 _15560_ (.A(net2324),
    .B(_02815_),
    .Y(_06989_));
 sg13g2_a22oi_1 _15561_ (.Y(_06990_),
    .B1(_06989_),
    .B2(net2150),
    .A2(_06988_),
    .A1(net4095));
 sg13g2_nor2_1 _15562_ (.A(net2343),
    .B(_06990_),
    .Y(_00818_));
 sg13g2_nor2_1 _15563_ (.A(net2324),
    .B(_02818_),
    .Y(_06991_));
 sg13g2_a22oi_1 _15564_ (.Y(_06992_),
    .B1(_06991_),
    .B2(net2150),
    .A2(_06988_),
    .A1(net4034));
 sg13g2_nor2_1 _15565_ (.A(net2344),
    .B(_06992_),
    .Y(_00819_));
 sg13g2_nor2_1 _15566_ (.A(net2324),
    .B(_02820_),
    .Y(_06993_));
 sg13g2_a22oi_1 _15567_ (.Y(_06994_),
    .B1(_06993_),
    .B2(net2150),
    .A2(_06988_),
    .A1(net4107));
 sg13g2_nor2_1 _15568_ (.A(net2343),
    .B(_06994_),
    .Y(_00820_));
 sg13g2_nor2_1 _15569_ (.A(_01163_),
    .B(_02824_),
    .Y(_06995_));
 sg13g2_a22oi_1 _15570_ (.Y(_06996_),
    .B1(_06995_),
    .B2(net2150),
    .A2(_06988_),
    .A1(net4108));
 sg13g2_nor2_1 _15571_ (.A(net2344),
    .B(_06996_),
    .Y(_00821_));
 sg13g2_nand2_2 _15572_ (.Y(_06997_),
    .A(_01346_),
    .B(net2303));
 sg13g2_nor2_1 _15573_ (.A(net2307),
    .B(_02815_),
    .Y(_06998_));
 sg13g2_a22oi_1 _15574_ (.Y(_06999_),
    .B1(_06998_),
    .B2(net2151),
    .A2(_06997_),
    .A1(net4124));
 sg13g2_nor2_1 _15575_ (.A(net2343),
    .B(_06999_),
    .Y(_00822_));
 sg13g2_nor2_1 _15576_ (.A(net2307),
    .B(_02818_),
    .Y(_07000_));
 sg13g2_a22oi_1 _15577_ (.Y(_07001_),
    .B1(_07000_),
    .B2(net2151),
    .A2(_06997_),
    .A1(net3590));
 sg13g2_nor2_1 _15578_ (.A(net2346),
    .B(_07001_),
    .Y(_00823_));
 sg13g2_nor2_1 _15579_ (.A(net2307),
    .B(_02820_),
    .Y(_07002_));
 sg13g2_a22oi_1 _15580_ (.Y(_07003_),
    .B1(_07002_),
    .B2(net2151),
    .A2(_06997_),
    .A1(net3688));
 sg13g2_nor2_1 _15581_ (.A(net2346),
    .B(_07003_),
    .Y(_00824_));
 sg13g2_nor2_1 _15582_ (.A(_01202_),
    .B(_02824_),
    .Y(_07004_));
 sg13g2_a22oi_1 _15583_ (.Y(_07005_),
    .B1(_07004_),
    .B2(net2151),
    .A2(_06997_),
    .A1(net3435));
 sg13g2_nor2_1 _15584_ (.A(net2343),
    .B(_07005_),
    .Y(_00825_));
 sg13g2_nand2_2 _15585_ (.Y(_07006_),
    .A(_01208_),
    .B(net2303));
 sg13g2_o21ai_1 _15586_ (.B1(net2496),
    .Y(_07007_),
    .A1(_02816_),
    .A2(_07006_));
 sg13g2_a21oi_1 _15587_ (.A1(_00962_),
    .A2(_07006_),
    .Y(_00826_),
    .B1(_07007_));
 sg13g2_o21ai_1 _15588_ (.B1(net2496),
    .Y(_07008_),
    .A1(_02817_),
    .A2(_07006_));
 sg13g2_a21oi_1 _15589_ (.A1(_00961_),
    .A2(_07006_),
    .Y(_00827_),
    .B1(_07008_));
 sg13g2_o21ai_1 _15590_ (.B1(net2496),
    .Y(_07009_),
    .A1(_02821_),
    .A2(_07006_));
 sg13g2_a21oi_1 _15591_ (.A1(_00960_),
    .A2(_07006_),
    .Y(_00828_),
    .B1(_07009_));
 sg13g2_o21ai_1 _15592_ (.B1(net2496),
    .Y(_07010_),
    .A1(_02823_),
    .A2(_07006_));
 sg13g2_a21oi_1 _15593_ (.A1(_00959_),
    .A2(_07006_),
    .Y(_00829_),
    .B1(_07010_));
 sg13g2_nand2_2 _15594_ (.Y(_07011_),
    .A(_01206_),
    .B(net2303));
 sg13g2_a21oi_2 _15595_ (.B1(_01405_),
    .Y(_07012_),
    .A2(_02001_),
    .A1(net2235));
 sg13g2_a22oi_1 _15596_ (.Y(_07013_),
    .B1(net2148),
    .B2(_06979_),
    .A2(_07011_),
    .A1(net4035));
 sg13g2_nor2_1 _15597_ (.A(net2345),
    .B(_07013_),
    .Y(_00830_));
 sg13g2_a22oi_1 _15598_ (.Y(_07014_),
    .B1(net2148),
    .B2(_06982_),
    .A2(_07011_),
    .A1(net3642));
 sg13g2_nor2_1 _15599_ (.A(net2345),
    .B(_07014_),
    .Y(_00831_));
 sg13g2_a22oi_1 _15600_ (.Y(_07015_),
    .B1(net2148),
    .B2(_06984_),
    .A2(_07011_),
    .A1(net3643));
 sg13g2_nor2_1 _15601_ (.A(net2347),
    .B(_07015_),
    .Y(_00832_));
 sg13g2_a22oi_1 _15602_ (.Y(_07016_),
    .B1(net2148),
    .B2(_06986_),
    .A2(_07011_),
    .A1(net3591));
 sg13g2_nor2_1 _15603_ (.A(net2345),
    .B(_07016_),
    .Y(_00833_));
 sg13g2_nand2_2 _15604_ (.Y(_07017_),
    .A(_01164_),
    .B(_01404_));
 sg13g2_a22oi_1 _15605_ (.Y(_07018_),
    .B1(_07017_),
    .B2(net3225),
    .A2(net2148),
    .A1(_06989_));
 sg13g2_nor2_1 _15606_ (.A(net2344),
    .B(_07018_),
    .Y(_00834_));
 sg13g2_a22oi_1 _15607_ (.Y(_07019_),
    .B1(_07017_),
    .B2(net3196),
    .A2(net2148),
    .A1(_06991_));
 sg13g2_nor2_1 _15608_ (.A(net2344),
    .B(_07019_),
    .Y(_00835_));
 sg13g2_a22oi_1 _15609_ (.Y(_07020_),
    .B1(_07017_),
    .B2(net3329),
    .A2(net2148),
    .A1(_06993_));
 sg13g2_nor2_1 _15610_ (.A(net2344),
    .B(_07020_),
    .Y(_00836_));
 sg13g2_a22oi_1 _15611_ (.Y(_07021_),
    .B1(_07017_),
    .B2(net3386),
    .A2(net2148),
    .A1(_06995_));
 sg13g2_nor2_1 _15612_ (.A(net2344),
    .B(_07021_),
    .Y(_00837_));
 sg13g2_nand2_2 _15613_ (.Y(_07022_),
    .A(_01385_),
    .B(_01404_));
 sg13g2_a22oi_1 _15614_ (.Y(_07023_),
    .B1(_07022_),
    .B2(net3229),
    .A2(net2149),
    .A1(_06998_));
 sg13g2_nor2_1 _15615_ (.A(net2343),
    .B(_07023_),
    .Y(_00838_));
 sg13g2_a22oi_1 _15616_ (.Y(_07024_),
    .B1(_07022_),
    .B2(net3317),
    .A2(net2149),
    .A1(_07000_));
 sg13g2_nor2_1 _15617_ (.A(net2343),
    .B(_07024_),
    .Y(_00839_));
 sg13g2_a22oi_1 _15618_ (.Y(_07025_),
    .B1(_07022_),
    .B2(net3327),
    .A2(net2149),
    .A1(_07002_));
 sg13g2_nor2_1 _15619_ (.A(net2343),
    .B(_07025_),
    .Y(_00840_));
 sg13g2_a22oi_1 _15620_ (.Y(_07026_),
    .B1(_07022_),
    .B2(net3281),
    .A2(net2149),
    .A1(_07004_));
 sg13g2_nor2_1 _15621_ (.A(net2343),
    .B(_07026_),
    .Y(_00841_));
 sg13g2_a21oi_1 _15622_ (.A1(net3732),
    .A2(net2232),
    .Y(_07027_),
    .B1(_01944_));
 sg13g2_nand2_1 _15623_ (.Y(_07028_),
    .A(_02635_),
    .B(_07027_));
 sg13g2_nor2_1 _15624_ (.A(net4051),
    .B(_07028_),
    .Y(_07029_));
 sg13g2_nor2_1 _15625_ (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .B(_02635_),
    .Y(_07030_));
 sg13g2_o21ai_1 _15626_ (.B1(net2494),
    .Y(_00842_),
    .A1(_07029_),
    .A2(_07030_));
 sg13g2_nor2_1 _15627_ (.A(\i_tinyqv.cpu.data_write_n[1] ),
    .B(_07028_),
    .Y(_07031_));
 sg13g2_nor2_1 _15628_ (.A(net4049),
    .B(_02635_),
    .Y(_07032_));
 sg13g2_o21ai_1 _15629_ (.B1(net2494),
    .Y(_00843_),
    .A1(_07031_),
    .A2(_07032_));
 sg13g2_a21oi_1 _15630_ (.A1(net2775),
    .A2(_01944_),
    .Y(_07033_),
    .B1(_02628_));
 sg13g2_nor2_1 _15631_ (.A(net3798),
    .B(net2123),
    .Y(_07034_));
 sg13g2_nor2_1 _15632_ (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .B(net2122),
    .Y(_07035_));
 sg13g2_o21ai_1 _15633_ (.B1(_07033_),
    .Y(_00844_),
    .A1(_07034_),
    .A2(_07035_));
 sg13g2_nor2_1 _15634_ (.A(net3800),
    .B(net2123),
    .Y(_07036_));
 sg13g2_nor2_1 _15635_ (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .B(net2122),
    .Y(_07037_));
 sg13g2_o21ai_1 _15636_ (.B1(_07033_),
    .Y(_00845_),
    .A1(_07036_),
    .A2(_07037_));
 sg13g2_nor4_1 _15637_ (.A(net3732),
    .B(_01907_),
    .C(_01944_),
    .D(_02634_),
    .Y(_07038_));
 sg13g2_a21oi_1 _15638_ (.A1(net4041),
    .A2(net2223),
    .Y(_07039_),
    .B1(_02635_));
 sg13g2_nor3_1 _15639_ (.A(net2229),
    .B(_07038_),
    .C(_07039_),
    .Y(_07040_));
 sg13g2_a21oi_1 _15640_ (.A1(net3713),
    .A2(net2229),
    .Y(_07041_),
    .B1(_07040_));
 sg13g2_nand2_1 _15641_ (.Y(_00846_),
    .A(net2494),
    .B(_07041_));
 sg13g2_a21oi_1 _15642_ (.A1(_00945_),
    .A2(_02632_),
    .Y(_00847_),
    .B1(_02628_));
 sg13g2_o21ai_1 _15643_ (.B1(net2489),
    .Y(_07042_),
    .A1(net3852),
    .A2(net2125));
 sg13g2_and2_1 _15644_ (.A(net3540),
    .B(net2222),
    .X(_07043_));
 sg13g2_a21oi_1 _15645_ (.A1(\i_tinyqv.cpu.i_core.mepc[0] ),
    .A2(net2186),
    .Y(_07044_),
    .B1(_07043_));
 sg13g2_a21oi_1 _15646_ (.A1(net2125),
    .A2(_07044_),
    .Y(_00848_),
    .B1(_07042_));
 sg13g2_o21ai_1 _15647_ (.B1(net2489),
    .Y(_07045_),
    .A1(net2122),
    .A2(_06271_));
 sg13g2_a21oi_1 _15648_ (.A1(_00944_),
    .A2(net2122),
    .Y(_00849_),
    .B1(_07045_));
 sg13g2_nand2_1 _15649_ (.Y(_07046_),
    .A(net3916),
    .B(_06276_));
 sg13g2_xnor2_1 _15650_ (.Y(_07047_),
    .A(net3916),
    .B(_06276_));
 sg13g2_o21ai_1 _15651_ (.B1(net2490),
    .Y(_07048_),
    .A1(net2388),
    .A2(net2123));
 sg13g2_a21oi_1 _15652_ (.A1(net2123),
    .A2(_07047_),
    .Y(_00850_),
    .B1(_07048_));
 sg13g2_xor2_1 _15653_ (.B(_06822_),
    .A(net2801),
    .X(_07049_));
 sg13g2_o21ai_1 _15654_ (.B1(net2123),
    .Y(_07050_),
    .A1(_07046_),
    .A2(_07049_));
 sg13g2_a21oi_1 _15655_ (.A1(_07046_),
    .A2(_07049_),
    .Y(_07051_),
    .B1(_07050_));
 sg13g2_o21ai_1 _15656_ (.B1(net2491),
    .Y(_07052_),
    .A1(net3975),
    .A2(net2123));
 sg13g2_nor2_1 _15657_ (.A(_07051_),
    .B(_07052_),
    .Y(_00851_));
 sg13g2_o21ai_1 _15658_ (.B1(net2489),
    .Y(_07053_),
    .A1(net2385),
    .A2(net2124));
 sg13g2_a21oi_1 _15659_ (.A1(net2124),
    .A2(_06829_),
    .Y(_00852_),
    .B1(_07053_));
 sg13g2_o21ai_1 _15660_ (.B1(net2491),
    .Y(_07054_),
    .A1(net4061),
    .A2(net2124));
 sg13g2_a21oi_1 _15661_ (.A1(net2124),
    .A2(_06838_),
    .Y(_00853_),
    .B1(_07054_));
 sg13g2_o21ai_1 _15662_ (.B1(net2491),
    .Y(_07055_),
    .A1(net2122),
    .A2(_06845_));
 sg13g2_a21oi_1 _15663_ (.A1(_00942_),
    .A2(net2122),
    .Y(_00854_),
    .B1(_07055_));
 sg13g2_o21ai_1 _15664_ (.B1(net2489),
    .Y(_07056_),
    .A1(net2122),
    .A2(_06853_));
 sg13g2_a21oi_1 _15665_ (.A1(_00941_),
    .A2(net2122),
    .Y(_00855_),
    .B1(_07056_));
 sg13g2_o21ai_1 _15666_ (.B1(net2483),
    .Y(_07057_),
    .A1(net4044),
    .A2(net2125));
 sg13g2_a21oi_1 _15667_ (.A1(net2125),
    .A2(_06860_),
    .Y(_00856_),
    .B1(_07057_));
 sg13g2_o21ai_1 _15668_ (.B1(net2489),
    .Y(_07058_),
    .A1(net3960),
    .A2(net2124));
 sg13g2_a21oi_1 _15669_ (.A1(net2124),
    .A2(_06868_),
    .Y(_00857_),
    .B1(_07058_));
 sg13g2_o21ai_1 _15670_ (.B1(net2484),
    .Y(_07059_),
    .A1(net2120),
    .A2(_06876_));
 sg13g2_a21oi_1 _15671_ (.A1(_00940_),
    .A2(net2120),
    .Y(_00858_),
    .B1(_07059_));
 sg13g2_o21ai_1 _15672_ (.B1(net2483),
    .Y(_07060_),
    .A1(net4005),
    .A2(net2125));
 sg13g2_a21oi_1 _15673_ (.A1(net2125),
    .A2(_06881_),
    .Y(_00859_),
    .B1(_07060_));
 sg13g2_o21ai_1 _15674_ (.B1(net2482),
    .Y(_07061_),
    .A1(net2117),
    .A2(_06890_));
 sg13g2_a21oi_1 _15675_ (.A1(_00939_),
    .A2(net2118),
    .Y(_00860_),
    .B1(_07061_));
 sg13g2_o21ai_1 _15676_ (.B1(net2483),
    .Y(_07062_),
    .A1(net2116),
    .A2(_06895_));
 sg13g2_a21oi_1 _15677_ (.A1(_00938_),
    .A2(net2118),
    .Y(_00861_),
    .B1(_07062_));
 sg13g2_o21ai_1 _15678_ (.B1(net2482),
    .Y(_07063_),
    .A1(net2116),
    .A2(_06904_));
 sg13g2_a21oi_1 _15679_ (.A1(_00937_),
    .A2(net2116),
    .Y(_00862_),
    .B1(_07063_));
 sg13g2_o21ai_1 _15680_ (.B1(net2482),
    .Y(_07064_),
    .A1(net2116),
    .A2(_06911_));
 sg13g2_a21oi_1 _15681_ (.A1(_00936_),
    .A2(net2116),
    .Y(_00863_),
    .B1(_07064_));
 sg13g2_o21ai_1 _15682_ (.B1(net2482),
    .Y(_07065_),
    .A1(net2119),
    .A2(_06916_));
 sg13g2_a21oi_1 _15683_ (.A1(_00935_),
    .A2(net2119),
    .Y(_00864_),
    .B1(_07065_));
 sg13g2_o21ai_1 _15684_ (.B1(net2482),
    .Y(_07066_),
    .A1(net2116),
    .A2(_06923_));
 sg13g2_a21oi_1 _15685_ (.A1(_00934_),
    .A2(net2117),
    .Y(_00865_),
    .B1(_07066_));
 sg13g2_o21ai_1 _15686_ (.B1(net2483),
    .Y(_07067_),
    .A1(net2116),
    .A2(_06927_));
 sg13g2_a21oi_1 _15687_ (.A1(_00933_),
    .A2(net2118),
    .Y(_00866_),
    .B1(_07067_));
 sg13g2_o21ai_1 _15688_ (.B1(net2482),
    .Y(_07068_),
    .A1(net2116),
    .A2(_06934_));
 sg13g2_a21oi_1 _15689_ (.A1(_00932_),
    .A2(net2117),
    .Y(_00867_),
    .B1(_07068_));
 sg13g2_o21ai_1 _15690_ (.B1(net2482),
    .Y(_07069_),
    .A1(net2117),
    .A2(_06941_));
 sg13g2_a21oi_1 _15691_ (.A1(_00931_),
    .A2(net2118),
    .Y(_00868_),
    .B1(_07069_));
 sg13g2_o21ai_1 _15692_ (.B1(net2482),
    .Y(_07070_),
    .A1(net2117),
    .A2(_06948_));
 sg13g2_a21oi_1 _15693_ (.A1(_00930_),
    .A2(net2118),
    .Y(_00869_),
    .B1(_07070_));
 sg13g2_o21ai_1 _15694_ (.B1(net2485),
    .Y(_07071_),
    .A1(net2120),
    .A2(_06955_));
 sg13g2_a21oi_1 _15695_ (.A1(_00929_),
    .A2(net2120),
    .Y(_00870_),
    .B1(_07071_));
 sg13g2_o21ai_1 _15696_ (.B1(net2485),
    .Y(_07072_),
    .A1(net2120),
    .A2(_06962_));
 sg13g2_a21oi_1 _15697_ (.A1(_00928_),
    .A2(net2120),
    .Y(_00871_),
    .B1(_07072_));
 sg13g2_nor2_1 _15698_ (.A(net2186),
    .B(net2121),
    .Y(_07073_));
 sg13g2_a22oi_1 _15699_ (.Y(_07074_),
    .B1(_07073_),
    .B2(net3651),
    .A2(net2120),
    .A1(net3789));
 sg13g2_nor2_1 _15700_ (.A(net2341),
    .B(_07074_),
    .Y(_00872_));
 sg13g2_a22oi_1 _15701_ (.Y(_07075_),
    .B1(_07073_),
    .B2(net3697),
    .A2(net2120),
    .A1(net3940));
 sg13g2_nor2_1 _15702_ (.A(net2341),
    .B(_07075_),
    .Y(_00873_));
 sg13g2_a22oi_1 _15703_ (.Y(_07076_),
    .B1(_07073_),
    .B2(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .A2(net2121),
    .A1(net4013));
 sg13g2_nor2_1 _15704_ (.A(net2341),
    .B(net4014),
    .Y(_00874_));
 sg13g2_a21oi_1 _15705_ (.A1(net4041),
    .A2(net2220),
    .Y(_07077_),
    .B1(net2119));
 sg13g2_o21ai_1 _15706_ (.B1(net2483),
    .Y(_07078_),
    .A1(net4085),
    .A2(net2125));
 sg13g2_nor2_1 _15707_ (.A(_07077_),
    .B(_07078_),
    .Y(_00875_));
 sg13g2_nor2_1 _15708_ (.A(net2341),
    .B(net2383),
    .Y(_00876_));
 sg13g2_nor3_1 _15709_ (.A(net2342),
    .B(net2315),
    .C(net2309),
    .Y(_00877_));
 sg13g2_nor2_1 _15710_ (.A(net2377),
    .B(net2312),
    .Y(_07079_));
 sg13g2_nor3_1 _15711_ (.A(net2347),
    .B(net2232),
    .C(_07079_),
    .Y(_00878_));
 sg13g2_nor3_1 _15712_ (.A(net2341),
    .B(_01957_),
    .C(_01958_),
    .Y(_00879_));
 sg13g2_nor2_2 _15713_ (.A(net2066),
    .B(net1814),
    .Y(_07080_));
 sg13g2_a22oi_1 _15714_ (.Y(_07081_),
    .B1(_06080_),
    .B2(_02778_),
    .A2(_06065_),
    .A1(_06062_));
 sg13g2_nor2_1 _15715_ (.A(_06044_),
    .B(_07081_),
    .Y(_07082_));
 sg13g2_a221oi_1 _15716_ (.B2(_02544_),
    .C1(_07082_),
    .B1(_07080_),
    .A1(net4144),
    .Y(_07083_),
    .A2(net1815));
 sg13g2_nor2_1 _15717_ (.A(net2348),
    .B(_07083_),
    .Y(_00880_));
 sg13g2_nor2b_1 _15718_ (.A(net2127),
    .B_N(_06066_),
    .Y(_07084_));
 sg13g2_nand2b_1 _15719_ (.Y(_07085_),
    .B(_06066_),
    .A_N(net2127));
 sg13g2_nand3b_1 _15720_ (.B(_02537_),
    .C(net2138),
    .Y(_07086_),
    .A_N(net2136));
 sg13g2_nor2_1 _15721_ (.A(net2066),
    .B(_07086_),
    .Y(_07087_));
 sg13g2_a22oi_1 _15722_ (.Y(_07088_),
    .B1(_07087_),
    .B2(_02542_),
    .A2(_07085_),
    .A1(_02771_));
 sg13g2_nor3_1 _15723_ (.A(_02753_),
    .B(_02757_),
    .C(_06120_),
    .Y(_07089_));
 sg13g2_nand3_1 _15724_ (.B(_07088_),
    .C(_07089_),
    .A(net1817),
    .Y(_07090_));
 sg13g2_o21ai_1 _15725_ (.B1(_07090_),
    .Y(_07091_),
    .A1(net3825),
    .A2(net1816));
 sg13g2_nor2_1 _15726_ (.A(net2348),
    .B(_07091_),
    .Y(_00881_));
 sg13g2_nor2_1 _15727_ (.A(net2134),
    .B(net1972),
    .Y(_07092_));
 sg13g2_a22oi_1 _15728_ (.Y(_07093_),
    .B1(_07080_),
    .B2(_07092_),
    .A2(net1814),
    .A1(net3700));
 sg13g2_nor2_1 _15729_ (.A(net2348),
    .B(_07093_),
    .Y(_00882_));
 sg13g2_nor2_1 _15730_ (.A(net2066),
    .B(_06051_),
    .Y(_07094_));
 sg13g2_a221oi_1 _15731_ (.B2(_02538_),
    .C1(_06078_),
    .B1(_07094_),
    .A1(_06062_),
    .Y(_07095_),
    .A2(_06064_));
 sg13g2_nand3_1 _15732_ (.B(net2493),
    .C(net1814),
    .A(net3442),
    .Y(_07096_));
 sg13g2_o21ai_1 _15733_ (.B1(_07096_),
    .Y(_00883_),
    .A1(net1782),
    .A2(_07095_));
 sg13g2_nor2_1 _15734_ (.A(_06051_),
    .B(_07086_),
    .Y(_07097_));
 sg13g2_o21ai_1 _15735_ (.B1(_02765_),
    .Y(_07098_),
    .A1(_02533_),
    .A2(_02544_));
 sg13g2_a221oi_1 _15736_ (.B2(net2068),
    .C1(_07098_),
    .B1(_07097_),
    .A1(_02771_),
    .Y(_07099_),
    .A2(_07084_));
 sg13g2_nand3_1 _15737_ (.B(net2492),
    .C(net1815),
    .A(net3062),
    .Y(_07100_));
 sg13g2_o21ai_1 _15738_ (.B1(_07100_),
    .Y(_00884_),
    .A1(net1782),
    .A2(_07099_));
 sg13g2_nor3_1 _15739_ (.A(net2066),
    .B(_06047_),
    .C(_06051_),
    .Y(_07101_));
 sg13g2_nor3_1 _15740_ (.A(net1814),
    .B(_06181_),
    .C(_07101_),
    .Y(_07102_));
 sg13g2_o21ai_1 _15741_ (.B1(net2492),
    .Y(_07103_),
    .A1(net3824),
    .A2(net1818));
 sg13g2_nor2_1 _15742_ (.A(_07102_),
    .B(_07103_),
    .Y(_00885_));
 sg13g2_or4_1 _15743_ (.A(net2066),
    .B(_02543_),
    .C(_02564_),
    .D(_07092_),
    .X(_07104_));
 sg13g2_o21ai_1 _15744_ (.B1(net1940),
    .Y(_07105_),
    .A1(net2066),
    .A2(_06170_));
 sg13g2_o21ai_1 _15745_ (.B1(net2493),
    .Y(_07106_),
    .A1(net1815),
    .A2(_07105_));
 sg13g2_a21oi_1 _15746_ (.A1(_00927_),
    .A2(net1815),
    .Y(_00886_),
    .B1(_07106_));
 sg13g2_nand3b_1 _15747_ (.B(_02564_),
    .C(_07080_),
    .Y(_07107_),
    .A_N(net2136));
 sg13g2_nor3_1 _15748_ (.A(_02546_),
    .B(net1814),
    .C(_06071_),
    .Y(_07108_));
 sg13g2_a21oi_1 _15749_ (.A1(net4008),
    .A2(net1814),
    .Y(_07109_),
    .B1(_07108_));
 sg13g2_a21oi_1 _15750_ (.A1(_07107_),
    .A2(_07109_),
    .Y(_00887_),
    .B1(net2348));
 sg13g2_o21ai_1 _15751_ (.B1(net2488),
    .Y(_07110_),
    .A1(_02566_),
    .A2(net1815));
 sg13g2_a21oi_1 _15752_ (.A1(_00925_),
    .A2(net1815),
    .Y(_00888_),
    .B1(_07110_));
 sg13g2_nor3_1 _15753_ (.A(net2066),
    .B(_02563_),
    .C(_07086_),
    .Y(_07111_));
 sg13g2_a221oi_1 _15754_ (.B2(_02498_),
    .C1(_07111_),
    .B1(_06090_),
    .A1(_02545_),
    .Y(_07112_),
    .A2(_06071_));
 sg13g2_o21ai_1 _15755_ (.B1(net2493),
    .Y(_07113_),
    .A1(net3843),
    .A2(net1817));
 sg13g2_a21oi_1 _15756_ (.A1(net1817),
    .A2(_07112_),
    .Y(_00889_),
    .B1(_07113_));
 sg13g2_nor2_1 _15757_ (.A(net3558),
    .B(net1816),
    .Y(_07114_));
 sg13g2_nor3_1 _15758_ (.A(net2348),
    .B(_07080_),
    .C(_07114_),
    .Y(_00890_));
 sg13g2_nand2_1 _15759_ (.Y(_07115_),
    .A(net3819),
    .B(net1814));
 sg13g2_nand3b_1 _15760_ (.B(_07115_),
    .C(net2494),
    .Y(_00891_),
    .A_N(_07080_));
 sg13g2_nand2_2 _15761_ (.Y(_07116_),
    .A(_06142_),
    .B(_07097_));
 sg13g2_nand2_1 _15762_ (.Y(_07117_),
    .A(_06170_),
    .B(_07116_));
 sg13g2_nor2_1 _15763_ (.A(net2127),
    .B(_07117_),
    .Y(_07118_));
 sg13g2_a21oi_1 _15764_ (.A1(_06170_),
    .A2(_07116_),
    .Y(_07119_),
    .B1(net2141));
 sg13g2_nor3_1 _15765_ (.A(_07104_),
    .B(_07118_),
    .C(_07119_),
    .Y(_07120_));
 sg13g2_o21ai_1 _15766_ (.B1(_02771_),
    .Y(_07121_),
    .A1(_06047_),
    .A2(_06067_));
 sg13g2_a21oi_1 _15767_ (.A1(_02563_),
    .A2(_07084_),
    .Y(_07122_),
    .B1(_07121_));
 sg13g2_nor3_1 _15768_ (.A(_02758_),
    .B(_07120_),
    .C(_07122_),
    .Y(_07123_));
 sg13g2_o21ai_1 _15769_ (.B1(net2492),
    .Y(_07124_),
    .A1(net3926),
    .A2(net1816));
 sg13g2_a21oi_1 _15770_ (.A1(net1816),
    .A2(_07123_),
    .Y(_00892_),
    .B1(_07124_));
 sg13g2_a21oi_1 _15771_ (.A1(_02525_),
    .A2(_06169_),
    .Y(_07125_),
    .B1(_07104_));
 sg13g2_o21ai_1 _15772_ (.B1(_07125_),
    .Y(_07126_),
    .A1(net2141),
    .A2(_07117_));
 sg13g2_o21ai_1 _15773_ (.B1(_06064_),
    .Y(_07127_),
    .A1(net2131),
    .A2(_07085_));
 sg13g2_o21ai_1 _15774_ (.B1(_07126_),
    .Y(_07128_),
    .A1(_07121_),
    .A2(_07127_));
 sg13g2_nor3_1 _15775_ (.A(_02764_),
    .B(net1814),
    .C(_07128_),
    .Y(_07129_));
 sg13g2_o21ai_1 _15776_ (.B1(net2493),
    .Y(_07130_),
    .A1(net2372),
    .A2(net1816));
 sg13g2_nor2_1 _15777_ (.A(_07129_),
    .B(_07130_),
    .Y(_00893_));
 sg13g2_nand2_1 _15778_ (.Y(_07131_),
    .A(_02525_),
    .B(_07116_));
 sg13g2_o21ai_1 _15779_ (.B1(_07131_),
    .Y(_07132_),
    .A1(_06147_),
    .A2(_07116_));
 sg13g2_nor3_1 _15780_ (.A(_06169_),
    .B(_07104_),
    .C(_07132_),
    .Y(_07133_));
 sg13g2_nand3_1 _15781_ (.B(_06169_),
    .C(_07132_),
    .A(net2068),
    .Y(_07134_));
 sg13g2_nand2_1 _15782_ (.Y(_07135_),
    .A(_02542_),
    .B(_07084_));
 sg13g2_a21oi_1 _15783_ (.A1(_02771_),
    .A2(_07135_),
    .Y(_07136_),
    .B1(_07133_));
 sg13g2_nand4_1 _15784_ (.B(net1940),
    .C(_07134_),
    .A(net1817),
    .Y(_07137_),
    .D(_07136_));
 sg13g2_o21ai_1 _15785_ (.B1(_07137_),
    .Y(_07138_),
    .A1(net2369),
    .A2(net1818));
 sg13g2_nor2_1 _15786_ (.A(net2339),
    .B(_07138_),
    .Y(_00894_));
 sg13g2_nor2b_1 _15787_ (.A(net2141),
    .B_N(net2126),
    .Y(_07139_));
 sg13g2_o21ai_1 _15788_ (.B1(_06160_),
    .Y(_07140_),
    .A1(net2135),
    .A2(_07139_));
 sg13g2_a221oi_1 _15789_ (.B2(_07140_),
    .C1(_07104_),
    .B1(_07116_),
    .A1(net2131),
    .Y(_07141_),
    .A2(_06052_));
 sg13g2_nand2_1 _15790_ (.Y(_07142_),
    .A(net2130),
    .B(_06065_));
 sg13g2_a21oi_1 _15791_ (.A1(_07135_),
    .A2(_07142_),
    .Y(_07143_),
    .B1(_02772_));
 sg13g2_nor3_2 _15792_ (.A(_02764_),
    .B(_07141_),
    .C(_07143_),
    .Y(_07144_));
 sg13g2_o21ai_1 _15793_ (.B1(net2488),
    .Y(_07145_),
    .A1(net4024),
    .A2(net1818));
 sg13g2_a21oi_1 _15794_ (.A1(net1818),
    .A2(_07144_),
    .Y(_00895_),
    .B1(_07145_));
 sg13g2_nand2_1 _15795_ (.Y(_07146_),
    .A(net3689),
    .B(net2123));
 sg13g2_and4_1 _15796_ (.A(net2490),
    .B(net2234),
    .C(_01945_),
    .D(_07146_),
    .X(_00896_));
 sg13g2_a21oi_2 _15797_ (.B1(_06078_),
    .Y(_07147_),
    .A2(_06080_),
    .A1(_02778_));
 sg13g2_and3_1 _15798_ (.X(_07148_),
    .A(net1940),
    .B(_06267_),
    .C(_07147_));
 sg13g2_nand2_1 _15799_ (.Y(_07149_),
    .A(net2141),
    .B(_02543_));
 sg13g2_nor2b_1 _15800_ (.A(_07149_),
    .B_N(net2128),
    .Y(_07150_));
 sg13g2_a221oi_1 _15801_ (.B2(_07149_),
    .C1(_07148_),
    .B1(_06184_),
    .A1(_02760_),
    .Y(_07151_),
    .A2(_02770_));
 sg13g2_mux2_1 _15802_ (.A0(_00946_),
    .A1(_07151_),
    .S(net1784),
    .X(_07152_));
 sg13g2_inv_1 _15803_ (.Y(_00897_),
    .A(_07152_));
 sg13g2_nand3b_1 _15804_ (.B(_07147_),
    .C(net1790),
    .Y(_07153_),
    .A_N(_06187_));
 sg13g2_o21ai_1 _15805_ (.B1(_07153_),
    .Y(_07154_),
    .A1(net4049),
    .A2(net1790));
 sg13g2_inv_1 _15806_ (.Y(_00898_),
    .A(_07154_));
 sg13g2_a21oi_1 _15807_ (.A1(net2131),
    .A2(net2130),
    .Y(_07155_),
    .B1(_06064_));
 sg13g2_nand4_1 _15808_ (.B(net1940),
    .C(_07147_),
    .A(net2064),
    .Y(_07156_),
    .D(_07155_));
 sg13g2_nor3_1 _15809_ (.A(net2128),
    .B(_02761_),
    .C(_06054_),
    .Y(_07157_));
 sg13g2_nor2_1 _15810_ (.A(_07150_),
    .B(_07157_),
    .Y(_07158_));
 sg13g2_nand3_1 _15811_ (.B(net2140),
    .C(_07158_),
    .A(net2069),
    .Y(_07159_));
 sg13g2_nand3_1 _15812_ (.B(_07156_),
    .C(_07159_),
    .A(net1790),
    .Y(_07160_));
 sg13g2_o21ai_1 _15813_ (.B1(_07160_),
    .Y(_07161_),
    .A1(net3964),
    .A2(net1790));
 sg13g2_inv_1 _15814_ (.Y(_00899_),
    .A(_07161_));
 sg13g2_nand2_1 _15815_ (.Y(_07162_),
    .A(net3866),
    .B(net1783));
 sg13g2_a21o_1 _15816_ (.A2(_02770_),
    .A1(_02559_),
    .B1(_06088_),
    .X(_07163_));
 sg13g2_a221oi_1 _15817_ (.B2(net2143),
    .C1(_02764_),
    .B1(_02757_),
    .A1(_02526_),
    .Y(_07164_),
    .A2(_02752_));
 sg13g2_o21ai_1 _15818_ (.B1(_02532_),
    .Y(_07165_),
    .A1(_02544_),
    .A2(net2128));
 sg13g2_nand3b_1 _15819_ (.B(_07164_),
    .C(_07165_),
    .Y(_07166_),
    .A_N(_07163_));
 sg13g2_nand2_1 _15820_ (.Y(_07167_),
    .A(_02775_),
    .B(_06082_));
 sg13g2_a221oi_1 _15821_ (.B2(_07166_),
    .C1(_07167_),
    .B1(_02551_),
    .A1(net2069),
    .Y(_07168_),
    .A2(_02528_));
 sg13g2_o21ai_1 _15822_ (.B1(_07162_),
    .Y(_00900_),
    .A1(net1783),
    .A2(_07168_));
 sg13g2_a21o_1 _15823_ (.A2(_06085_),
    .A1(_02766_),
    .B1(net2142),
    .X(_07169_));
 sg13g2_nand4_1 _15824_ (.B(_02762_),
    .C(_02775_),
    .A(net2065),
    .Y(_07170_),
    .D(_06084_));
 sg13g2_a21oi_1 _15825_ (.A1(net2129),
    .A2(_07166_),
    .Y(_07171_),
    .B1(_07170_));
 sg13g2_a221oi_1 _15826_ (.B2(_07171_),
    .C1(net1780),
    .B1(_07169_),
    .A1(net2069),
    .Y(_07172_),
    .A2(_06200_));
 sg13g2_a21o_1 _15827_ (.A2(net1783),
    .A1(net3970),
    .B1(_07172_),
    .X(_00901_));
 sg13g2_a22oi_1 _15828_ (.Y(_07173_),
    .B1(_07166_),
    .B2(_02548_),
    .A2(_02760_),
    .A1(net2144));
 sg13g2_nor2_1 _15829_ (.A(net2069),
    .B(_07173_),
    .Y(_07174_));
 sg13g2_nor2_1 _15830_ (.A(_06211_),
    .B(_07174_),
    .Y(_07175_));
 sg13g2_nor2_1 _15831_ (.A(net3914),
    .B(net1793),
    .Y(_07176_));
 sg13g2_a21oi_1 _15832_ (.A1(net1793),
    .A2(_07175_),
    .Y(_00902_),
    .B1(_07176_));
 sg13g2_o21ai_1 _15833_ (.B1(_07166_),
    .Y(_07177_),
    .A1(net2130),
    .A2(_07163_));
 sg13g2_nand3_1 _15834_ (.B(_06218_),
    .C(_07177_),
    .A(net1791),
    .Y(_07178_));
 sg13g2_o21ai_1 _15835_ (.B1(_07178_),
    .Y(_07179_),
    .A1(net4075),
    .A2(net1793));
 sg13g2_inv_1 _15836_ (.Y(_00903_),
    .A(_07179_));
 sg13g2_a21oi_1 _15837_ (.A1(_02782_),
    .A2(net1940),
    .Y(_07180_),
    .B1(_06229_));
 sg13g2_a21oi_1 _15838_ (.A1(_06082_),
    .A2(_07180_),
    .Y(_07181_),
    .B1(net1850));
 sg13g2_xor2_1 _15839_ (.B(net3699),
    .A(net2361),
    .X(_07182_));
 sg13g2_a21oi_1 _15840_ (.A1(net1850),
    .A2(_07182_),
    .Y(_07183_),
    .B1(_07181_));
 sg13g2_nand2_1 _15841_ (.Y(_07184_),
    .A(net2361),
    .B(net1805));
 sg13g2_o21ai_1 _15842_ (.B1(_07184_),
    .Y(_00904_),
    .A1(net1805),
    .A2(_07183_));
 sg13g2_nand3_1 _15843_ (.B(net1940),
    .C(_06082_),
    .A(_02531_),
    .Y(_07185_));
 sg13g2_a21oi_1 _15844_ (.A1(net1940),
    .A2(_06082_),
    .Y(_07186_),
    .B1(net2144));
 sg13g2_o21ai_1 _15845_ (.B1(_06232_),
    .Y(_07187_),
    .A1(_02787_),
    .A2(_07186_));
 sg13g2_nand3_1 _15846_ (.B(net2361),
    .C(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A(net2360),
    .Y(_07188_));
 sg13g2_a21o_1 _15847_ (.A2(\i_tinyqv.cpu.mem_op_increment_reg ),
    .A1(net2361),
    .B1(net2360),
    .X(_07189_));
 sg13g2_a21o_1 _15848_ (.A2(_07189_),
    .A1(_07188_),
    .B1(_02480_),
    .X(_07190_));
 sg13g2_o21ai_1 _15849_ (.B1(_07190_),
    .Y(_07191_),
    .A1(net1851),
    .A2(_07187_));
 sg13g2_nand2_1 _15850_ (.Y(_07192_),
    .A(net2360),
    .B(net1805));
 sg13g2_o21ai_1 _15851_ (.B1(_07192_),
    .Y(_00905_),
    .A1(net1805),
    .A2(_07191_));
 sg13g2_nand4_1 _15852_ (.B(net2360),
    .C(net2361),
    .A(net2359),
    .Y(_07193_),
    .D(net3699));
 sg13g2_nand2b_1 _15853_ (.Y(_07194_),
    .B(_07188_),
    .A_N(net2359));
 sg13g2_a21o_1 _15854_ (.A2(_07194_),
    .A1(_07193_),
    .B1(_02480_),
    .X(_07195_));
 sg13g2_o21ai_1 _15855_ (.B1(_06235_),
    .Y(_07196_),
    .A1(_02793_),
    .A2(_07186_));
 sg13g2_o21ai_1 _15856_ (.B1(_07195_),
    .Y(_07197_),
    .A1(net1851),
    .A2(_07196_));
 sg13g2_nand2_1 _15857_ (.Y(_07198_),
    .A(net2359),
    .B(net1806));
 sg13g2_o21ai_1 _15858_ (.B1(_07198_),
    .Y(_00906_),
    .A1(net1806),
    .A2(_07197_));
 sg13g2_o21ai_1 _15859_ (.B1(net2135),
    .Y(_07199_),
    .A1(_02530_),
    .A2(_06081_));
 sg13g2_a21oi_1 _15860_ (.A1(_07185_),
    .A2(_07199_),
    .Y(_07200_),
    .B1(net2070));
 sg13g2_nor2_1 _15861_ (.A(net1851),
    .B(_07200_),
    .Y(_07201_));
 sg13g2_xor2_1 _15862_ (.B(_07193_),
    .A(net4042),
    .X(_07202_));
 sg13g2_a221oi_1 _15863_ (.B2(net1851),
    .C1(net1805),
    .B1(_07202_),
    .A1(_06238_),
    .Y(_07203_),
    .A2(_07201_));
 sg13g2_a21o_1 _15864_ (.A2(net1805),
    .A1(net4042),
    .B1(_07203_),
    .X(_00907_));
 sg13g2_a221oi_1 _15865_ (.B2(_02536_),
    .C1(net2069),
    .B1(_06081_),
    .A1(_02551_),
    .Y(_07204_),
    .A2(_02774_));
 sg13g2_a21oi_1 _15866_ (.A1(net2069),
    .A2(_07158_),
    .Y(_07205_),
    .B1(_07204_));
 sg13g2_o21ai_1 _15867_ (.B1(net2498),
    .Y(_07206_),
    .A1(net4012),
    .A2(net1851));
 sg13g2_a21oi_1 _15868_ (.A1(net4012),
    .A2(_02750_),
    .Y(_07207_),
    .B1(_07206_));
 sg13g2_a21o_1 _15869_ (.A2(_07205_),
    .A1(net1793),
    .B1(_07207_),
    .X(_00908_));
 sg13g2_and2_1 _15870_ (.A(net3839),
    .B(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .X(_07208_));
 sg13g2_o21ai_1 _15871_ (.B1(_01433_),
    .Y(_07209_),
    .A1(net3839),
    .A2(\i_tinyqv.cpu.additional_mem_ops[0] ));
 sg13g2_nand3_1 _15872_ (.B(net2139),
    .C(_07150_),
    .A(net2069),
    .Y(_07210_));
 sg13g2_a22oi_1 _15873_ (.Y(_07211_),
    .B1(_02788_),
    .B2(_06081_),
    .A2(_02774_),
    .A1(_02550_));
 sg13g2_nand2_1 _15874_ (.Y(_07212_),
    .A(net2069),
    .B(_07157_));
 sg13g2_nand4_1 _15875_ (.B(_07210_),
    .C(_07211_),
    .A(_02480_),
    .Y(_07213_),
    .D(_07212_));
 sg13g2_o21ai_1 _15876_ (.B1(_07213_),
    .Y(_07214_),
    .A1(_07208_),
    .A2(_07209_));
 sg13g2_o21ai_1 _15877_ (.B1(net2498),
    .Y(_07215_),
    .A1(net3839),
    .A2(_02750_));
 sg13g2_a21oi_1 _15878_ (.A1(_02750_),
    .A2(_07214_),
    .Y(_00909_),
    .B1(_07215_));
 sg13g2_a22oi_1 _15879_ (.Y(_07216_),
    .B1(_06081_),
    .B2(_02534_),
    .A2(_02774_),
    .A1(_02548_));
 sg13g2_nand2_1 _15880_ (.Y(_07217_),
    .A(_02750_),
    .B(_07209_));
 sg13g2_nand3_1 _15881_ (.B(net2498),
    .C(_07217_),
    .A(net2857),
    .Y(_07218_));
 sg13g2_o21ai_1 _15882_ (.B1(net2858),
    .Y(_00910_),
    .A1(net1783),
    .A2(_07216_));
 sg13g2_a21o_1 _15883_ (.A2(net1852),
    .A1(net3916),
    .B1(net1818),
    .X(_07219_));
 sg13g2_o21ai_1 _15884_ (.B1(net2488),
    .Y(_07220_),
    .A1(net3916),
    .A2(net1852));
 sg13g2_nor2_1 _15885_ (.A(_07219_),
    .B(_07220_),
    .Y(_00911_));
 sg13g2_a21oi_1 _15886_ (.A1(\i_tinyqv.cpu.addr_offset[2] ),
    .A2(net1852),
    .Y(_07221_),
    .B1(net2801));
 sg13g2_nand2b_1 _15887_ (.Y(_07222_),
    .B(net2490),
    .A_N(_07221_));
 sg13g2_a21oi_1 _15888_ (.A1(net2801),
    .A2(_07219_),
    .Y(_00912_),
    .B1(_07222_));
 sg13g2_mux2_1 _15889_ (.A0(net3699),
    .A1(_07212_),
    .S(net1793),
    .X(_00913_));
 sg13g2_a21oi_1 _15890_ (.A1(net3476),
    .A2(_06042_),
    .Y(_07223_),
    .B1(_02747_));
 sg13g2_nor2_1 _15891_ (.A(net2340),
    .B(_07223_),
    .Y(_00914_));
 sg13g2_nor3_1 _15892_ (.A(_02512_),
    .B(_02555_),
    .C(_02747_),
    .Y(_07224_));
 sg13g2_nor2_1 _15893_ (.A(_06042_),
    .B(_07224_),
    .Y(_07225_));
 sg13g2_and2_1 _15894_ (.A(_00923_),
    .B(_06042_),
    .X(_07226_));
 sg13g2_nor3_1 _15895_ (.A(net2339),
    .B(_07225_),
    .C(_07226_),
    .Y(_00915_));
 sg13g2_nand2b_2 _15896_ (.Y(_07227_),
    .B(net2271),
    .A_N(_02834_));
 sg13g2_nor2_1 _15897_ (.A(net2737),
    .B(net2254),
    .Y(_00916_));
 sg13g2_or2_1 _15898_ (.X(_07228_),
    .B(net4081),
    .A(net2737));
 sg13g2_and3_1 _15899_ (.X(_00917_),
    .A(net2271),
    .B(_02827_),
    .C(_07228_));
 sg13g2_nand3_1 _15900_ (.B(net4169),
    .C(net3983),
    .A(net2737),
    .Y(_07229_));
 sg13g2_xnor2_1 _15901_ (.Y(_07230_),
    .A(_01107_),
    .B(_02827_));
 sg13g2_nor2_1 _15902_ (.A(_07227_),
    .B(net3984),
    .Y(_00918_));
 sg13g2_nor2_1 _15903_ (.A(_01108_),
    .B(_07229_),
    .Y(_07231_));
 sg13g2_and2_1 _15904_ (.A(_01108_),
    .B(_07229_),
    .X(_07232_));
 sg13g2_nor3_1 _15905_ (.A(_07227_),
    .B(_07231_),
    .C(net4021),
    .Y(_00919_));
 sg13g2_and2_1 _15906_ (.A(net3431),
    .B(_07231_),
    .X(_07233_));
 sg13g2_nor2_1 _15907_ (.A(net3431),
    .B(_07231_),
    .Y(_07234_));
 sg13g2_nor3_1 _15908_ (.A(_07227_),
    .B(_07233_),
    .C(net3432),
    .Y(_00920_));
 sg13g2_nand2_1 _15909_ (.Y(_07235_),
    .A(net3506),
    .B(_07233_));
 sg13g2_xnor2_1 _15910_ (.Y(_07236_),
    .A(net3506),
    .B(_07233_));
 sg13g2_nor2_1 _15911_ (.A(_07227_),
    .B(net3507),
    .Y(_00921_));
 sg13g2_xor2_1 _15912_ (.B(_07235_),
    .A(net3701),
    .X(_07237_));
 sg13g2_nor2_1 _15913_ (.A(_07227_),
    .B(_07237_),
    .Y(_00922_));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_dfrbpq_2 _15915_ (.RESET_B(net1422),
    .D(_00077_),
    .Q(\i_tinyqv.cpu.instr_write_offset[3] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_1 _15916_ (.RESET_B(net1256),
    .D(net3405),
    .Q(\i_tinyqv.cpu.instr_data[1][2] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _15917_ (.RESET_B(net1255),
    .D(net3457),
    .Q(\i_tinyqv.cpu.instr_data[1][3] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _15918_ (.RESET_B(net1254),
    .D(_00080_),
    .Q(\i_tinyqv.cpu.instr_data[1][4] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _15919_ (.RESET_B(net1253),
    .D(net3347),
    .Q(\i_tinyqv.cpu.instr_data[1][5] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _15920_ (.RESET_B(net1252),
    .D(net3411),
    .Q(\i_tinyqv.cpu.instr_data[1][6] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _15921_ (.RESET_B(net1251),
    .D(net3128),
    .Q(\i_tinyqv.cpu.instr_data[1][7] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _15922_ (.RESET_B(net1250),
    .D(net3528),
    .Q(\i_tinyqv.cpu.instr_data[1][8] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _15923_ (.RESET_B(net1249),
    .D(net3121),
    .Q(\i_tinyqv.cpu.instr_data[1][9] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _15924_ (.RESET_B(net1248),
    .D(net3374),
    .Q(\i_tinyqv.cpu.instr_data[1][10] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _15925_ (.RESET_B(net1247),
    .D(net3143),
    .Q(\i_tinyqv.cpu.instr_data[1][11] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _15926_ (.RESET_B(net1246),
    .D(net3624),
    .Q(\i_tinyqv.cpu.instr_data[1][12] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _15927_ (.RESET_B(net1245),
    .D(net3090),
    .Q(\i_tinyqv.cpu.instr_data[1][13] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _15928_ (.RESET_B(net1244),
    .D(net3058),
    .Q(\i_tinyqv.cpu.instr_data[1][14] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _15929_ (.RESET_B(net1423),
    .D(net3384),
    .Q(\i_tinyqv.cpu.instr_data[1][15] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _15930_ (.RESET_B(net1424),
    .D(net1486),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_2 _15931_ (.RESET_B(net1425),
    .D(net2514),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_2 _15932_ (.RESET_B(net1426),
    .D(net2651),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_2 _15933_ (.RESET_B(net1427),
    .D(net1520),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _15934_ (.RESET_B(net1428),
    .D(net1608),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _15935_ (.RESET_B(net1429),
    .D(net1575),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _15936_ (.RESET_B(net1430),
    .D(net1478),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _15937_ (.RESET_B(net1431),
    .D(net2591),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _15938_ (.RESET_B(net1432),
    .D(net2531),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15939_ (.RESET_B(net1433),
    .D(net2561),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _15940_ (.RESET_B(net14),
    .D(net2544),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _15941_ (.RESET_B(net15),
    .D(net2527),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _15942_ (.RESET_B(net16),
    .D(net1544),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15943_ (.RESET_B(net17),
    .D(net1570),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15944_ (.RESET_B(net18),
    .D(net2584),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _15945_ (.RESET_B(net19),
    .D(net1676),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _15946_ (.RESET_B(net20),
    .D(net2564),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15947_ (.RESET_B(net21),
    .D(net2632),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15948_ (.RESET_B(net22),
    .D(net1535),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _15949_ (.RESET_B(net23),
    .D(net2533),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _15950_ (.RESET_B(net24),
    .D(net2537),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15951_ (.RESET_B(net25),
    .D(net2511),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _15952_ (.RESET_B(net26),
    .D(net2660),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _15953_ (.RESET_B(net27),
    .D(net1645),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _15954_ (.RESET_B(net28),
    .D(net1637),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _15955_ (.RESET_B(net29),
    .D(net1634),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15956_ (.RESET_B(net35),
    .D(net2530),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _15957_ (.RESET_B(net1243),
    .D(net2665),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _15958_ (.RESET_B(net1242),
    .D(net4069),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _15959_ (.RESET_B(net1241),
    .D(net4047),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _15960_ (.RESET_B(net1240),
    .D(net3731),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _15961_ (.RESET_B(net1239),
    .D(_00095_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _15962_ (.RESET_B(net36),
    .D(net3255),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.cy ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _15963_ (.RESET_B(net37),
    .D(net2695),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[0] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _15964_ (.RESET_B(net38),
    .D(net2698),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _15965_ (.RESET_B(net39),
    .D(net2735),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_2 _15966_ (.RESET_B(net40),
    .D(net2666),
    .Q(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _15967_ (.RESET_B(net41),
    .D(net1522),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _15968_ (.RESET_B(net42),
    .D(net2676),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_2 _15969_ (.RESET_B(net43),
    .D(net1514),
    .Q(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15970_ (.RESET_B(net44),
    .D(net2552),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _15971_ (.RESET_B(net45),
    .D(net1668),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _15972_ (.RESET_B(net46),
    .D(net2610),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _15973_ (.RESET_B(net47),
    .D(net2541),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15974_ (.RESET_B(net48),
    .D(net1578),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15975_ (.RESET_B(net49),
    .D(net2686),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _15976_ (.RESET_B(net50),
    .D(net2573),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _15977_ (.RESET_B(net51),
    .D(net1627),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15978_ (.RESET_B(net52),
    .D(net1611),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15979_ (.RESET_B(net53),
    .D(net2589),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _15980_ (.RESET_B(net54),
    .D(net1642),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _15981_ (.RESET_B(net55),
    .D(net1468),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15982_ (.RESET_B(net56),
    .D(net1606),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15983_ (.RESET_B(net57),
    .D(net1619),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _15984_ (.RESET_B(net58),
    .D(net1530),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _15985_ (.RESET_B(net59),
    .D(net1560),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _15986_ (.RESET_B(net60),
    .D(net1469),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .CLK(clknet_leaf_166_clk_regs));
 sg13g2_dfrbpq_1 _15987_ (.RESET_B(net61),
    .D(net2641),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _15988_ (.RESET_B(net62),
    .D(net1590),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _15989_ (.RESET_B(net69),
    .D(net1554),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _15990_ (.RESET_B(net1238),
    .D(net1664),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _15991_ (.RESET_B(net1237),
    .D(_00097_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _15992_ (.RESET_B(net1236),
    .D(_00098_),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _15993_ (.RESET_B(net1235),
    .D(net3890),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .CLK(clknet_leaf_162_clk_regs));
 sg13g2_dfrbpq_1 _15994_ (.RESET_B(net1234),
    .D(_00100_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _15995_ (.RESET_B(net1233),
    .D(net3901),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .CLK(clknet_leaf_167_clk_regs));
 sg13g2_dfrbpq_1 _15996_ (.RESET_B(net70),
    .D(_00102_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _15997_ (.RESET_B(net71),
    .D(net2731),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_2 _15998_ (.RESET_B(net72),
    .D(net2718),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_1 _15999_ (.RESET_B(net73),
    .D(net2732),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16000_ (.RESET_B(net74),
    .D(net2733),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16001_ (.RESET_B(net75),
    .D(net2547),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_2 _16002_ (.RESET_B(net76),
    .D(net2543),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_2 _16003_ (.RESET_B(net77),
    .D(net1661),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_2 _16004_ (.RESET_B(net78),
    .D(net1604),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16005_ (.RESET_B(net79),
    .D(net1456),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16006_ (.RESET_B(net80),
    .D(net1665),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16007_ (.RESET_B(net81),
    .D(net2667),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16008_ (.RESET_B(net82),
    .D(net2586),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16009_ (.RESET_B(net83),
    .D(net1548),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _16010_ (.RESET_B(net84),
    .D(net1643),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16011_ (.RESET_B(net85),
    .D(net2515),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16012_ (.RESET_B(net86),
    .D(net1505),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16013_ (.RESET_B(net87),
    .D(net2582),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _16014_ (.RESET_B(net88),
    .D(net2648),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _16015_ (.RESET_B(net89),
    .D(net1495),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16016_ (.RESET_B(net90),
    .D(net1497),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16017_ (.RESET_B(net91),
    .D(net1675),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16018_ (.RESET_B(net92),
    .D(net1603),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _16019_ (.RESET_B(net93),
    .D(net1545),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16020_ (.RESET_B(net94),
    .D(net1481),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16021_ (.RESET_B(net95),
    .D(net2600),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16022_ (.RESET_B(net96),
    .D(net2596),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _16023_ (.RESET_B(net97),
    .D(net2538),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16024_ (.RESET_B(net98),
    .D(net1656),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16025_ (.RESET_B(net99),
    .D(_00041_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16026_ (.RESET_B(net100),
    .D(_00042_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16027_ (.RESET_B(net101),
    .D(_00043_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16028_ (.RESET_B(net102),
    .D(_00044_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_2 _16029_ (.RESET_B(net103),
    .D(net2700),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16030_ (.RESET_B(net104),
    .D(net2717),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_2 _16031_ (.RESET_B(net105),
    .D(net2716),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_2 _16032_ (.RESET_B(net106),
    .D(net2704),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _16033_ (.RESET_B(net107),
    .D(net1475),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16034_ (.RESET_B(net108),
    .D(net1436),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16035_ (.RESET_B(net109),
    .D(net1595),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16036_ (.RESET_B(net110),
    .D(net1538),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16037_ (.RESET_B(net111),
    .D(net2635),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_1 _16038_ (.RESET_B(net112),
    .D(net2678),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16039_ (.RESET_B(net113),
    .D(net1591),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16040_ (.RESET_B(net114),
    .D(net1667),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16041_ (.RESET_B(net115),
    .D(net1636),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16042_ (.RESET_B(net116),
    .D(net1439),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16043_ (.RESET_B(net117),
    .D(net1465),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16044_ (.RESET_B(net118),
    .D(net2611),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16045_ (.RESET_B(net119),
    .D(net1489),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16046_ (.RESET_B(net120),
    .D(net2677),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16047_ (.RESET_B(net121),
    .D(net1440),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _16048_ (.RESET_B(net122),
    .D(net1556),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16049_ (.RESET_B(net123),
    .D(net2597),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16050_ (.RESET_B(net124),
    .D(net1466),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16051_ (.RESET_B(net125),
    .D(net2672),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16052_ (.RESET_B(net126),
    .D(net2513),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16053_ (.RESET_B(net127),
    .D(net1510),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16054_ (.RESET_B(net128),
    .D(net1580),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _16055_ (.RESET_B(net129),
    .D(net2560),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _16056_ (.RESET_B(net130),
    .D(net1574),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16057_ (.RESET_B(net131),
    .D(_00037_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16058_ (.RESET_B(net132),
    .D(_00038_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _16059_ (.RESET_B(net133),
    .D(_00039_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _16060_ (.RESET_B(net134),
    .D(_00040_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_2 _16061_ (.RESET_B(net135),
    .D(net1612),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16062_ (.RESET_B(net136),
    .D(net2687),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_2 _16063_ (.RESET_B(net137),
    .D(net1558),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_2 _16064_ (.RESET_B(net138),
    .D(net2680),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16065_ (.RESET_B(net139),
    .D(net2570),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16066_ (.RESET_B(net140),
    .D(net2617),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16067_ (.RESET_B(net141),
    .D(net1641),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _16068_ (.RESET_B(net142),
    .D(net2642),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16069_ (.RESET_B(net143),
    .D(net1516),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16070_ (.RESET_B(net144),
    .D(net2545),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16071_ (.RESET_B(net145),
    .D(net2606),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16072_ (.RESET_B(net146),
    .D(net2621),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16073_ (.RESET_B(net147),
    .D(net1536),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16074_ (.RESET_B(net148),
    .D(net1512),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16075_ (.RESET_B(net149),
    .D(net1500),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16076_ (.RESET_B(net150),
    .D(net1458),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16077_ (.RESET_B(net151),
    .D(net2566),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16078_ (.RESET_B(net152),
    .D(net1451),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16079_ (.RESET_B(net153),
    .D(net2540),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16080_ (.RESET_B(net154),
    .D(net1657),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16081_ (.RESET_B(net155),
    .D(net2571),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16082_ (.RESET_B(net156),
    .D(net2623),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _16083_ (.RESET_B(net157),
    .D(net2601),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16084_ (.RESET_B(net158),
    .D(net1506),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16085_ (.RESET_B(net159),
    .D(net2572),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16086_ (.RESET_B(net160),
    .D(net1477),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _16087_ (.RESET_B(net161),
    .D(net1537),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16088_ (.RESET_B(net162),
    .D(net1607),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16089_ (.RESET_B(net163),
    .D(_00033_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16090_ (.RESET_B(net164),
    .D(_00034_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_165_clk_regs));
 sg13g2_dfrbpq_1 _16091_ (.RESET_B(net165),
    .D(_00035_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16092_ (.RESET_B(net166),
    .D(_00036_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16093_ (.RESET_B(net167),
    .D(net2719),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_2 _16094_ (.RESET_B(net168),
    .D(net2714),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16095_ (.RESET_B(net169),
    .D(net2702),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_2 _16096_ (.RESET_B(net170),
    .D(net2712),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16097_ (.RESET_B(net171),
    .D(net2594),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16098_ (.RESET_B(net172),
    .D(net2637),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16099_ (.RESET_B(net173),
    .D(net2549),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16100_ (.RESET_B(net174),
    .D(net1639),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16101_ (.RESET_B(net175),
    .D(net2528),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16102_ (.RESET_B(net176),
    .D(net2542),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16103_ (.RESET_B(net177),
    .D(net2517),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16104_ (.RESET_B(net178),
    .D(net2624),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16105_ (.RESET_B(net179),
    .D(net1467),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16106_ (.RESET_B(net180),
    .D(net1633),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16107_ (.RESET_B(net181),
    .D(net2526),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16108_ (.RESET_B(net182),
    .D(net1566),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16109_ (.RESET_B(net183),
    .D(net1519),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16110_ (.RESET_B(net184),
    .D(net1483),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16111_ (.RESET_B(net185),
    .D(net1623),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_127_clk_regs));
 sg13g2_dfrbpq_1 _16112_ (.RESET_B(net186),
    .D(net2551),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16113_ (.RESET_B(net187),
    .D(net1582),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16114_ (.RESET_B(net188),
    .D(net1593),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16115_ (.RESET_B(net189),
    .D(net1553),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16116_ (.RESET_B(net190),
    .D(net1551),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16117_ (.RESET_B(net191),
    .D(net1602),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16118_ (.RESET_B(net192),
    .D(net1504),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16119_ (.RESET_B(net193),
    .D(net2585),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16120_ (.RESET_B(net194),
    .D(net2520),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16121_ (.RESET_B(net195),
    .D(_00029_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16122_ (.RESET_B(net196),
    .D(_00030_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16123_ (.RESET_B(net197),
    .D(_00031_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16124_ (.RESET_B(net198),
    .D(_00032_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_2 _16125_ (.RESET_B(net199),
    .D(net2724),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16126_ (.RESET_B(net200),
    .D(net2647),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_2 _16127_ (.RESET_B(net201),
    .D(net2644),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_2 _16128_ (.RESET_B(net202),
    .D(net2736),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .CLK(clknet_leaf_126_clk_regs));
 sg13g2_dfrbpq_1 _16129_ (.RESET_B(net203),
    .D(net1658),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16130_ (.RESET_B(net204),
    .D(net2519),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16131_ (.RESET_B(net205),
    .D(net1592),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_2 _16132_ (.RESET_B(net206),
    .D(net1473),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16133_ (.RESET_B(net207),
    .D(net2592),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16134_ (.RESET_B(net208),
    .D(net1654),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16135_ (.RESET_B(net209),
    .D(net1681),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _16136_ (.RESET_B(net210),
    .D(net2603),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16137_ (.RESET_B(net211),
    .D(net2605),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16138_ (.RESET_B(net212),
    .D(net1618),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16139_ (.RESET_B(net213),
    .D(net1470),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16140_ (.RESET_B(net214),
    .D(net1472),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16141_ (.RESET_B(net215),
    .D(net2508),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16142_ (.RESET_B(net216),
    .D(net2593),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16143_ (.RESET_B(net217),
    .D(net1626),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16144_ (.RESET_B(net218),
    .D(net1515),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16145_ (.RESET_B(net219),
    .D(net1565),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16146_ (.RESET_B(net220),
    .D(net1487),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16147_ (.RESET_B(net221),
    .D(net1494),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16148_ (.RESET_B(net222),
    .D(net1543),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16149_ (.RESET_B(net223),
    .D(net1674),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_1 _16150_ (.RESET_B(net224),
    .D(net1650),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16151_ (.RESET_B(net225),
    .D(net1525),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16152_ (.RESET_B(net226),
    .D(net1550),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16153_ (.RESET_B(net227),
    .D(_00025_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16154_ (.RESET_B(net228),
    .D(_00026_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16155_ (.RESET_B(net229),
    .D(_00027_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16156_ (.RESET_B(net230),
    .D(_00028_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_2 _16157_ (.RESET_B(net231),
    .D(net2691),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16158_ (.RESET_B(net232),
    .D(net2725),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_2 _16159_ (.RESET_B(net233),
    .D(net2705),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_2 _16160_ (.RESET_B(net234),
    .D(net2723),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _16161_ (.RESET_B(net235),
    .D(net1583),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_2 _16162_ (.RESET_B(net236),
    .D(net1646),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16163_ (.RESET_B(net237),
    .D(net2640),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16164_ (.RESET_B(net238),
    .D(net2536),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16165_ (.RESET_B(net239),
    .D(net2557),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _16166_ (.RESET_B(net240),
    .D(net1480),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16167_ (.RESET_B(net241),
    .D(net2563),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16168_ (.RESET_B(net242),
    .D(net2631),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16169_ (.RESET_B(net243),
    .D(net2558),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _16170_ (.RESET_B(net244),
    .D(net2620),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16171_ (.RESET_B(net245),
    .D(net1445),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16172_ (.RESET_B(net246),
    .D(net1531),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16173_ (.RESET_B(net247),
    .D(net2580),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _16174_ (.RESET_B(net248),
    .D(net2655),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16175_ (.RESET_B(net249),
    .D(net1640),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16176_ (.RESET_B(net250),
    .D(net1529),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16177_ (.RESET_B(net251),
    .D(net1586),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _16178_ (.RESET_B(net252),
    .D(net2569),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16179_ (.RESET_B(net253),
    .D(net2523),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16180_ (.RESET_B(net254),
    .D(net1485),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16181_ (.RESET_B(net255),
    .D(net2658),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _16182_ (.RESET_B(net256),
    .D(net1555),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16183_ (.RESET_B(net257),
    .D(net1569),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16184_ (.RESET_B(net258),
    .D(net1613),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16185_ (.RESET_B(net259),
    .D(_00021_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16186_ (.RESET_B(net260),
    .D(_00022_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16187_ (.RESET_B(net261),
    .D(_00023_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16188_ (.RESET_B(net262),
    .D(_00024_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16189_ (.RESET_B(net263),
    .D(net2709),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16190_ (.RESET_B(net264),
    .D(net2730),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .CLK(clknet_leaf_128_clk_regs));
 sg13g2_dfrbpq_2 _16191_ (.RESET_B(net265),
    .D(net2693),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_2 _16192_ (.RESET_B(net266),
    .D(net2697),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16193_ (.RESET_B(net267),
    .D(net2525),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16194_ (.RESET_B(net268),
    .D(net2516),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16195_ (.RESET_B(net269),
    .D(net1629),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16196_ (.RESET_B(net270),
    .D(net2634),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16197_ (.RESET_B(net271),
    .D(net1464),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_125_clk_regs));
 sg13g2_dfrbpq_1 _16198_ (.RESET_B(net272),
    .D(net1679),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16199_ (.RESET_B(net273),
    .D(net1453),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16200_ (.RESET_B(net274),
    .D(net1461),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16201_ (.RESET_B(net275),
    .D(net2618),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16202_ (.RESET_B(net276),
    .D(net1476),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16203_ (.RESET_B(net277),
    .D(net2507),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16204_ (.RESET_B(net278),
    .D(net2616),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16205_ (.RESET_B(net279),
    .D(net1511),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16206_ (.RESET_B(net280),
    .D(net1549),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16207_ (.RESET_B(net281),
    .D(net1521),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16208_ (.RESET_B(net282),
    .D(net1462),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_120_clk_regs));
 sg13g2_dfrbpq_1 _16209_ (.RESET_B(net283),
    .D(net2652),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16210_ (.RESET_B(net284),
    .D(net1474),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_119_clk_regs));
 sg13g2_dfrbpq_1 _16211_ (.RESET_B(net285),
    .D(net1625),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16212_ (.RESET_B(net286),
    .D(net1609),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16213_ (.RESET_B(net287),
    .D(net1517),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16214_ (.RESET_B(net288),
    .D(net2567),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_121_clk_regs));
 sg13g2_dfrbpq_1 _16215_ (.RESET_B(net289),
    .D(net2534),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16216_ (.RESET_B(net290),
    .D(net1638),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_123_clk_regs));
 sg13g2_dfrbpq_1 _16217_ (.RESET_B(net291),
    .D(_00069_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16218_ (.RESET_B(net292),
    .D(_00070_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_122_clk_regs));
 sg13g2_dfrbpq_1 _16219_ (.RESET_B(net293),
    .D(_00071_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _16220_ (.RESET_B(net294),
    .D(_00072_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_124_clk_regs));
 sg13g2_dfrbpq_2 _16221_ (.RESET_B(net295),
    .D(net2722),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16222_ (.RESET_B(net296),
    .D(net2703),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_2 _16223_ (.RESET_B(net297),
    .D(net2728),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_2 _16224_ (.RESET_B(net298),
    .D(net2721),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_2 _16225_ (.RESET_B(net299),
    .D(net1455),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16226_ (.RESET_B(net300),
    .D(net1492),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_2 _16227_ (.RESET_B(net301),
    .D(net1663),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16228_ (.RESET_B(net302),
    .D(net1678),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16229_ (.RESET_B(net303),
    .D(net2645),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16230_ (.RESET_B(net304),
    .D(net1540),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16231_ (.RESET_B(net305),
    .D(net2649),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16232_ (.RESET_B(net306),
    .D(net2607),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16233_ (.RESET_B(net307),
    .D(net2622),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16234_ (.RESET_B(net308),
    .D(net2550),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16235_ (.RESET_B(net309),
    .D(net1649),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16236_ (.RESET_B(net310),
    .D(net2614),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16237_ (.RESET_B(net311),
    .D(net1579),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16238_ (.RESET_B(net312),
    .D(net2535),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16239_ (.RESET_B(net313),
    .D(net2518),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_116_clk_regs));
 sg13g2_dfrbpq_1 _16240_ (.RESET_B(net314),
    .D(net1454),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16241_ (.RESET_B(net315),
    .D(net1471),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_115_clk_regs));
 sg13g2_dfrbpq_1 _16242_ (.RESET_B(net316),
    .D(net1513),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16243_ (.RESET_B(net317),
    .D(net1463),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_117_clk_regs));
 sg13g2_dfrbpq_1 _16244_ (.RESET_B(net318),
    .D(net2529),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16245_ (.RESET_B(net319),
    .D(net1572),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _16246_ (.RESET_B(net320),
    .D(net1588),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16247_ (.RESET_B(net321),
    .D(net2548),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16248_ (.RESET_B(net322),
    .D(net2659),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16249_ (.RESET_B(net323),
    .D(_00065_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _16250_ (.RESET_B(net324),
    .D(_00066_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_113_clk_regs));
 sg13g2_dfrbpq_1 _16251_ (.RESET_B(net325),
    .D(_00067_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_114_clk_regs));
 sg13g2_dfrbpq_1 _16252_ (.RESET_B(net326),
    .D(_00068_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_118_clk_regs));
 sg13g2_dfrbpq_1 _16253_ (.RESET_B(net327),
    .D(net2715),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _16254_ (.RESET_B(net328),
    .D(net2726),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_2 _16255_ (.RESET_B(net329),
    .D(net2713),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _16256_ (.RESET_B(net330),
    .D(net2727),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16257_ (.RESET_B(net331),
    .D(net1610),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16258_ (.RESET_B(net332),
    .D(net1666),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16259_ (.RESET_B(net333),
    .D(net2674),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16260_ (.RESET_B(net334),
    .D(net2626),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16261_ (.RESET_B(net335),
    .D(net1541),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16262_ (.RESET_B(net336),
    .D(net1482),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16263_ (.RESET_B(net337),
    .D(net1587),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16264_ (.RESET_B(net338),
    .D(net1490),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_106_clk_regs));
 sg13g2_dfrbpq_1 _16265_ (.RESET_B(net339),
    .D(net2568),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16266_ (.RESET_B(net340),
    .D(net1653),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16267_ (.RESET_B(net341),
    .D(net1438),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_105_clk_regs));
 sg13g2_dfrbpq_1 _16268_ (.RESET_B(net342),
    .D(net2559),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16269_ (.RESET_B(net343),
    .D(net2562),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16270_ (.RESET_B(net344),
    .D(net1669),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16271_ (.RESET_B(net345),
    .D(net2604),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16272_ (.RESET_B(net346),
    .D(net1496),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16273_ (.RESET_B(net347),
    .D(net2675),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16274_ (.RESET_B(net348),
    .D(net1584),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16275_ (.RESET_B(net349),
    .D(net1503),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16276_ (.RESET_B(net350),
    .D(net1630),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16277_ (.RESET_B(net351),
    .D(net1443),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _16278_ (.RESET_B(net352),
    .D(net2555),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16279_ (.RESET_B(net353),
    .D(net1576),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16280_ (.RESET_B(net354),
    .D(net2669),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_107_clk_regs));
 sg13g2_dfrbpq_1 _16281_ (.RESET_B(net355),
    .D(_00061_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_103_clk_regs));
 sg13g2_dfrbpq_1 _16282_ (.RESET_B(net356),
    .D(_00062_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_1 _16283_ (.RESET_B(net357),
    .D(_00063_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_1 _16284_ (.RESET_B(net358),
    .D(_00064_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_108_clk_regs));
 sg13g2_dfrbpq_2 _16285_ (.RESET_B(net359),
    .D(net1628),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _16286_ (.RESET_B(net360),
    .D(net2708),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _16287_ (.RESET_B(net361),
    .D(net2688),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_2 _16288_ (.RESET_B(net362),
    .D(net2720),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _16289_ (.RESET_B(net363),
    .D(net2692),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _16290_ (.RESET_B(net364),
    .D(net1632),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _16291_ (.RESET_B(net365),
    .D(net2671),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_104_clk_regs));
 sg13g2_dfrbpq_2 _16292_ (.RESET_B(net366),
    .D(net1532),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16293_ (.RESET_B(net367),
    .D(net1444),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _16294_ (.RESET_B(net368),
    .D(net2630),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _16295_ (.RESET_B(net369),
    .D(net1457),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _16296_ (.RESET_B(net370),
    .D(net2650),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_109_clk_regs));
 sg13g2_dfrbpq_1 _16297_ (.RESET_B(net371),
    .D(net2581),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16298_ (.RESET_B(net372),
    .D(net2532),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _16299_ (.RESET_B(net373),
    .D(net2639),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _16300_ (.RESET_B(net374),
    .D(net1652),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16301_ (.RESET_B(net375),
    .D(net2512),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16302_ (.RESET_B(net376),
    .D(net1615),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_102_clk_regs));
 sg13g2_dfrbpq_1 _16303_ (.RESET_B(net377),
    .D(net1585),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _16304_ (.RESET_B(net378),
    .D(net1651),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16305_ (.RESET_B(net379),
    .D(net2629),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16306_ (.RESET_B(net380),
    .D(net1573),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _16307_ (.RESET_B(net381),
    .D(net2574),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _16308_ (.RESET_B(net382),
    .D(net1561),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16309_ (.RESET_B(net383),
    .D(net2664),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16310_ (.RESET_B(net384),
    .D(net1459),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _16311_ (.RESET_B(net385),
    .D(net2546),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _16312_ (.RESET_B(net386),
    .D(net2575),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_110_clk_regs));
 sg13g2_dfrbpq_1 _16313_ (.RESET_B(net387),
    .D(_00057_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _16314_ (.RESET_B(net388),
    .D(_00058_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _16315_ (.RESET_B(net389),
    .D(_00059_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_101_clk_regs));
 sg13g2_dfrbpq_1 _16316_ (.RESET_B(net390),
    .D(_00060_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _16317_ (.RESET_B(net391),
    .D(net1648),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_1 _16318_ (.RESET_B(net392),
    .D(net2682),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .CLK(clknet_leaf_131_clk_regs));
 sg13g2_dfrbpq_2 _16319_ (.RESET_B(net393),
    .D(net2627),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_2 _16320_ (.RESET_B(net394),
    .D(net2662),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_1 _16321_ (.RESET_B(net395),
    .D(net1616),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _16322_ (.RESET_B(net396),
    .D(net2628),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_112_clk_regs));
 sg13g2_dfrbpq_1 _16323_ (.RESET_B(net397),
    .D(net1647),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_1 _16324_ (.RESET_B(net398),
    .D(net2663),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_133_clk_regs));
 sg13g2_dfrbpq_1 _16325_ (.RESET_B(net399),
    .D(net1508),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16326_ (.RESET_B(net400),
    .D(net2643),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_111_clk_regs));
 sg13g2_dfrbpq_1 _16327_ (.RESET_B(net401),
    .D(net1594),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16328_ (.RESET_B(net402),
    .D(net2612),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16329_ (.RESET_B(net403),
    .D(net1624),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16330_ (.RESET_B(net404),
    .D(net1680),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16331_ (.RESET_B(net405),
    .D(net1534),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16332_ (.RESET_B(net406),
    .D(net1509),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16333_ (.RESET_B(net407),
    .D(net1601),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16334_ (.RESET_B(net408),
    .D(net1655),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16335_ (.RESET_B(net409),
    .D(net1527),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16336_ (.RESET_B(net410),
    .D(net1597),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_134_clk_regs));
 sg13g2_dfrbpq_1 _16337_ (.RESET_B(net411),
    .D(net1622),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16338_ (.RESET_B(net412),
    .D(net2595),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_130_clk_regs));
 sg13g2_dfrbpq_1 _16339_ (.RESET_B(net413),
    .D(net1484),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16340_ (.RESET_B(net414),
    .D(net1581),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16341_ (.RESET_B(net415),
    .D(net1677),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16342_ (.RESET_B(net416),
    .D(net1567),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16343_ (.RESET_B(net417),
    .D(net2522),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _16344_ (.RESET_B(net418),
    .D(net2653),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16345_ (.RESET_B(net419),
    .D(_00053_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16346_ (.RESET_B(net420),
    .D(_00054_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_129_clk_regs));
 sg13g2_dfrbpq_1 _16347_ (.RESET_B(net421),
    .D(_00055_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _16348_ (.RESET_B(net422),
    .D(_00056_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_2 _16349_ (.RESET_B(net423),
    .D(net2670),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .CLK(clknet_leaf_132_clk_regs));
 sg13g2_dfrbpq_2 _16350_ (.RESET_B(net424),
    .D(net2689),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_2 _16351_ (.RESET_B(net425),
    .D(net1605),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .CLK(clknet_leaf_137_clk_regs));
 sg13g2_dfrbpq_2 _16352_ (.RESET_B(net426),
    .D(net1488),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _16353_ (.RESET_B(net427),
    .D(net1546),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16354_ (.RESET_B(net428),
    .D(net1559),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16355_ (.RESET_B(net429),
    .D(net1614),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16356_ (.RESET_B(net430),
    .D(net1499),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16357_ (.RESET_B(net431),
    .D(net1528),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16358_ (.RESET_B(net432),
    .D(net2646),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_139_clk_regs));
 sg13g2_dfrbpq_1 _16359_ (.RESET_B(net433),
    .D(net1598),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_142_clk_regs));
 sg13g2_dfrbpq_1 _16360_ (.RESET_B(net434),
    .D(net1523),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16361_ (.RESET_B(net435),
    .D(net2608),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_135_clk_regs));
 sg13g2_dfrbpq_1 _16362_ (.RESET_B(net436),
    .D(net1617),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16363_ (.RESET_B(net437),
    .D(net1491),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16364_ (.RESET_B(net438),
    .D(net1533),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16365_ (.RESET_B(net439),
    .D(net2556),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16366_ (.RESET_B(net440),
    .D(net1450),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_140_clk_regs));
 sg13g2_dfrbpq_1 _16367_ (.RESET_B(net441),
    .D(net1552),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16368_ (.RESET_B(net442),
    .D(net2509),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_143_clk_regs));
 sg13g2_dfrbpq_1 _16369_ (.RESET_B(net443),
    .D(net2524),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_136_clk_regs));
 sg13g2_dfrbpq_1 _16370_ (.RESET_B(net444),
    .D(net2619),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _16371_ (.RESET_B(net445),
    .D(net1524),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16372_ (.RESET_B(net446),
    .D(net1501),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16373_ (.RESET_B(net447),
    .D(net1507),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16374_ (.RESET_B(net448),
    .D(net2657),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_164_clk_regs));
 sg13g2_dfrbpq_1 _16375_ (.RESET_B(net449),
    .D(net1479),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_141_clk_regs));
 sg13g2_dfrbpq_1 _16376_ (.RESET_B(net450),
    .D(net1449),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16377_ (.RESET_B(net451),
    .D(_00049_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_138_clk_regs));
 sg13g2_dfrbpq_1 _16378_ (.RESET_B(net452),
    .D(_00050_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _16379_ (.RESET_B(net453),
    .D(_00051_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_163_clk_regs));
 sg13g2_dfrbpq_1 _16380_ (.RESET_B(net454),
    .D(_00052_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_2 _16381_ (.RESET_B(net455),
    .D(net1671),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_2 _16382_ (.RESET_B(net456),
    .D(net2739),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_2 _16383_ (.RESET_B(net457),
    .D(net2746),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_2 _16384_ (.RESET_B(net458),
    .D(net2747),
    .Q(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16385_ (.RESET_B(net459),
    .D(net2740),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_2 _16386_ (.RESET_B(net460),
    .D(net2734),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _16387_ (.RESET_B(net461),
    .D(net2729),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _16388_ (.RESET_B(net462),
    .D(net2707),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _16389_ (.RESET_B(net463),
    .D(net2699),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _16390_ (.RESET_B(net464),
    .D(net2673),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _16391_ (.RESET_B(net465),
    .D(net2694),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16392_ (.RESET_B(net466),
    .D(net2696),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16393_ (.RESET_B(net467),
    .D(net2681),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _16394_ (.RESET_B(net468),
    .D(net2683),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16395_ (.RESET_B(net469),
    .D(net2711),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16396_ (.RESET_B(net470),
    .D(net2690),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _16397_ (.RESET_B(net471),
    .D(net2685),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16398_ (.RESET_B(net472),
    .D(net2710),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16399_ (.RESET_B(net473),
    .D(net2706),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _16400_ (.RESET_B(net474),
    .D(net2701),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _16401_ (.RESET_B(net475),
    .D(net2738),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16402_ (.RESET_B(net476),
    .D(net2743),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16403_ (.RESET_B(net477),
    .D(net2741),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _16404_ (.RESET_B(net478),
    .D(net2742),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _16405_ (.RESET_B(net479),
    .D(net1673),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_2 _16406_ (.RESET_B(net480),
    .D(net2588),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_2 _16407_ (.RESET_B(net481),
    .D(net2656),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_2 _16408_ (.RESET_B(net489),
    .D(net2613),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16409_ (.RESET_B(net1232),
    .D(\i_tinyqv.cpu.i_core.cy_out ),
    .Q(\i_tinyqv.cpu.i_core.cy ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _16410_ (.RESET_B(net1231),
    .D(_00103_),
    .Q(\i_tinyqv.cpu.i_core.load_done ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _16411_ (.RESET_B(net1230),
    .D(_00104_),
    .Q(\i_tinyqv.cpu.i_core.cycle[0] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _16412_ (.RESET_B(net1228),
    .D(net3578),
    .Q(\i_tinyqv.cpu.i_core.cycle[1] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _16413_ (.RESET_B(net1226),
    .D(_00106_),
    .Q(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_1 _16414_ (.RESET_B(net1225),
    .D(_00107_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _16415_ (.RESET_B(net1223),
    .D(_00108_),
    .Q(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .CLK(clknet_leaf_168_clk_regs));
 sg13g2_dfrbpq_1 _16416_ (.RESET_B(net503),
    .D(net2998),
    .Q(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _16417_ (.RESET_B(net1221),
    .D(_00020_),
    .Q(\i_tinyqv.cpu.i_core.i_instrret.add ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _16418_ (.RESET_B(net1219),
    .D(net3781),
    .Q(\i_tinyqv.cpu.i_core.mcause[0] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16419_ (.RESET_B(net1217),
    .D(net3469),
    .Q(\i_tinyqv.cpu.i_core.mcause[1] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _16420_ (.RESET_B(net1215),
    .D(_00112_),
    .Q(\i_tinyqv.cpu.i_core.mcause[2] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _16421_ (.RESET_B(net1213),
    .D(_00113_),
    .Q(\i_tinyqv.cpu.i_core.mcause[3] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _16422_ (.RESET_B(net1211),
    .D(_00114_),
    .Q(\i_tinyqv.cpu.i_core.mcause[4] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_1 _16423_ (.RESET_B(net1209),
    .D(_00115_),
    .Q(\i_tinyqv.cpu.i_core.mcause[5] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_2 _16424_ (.RESET_B(net2487),
    .D(_00116_),
    .Q(_00074_),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _16425_ (.RESET_B(net1205),
    .D(net2838),
    .Q(\i_tinyqv.cpu.i_core.mepc[20] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16426_ (.RESET_B(net1203),
    .D(net2862),
    .Q(\i_tinyqv.cpu.i_core.mepc[21] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16427_ (.RESET_B(net1201),
    .D(net2860),
    .Q(\i_tinyqv.cpu.i_core.mepc[22] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _16428_ (.RESET_B(net1199),
    .D(net2829),
    .Q(\i_tinyqv.cpu.i_core.mepc[23] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _16429_ (.RESET_B(net1197),
    .D(net3130),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _16430_ (.RESET_B(net511),
    .D(net3141),
    .Q(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _16431_ (.RESET_B(net1196),
    .D(\i_tinyqv.cpu.i_core.cmp_out ),
    .Q(\i_tinyqv.cpu.i_core.cmp ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_1 _16432_ (.RESET_B(net1195),
    .D(net3098),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _16433_ (.RESET_B(net1193),
    .D(_00124_),
    .Q(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _16434_ (.RESET_B(net1191),
    .D(_00125_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_2 _16435_ (.RESET_B(net1190),
    .D(_00126_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_2 _16436_ (.RESET_B(net1189),
    .D(_00127_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_2 _16437_ (.RESET_B(net1188),
    .D(_00128_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_1 _16438_ (.RESET_B(net512),
    .D(net2782),
    .Q(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16439_ (.RESET_B(net513),
    .D(_00045_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_1 _16440_ (.RESET_B(net514),
    .D(net3641),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_1 _16441_ (.RESET_B(net515),
    .D(_00047_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _16442_ (.RESET_B(net516),
    .D(_00048_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .CLK(clknet_leaf_149_clk_regs));
 sg13g2_dfrbpq_2 _16443_ (.RESET_B(net517),
    .D(net1460),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.data[0] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_2 _16444_ (.RESET_B(net518),
    .D(net2554),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.data[1] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_2 _16445_ (.RESET_B(net519),
    .D(net1437),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.data[2] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_2 _16446_ (.RESET_B(net520),
    .D(net1557),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.data[3] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16447_ (.RESET_B(net521),
    .D(net1498),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[4] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16448_ (.RESET_B(net522),
    .D(net1660),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[5] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16449_ (.RESET_B(net523),
    .D(net2679),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[6] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16450_ (.RESET_B(net524),
    .D(net2638),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[7] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16451_ (.RESET_B(net525),
    .D(net1662),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[8] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16452_ (.RESET_B(net526),
    .D(net1577),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[9] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16453_ (.RESET_B(net527),
    .D(net1441),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[10] ),
    .CLK(clknet_leaf_99_clk_regs));
 sg13g2_dfrbpq_1 _16454_ (.RESET_B(net528),
    .D(net1452),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[11] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16455_ (.RESET_B(net529),
    .D(net2661),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[12] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16456_ (.RESET_B(net530),
    .D(net2521),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[13] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16457_ (.RESET_B(net531),
    .D(net1518),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[14] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _16458_ (.RESET_B(net532),
    .D(net1644),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[15] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16459_ (.RESET_B(net533),
    .D(net2599),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[16] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16460_ (.RESET_B(net534),
    .D(net1635),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[17] ),
    .CLK(clknet_leaf_100_clk_regs));
 sg13g2_dfrbpq_1 _16461_ (.RESET_B(net535),
    .D(net1502),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[18] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _16462_ (.RESET_B(net536),
    .D(net1542),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[19] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16463_ (.RESET_B(net537),
    .D(net2587),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[20] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16464_ (.RESET_B(net538),
    .D(net1526),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[21] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _16465_ (.RESET_B(net539),
    .D(net1659),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[22] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _16466_ (.RESET_B(net540),
    .D(net1670),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[23] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16467_ (.RESET_B(net541),
    .D(net1447),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[24] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16468_ (.RESET_B(net542),
    .D(net1547),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[25] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _16469_ (.RESET_B(net555),
    .D(net1563),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[26] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _16470_ (.RESET_B(net1187),
    .D(net2510),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[27] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_1 _16471_ (.RESET_B(net1185),
    .D(_00130_),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[0] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _16472_ (.RESET_B(net1184),
    .D(_00131_),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[1] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16473_ (.RESET_B(net1183),
    .D(_00132_),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[2] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16474_ (.RESET_B(net1182),
    .D(_00133_),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[3] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _16475_ (.RESET_B(net1181),
    .D(net3762),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.cy ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16476_ (.RESET_B(net1180),
    .D(net4039),
    .Q(\i_tinyqv.cpu.i_timer.cy ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _16477_ (.RESET_B(net1179),
    .D(net3974),
    .Q(\i_tinyqv.cpu.i_core.mip[16] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16478_ (.RESET_B(net1178),
    .D(_00137_),
    .Q(\i_tinyqv.cpu.i_timer.time_pulse_r ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _16479_ (.RESET_B(net1177),
    .D(_00138_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[12] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16480_ (.RESET_B(net1176),
    .D(_00139_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[13] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16481_ (.RESET_B(net1175),
    .D(_00140_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[14] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_1 _16482_ (.RESET_B(net556),
    .D(_00141_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[15] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16483_ (.RESET_B(net557),
    .D(net1672),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[4] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_2 _16484_ (.RESET_B(net558),
    .D(net2577),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[5] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_2 _16485_ (.RESET_B(net559),
    .D(net2684),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[6] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_2 _16486_ (.RESET_B(net560),
    .D(net1562),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[7] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _16487_ (.RESET_B(net561),
    .D(net1493),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[8] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16488_ (.RESET_B(net562),
    .D(net2579),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[9] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16489_ (.RESET_B(net563),
    .D(net2576),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[10] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16490_ (.RESET_B(net564),
    .D(net1442),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[11] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _16491_ (.RESET_B(net565),
    .D(net1631),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[12] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16492_ (.RESET_B(net566),
    .D(net2578),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[13] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16493_ (.RESET_B(net567),
    .D(net2615),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[14] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16494_ (.RESET_B(net568),
    .D(net2598),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[15] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _16495_ (.RESET_B(net569),
    .D(net2539),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[16] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16496_ (.RESET_B(net570),
    .D(net2625),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[17] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16497_ (.RESET_B(net571),
    .D(net2609),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[18] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_1 _16498_ (.RESET_B(net572),
    .D(net1568),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[19] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _16499_ (.RESET_B(net573),
    .D(net2565),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[20] ),
    .CLK(clknet_leaf_97_clk_regs));
 sg13g2_dfrbpq_1 _16500_ (.RESET_B(net574),
    .D(net2602),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[21] ),
    .CLK(clknet_leaf_98_clk_regs));
 sg13g2_dfrbpq_1 _16501_ (.RESET_B(net575),
    .D(net2590),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[22] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16502_ (.RESET_B(net576),
    .D(net2583),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[23] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _16503_ (.RESET_B(net577),
    .D(net2654),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[24] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _16504_ (.RESET_B(net578),
    .D(net1596),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[25] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16505_ (.RESET_B(net579),
    .D(net1448),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[26] ),
    .CLK(clknet_leaf_144_clk_regs));
 sg13g2_dfrbpq_1 _16506_ (.RESET_B(net580),
    .D(net1620),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[27] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _16507_ (.RESET_B(net581),
    .D(net1446),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[28] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16508_ (.RESET_B(net582),
    .D(net1621),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[29] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16509_ (.RESET_B(net583),
    .D(net2636),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[30] ),
    .CLK(clknet_leaf_160_clk_regs));
 sg13g2_dfrbpq_1 _16510_ (.RESET_B(net897),
    .D(net1589),
    .Q(\i_tinyqv.cpu.i_timer.mtimecmp[31] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _16511_ (.RESET_B(net1174),
    .D(net2278),
    .Q(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _16512_ (.RESET_B(net1173),
    .D(_00142_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[0] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _16513_ (.RESET_B(net1171),
    .D(_00143_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[1] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _16514_ (.RESET_B(net1169),
    .D(net3744),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[2] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _16515_ (.RESET_B(net1167),
    .D(_00145_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[3] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_2 _16516_ (.RESET_B(net1165),
    .D(_00146_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[4] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _16517_ (.RESET_B(net1163),
    .D(net3505),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[5] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_2 _16518_ (.RESET_B(net1161),
    .D(net3693),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[6] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_2 _16519_ (.RESET_B(net1159),
    .D(_00149_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[7] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _16520_ (.RESET_B(net1157),
    .D(net3680),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[8] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_2 _16521_ (.RESET_B(net1155),
    .D(_00151_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[9] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _16522_ (.RESET_B(net1153),
    .D(_00152_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[10] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_1 _16523_ (.RESET_B(net1151),
    .D(net3734),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[11] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _16524_ (.RESET_B(net1149),
    .D(net3663),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[12] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _16525_ (.RESET_B(net1146),
    .D(net3876),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[13] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _16526_ (.RESET_B(net1144),
    .D(net3851),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[14] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _16527_ (.RESET_B(net1142),
    .D(_00157_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[15] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _16528_ (.RESET_B(net1140),
    .D(net3856),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[16] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _16529_ (.RESET_B(net1138),
    .D(net3859),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[17] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _16530_ (.RESET_B(net1136),
    .D(_00160_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[18] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _16531_ (.RESET_B(net1134),
    .D(net3769),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[19] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _16532_ (.RESET_B(net1132),
    .D(net3791),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[20] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _16533_ (.RESET_B(net1130),
    .D(net3718),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[21] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _16534_ (.RESET_B(net1128),
    .D(_00164_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[22] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_1 _16535_ (.RESET_B(net1126),
    .D(_00165_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[23] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _16536_ (.RESET_B(net1124),
    .D(_00166_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[24] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _16537_ (.RESET_B(net1122),
    .D(net3906),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[25] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _16538_ (.RESET_B(net1120),
    .D(net3953),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[26] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _16539_ (.RESET_B(net1118),
    .D(_00169_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[27] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_1 _16540_ (.RESET_B(net1116),
    .D(_00170_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[28] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _16541_ (.RESET_B(net1114),
    .D(_00171_),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[29] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _16542_ (.RESET_B(net1112),
    .D(net3715),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[30] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _16543_ (.RESET_B(net1110),
    .D(net2836),
    .Q(\i_peripherals.i_user_peri39.math_result_reg[31] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _16544_ (.RESET_B(net1108),
    .D(_00174_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[0] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_2 _16545_ (.RESET_B(net1106),
    .D(_00175_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[1] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_1 _16546_ (.RESET_B(net1104),
    .D(net3842),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[2] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _16547_ (.RESET_B(net1102),
    .D(_00177_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[3] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_1 _16548_ (.RESET_B(net1100),
    .D(net3872),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[4] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_2 _16549_ (.RESET_B(net1098),
    .D(_00179_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[5] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _16550_ (.RESET_B(net1096),
    .D(net3804),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[6] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_2 _16551_ (.RESET_B(net1094),
    .D(_00181_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[7] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16552_ (.RESET_B(net1092),
    .D(_00182_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[8] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16553_ (.RESET_B(net1090),
    .D(_00183_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[9] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _16554_ (.RESET_B(net1088),
    .D(_00184_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[10] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16555_ (.RESET_B(net1086),
    .D(_00185_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[11] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _16556_ (.RESET_B(net1084),
    .D(_00186_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[12] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _16557_ (.RESET_B(net1082),
    .D(_00187_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[13] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16558_ (.RESET_B(net1080),
    .D(_00188_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[14] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _16559_ (.RESET_B(net1078),
    .D(_00189_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[15] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _16560_ (.RESET_B(net1076),
    .D(_00190_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[16] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16561_ (.RESET_B(net1074),
    .D(_00191_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[17] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16562_ (.RESET_B(net1072),
    .D(_00192_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[18] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16563_ (.RESET_B(net1070),
    .D(_00193_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[19] ),
    .CLK(clknet_leaf_86_clk_regs));
 sg13g2_dfrbpq_2 _16564_ (.RESET_B(net1068),
    .D(_00194_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[20] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_2 _16565_ (.RESET_B(net1066),
    .D(_00195_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[21] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _16566_ (.RESET_B(net1064),
    .D(net3004),
    .Q(\i_peripherals.i_user_peri39.instr[0] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16567_ (.RESET_B(net1062),
    .D(net3503),
    .Q(\i_peripherals.i_user_peri39.instr[1] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _16568_ (.RESET_B(net1060),
    .D(net3587),
    .Q(\i_peripherals.i_user_peri39.instr[2] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _16569_ (.RESET_B(net1058),
    .D(net3447),
    .Q(\i_peripherals.i_user_peri39.instr[3] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _16570_ (.RESET_B(net1056),
    .D(net3394),
    .Q(\i_peripherals.i_user_peri39.instr[4] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _16571_ (.RESET_B(net1054),
    .D(_00201_),
    .Q(\i_peripherals.i_user_peri39.instr[5] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _16572_ (.RESET_B(net1052),
    .D(net3550),
    .Q(\i_peripherals.i_user_peri39.instr[6] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_1 _16573_ (.RESET_B(net1050),
    .D(net3512),
    .Q(\i_peripherals.i_user_peri39.instr[7] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _16574_ (.RESET_B(net1048),
    .D(net2772),
    .Q(\i_peripherals.i_user_peri39.instr[8] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16575_ (.RESET_B(net1046),
    .D(net3464),
    .Q(\i_peripherals.i_user_peri39.instr[9] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _16576_ (.RESET_B(net1044),
    .D(net2752),
    .Q(\i_peripherals.i_user_peri39.instr[10] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _16577_ (.RESET_B(net1042),
    .D(net2780),
    .Q(\i_peripherals.i_user_peri39.instr[11] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_1 _16578_ (.RESET_B(net1040),
    .D(net2806),
    .Q(\i_peripherals.i_user_peri39.instr[12] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16579_ (.RESET_B(net1038),
    .D(_00209_),
    .Q(\i_peripherals.i_user_peri39.instr[13] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _16580_ (.RESET_B(net1036),
    .D(net3371),
    .Q(\i_peripherals.i_user_peri39.instr[14] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _16581_ (.RESET_B(net1034),
    .D(net3436),
    .Q(\i_peripherals.i_user_peri39.instr[15] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16582_ (.RESET_B(net1032),
    .D(net3675),
    .Q(\i_peripherals.i_user_peri39.instr[16] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _16583_ (.RESET_B(net1030),
    .D(net3481),
    .Q(\i_peripherals.i_user_peri39.instr[17] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16584_ (.RESET_B(net1028),
    .D(net3608),
    .Q(\i_peripherals.i_user_peri39.instr[18] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _16585_ (.RESET_B(net1026),
    .D(net3773),
    .Q(\i_peripherals.i_user_peri39.instr[19] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_2 _16586_ (.RESET_B(net1024),
    .D(net3748),
    .Q(\i_peripherals.i_user_peri39.instr[20] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16587_ (.RESET_B(net1022),
    .D(_00217_),
    .Q(\i_peripherals.i_user_peri39.instr[21] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_2 _16588_ (.RESET_B(net1020),
    .D(net3644),
    .Q(\i_peripherals.i_user_peri39.instr[22] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16589_ (.RESET_B(net1018),
    .D(net3592),
    .Q(\i_peripherals.i_user_peri39.instr[23] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16590_ (.RESET_B(net1016),
    .D(_00220_),
    .Q(\i_peripherals.i_user_peri39.instr[24] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _16591_ (.RESET_B(net1014),
    .D(_00221_),
    .Q(\i_peripherals.i_user_peri39.instr[25] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _16592_ (.RESET_B(net1012),
    .D(net3330),
    .Q(\i_peripherals.i_user_peri39.instr[26] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _16593_ (.RESET_B(net1010),
    .D(_00223_),
    .Q(\i_peripherals.i_user_peri39.instr[27] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _16594_ (.RESET_B(net1008),
    .D(_00224_),
    .Q(\i_peripherals.i_user_peri39.instr[28] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _16595_ (.RESET_B(net1006),
    .D(_00225_),
    .Q(\i_peripherals.i_user_peri39.instr[29] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _16596_ (.RESET_B(net1004),
    .D(_00226_),
    .Q(\i_peripherals.i_user_peri39.instr[30] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _16597_ (.RESET_B(net1002),
    .D(_00227_),
    .Q(\i_peripherals.i_user_peri39.instr[31] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _16598_ (.RESET_B(net1000),
    .D(_00228_),
    .Q(\i_peripherals.i_uart.i_uart_tx.txd_reg ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _16599_ (.RESET_B(net999),
    .D(_00229_),
    .Q(\i_peripherals.i_user_peri39._GEN[0] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _16600_ (.RESET_B(net998),
    .D(net3073),
    .Q(\i_peripherals.i_user_peri39._GEN[1] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _16601_ (.RESET_B(net997),
    .D(net2963),
    .Q(\i_peripherals.i_user_peri39._GEN[2] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _16602_ (.RESET_B(net996),
    .D(net3125),
    .Q(\i_peripherals.i_user_peri39._GEN[3] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _16603_ (.RESET_B(net995),
    .D(net3031),
    .Q(\i_peripherals.i_user_peri39._GEN[100] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _16604_ (.RESET_B(net994),
    .D(_00234_),
    .Q(\i_peripherals.i_user_peri39._GEN[101] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _16605_ (.RESET_B(net993),
    .D(net2996),
    .Q(\i_peripherals.i_user_peri39._GEN[102] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _16606_ (.RESET_B(net992),
    .D(net2923),
    .Q(\i_peripherals.i_user_peri39._GEN[103] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _16607_ (.RESET_B(net991),
    .D(net3585),
    .Q(\i_peripherals.i_user_peri39._GEN[104] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _16608_ (.RESET_B(net990),
    .D(net2994),
    .Q(\i_peripherals.i_user_peri39._GEN[105] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _16609_ (.RESET_B(net989),
    .D(net3564),
    .Q(\i_peripherals.i_user_peri39._GEN[106] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _16610_ (.RESET_B(net988),
    .D(net3560),
    .Q(\i_peripherals.i_user_peri39._GEN[107] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _16611_ (.RESET_B(net987),
    .D(net3635),
    .Q(\i_peripherals.i_user_peri39._GEN[108] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _16612_ (.RESET_B(net986),
    .D(net2978),
    .Q(\i_peripherals.i_user_peri39._GEN[109] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _16613_ (.RESET_B(net985),
    .D(net3027),
    .Q(\i_peripherals.i_user_peri39._GEN[110] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _16614_ (.RESET_B(net984),
    .D(net3109),
    .Q(\i_peripherals.i_user_peri39._GEN[111] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16615_ (.RESET_B(net983),
    .D(net2927),
    .Q(\i_peripherals.i_user_peri39._GEN[112] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_2 _16616_ (.RESET_B(net982),
    .D(net3086),
    .Q(\i_peripherals.i_user_peri39._GEN[113] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_2 _16617_ (.RESET_B(net981),
    .D(net2873),
    .Q(\i_peripherals.i_user_peri39._GEN[114] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _16618_ (.RESET_B(net980),
    .D(net3002),
    .Q(\i_peripherals.i_user_peri39._GEN[115] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _16619_ (.RESET_B(net979),
    .D(net3684),
    .Q(\i_peripherals.i_user_peri39._GEN[116] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _16620_ (.RESET_B(net978),
    .D(net2952),
    .Q(\i_peripherals.i_user_peri39._GEN[117] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _16621_ (.RESET_B(net977),
    .D(net3151),
    .Q(\i_peripherals.i_user_peri39._GEN[118] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _16622_ (.RESET_B(net976),
    .D(net3012),
    .Q(\i_peripherals.i_user_peri39._GEN[119] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_2 _16623_ (.RESET_B(net975),
    .D(net2940),
    .Q(\i_peripherals.i_user_peri39._GEN[120] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_1 _16624_ (.RESET_B(net974),
    .D(_00254_),
    .Q(\i_peripherals.i_user_peri39._GEN[121] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_2 _16625_ (.RESET_B(net973),
    .D(net2887),
    .Q(\i_peripherals.i_user_peri39._GEN[122] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _16626_ (.RESET_B(net972),
    .D(net2925),
    .Q(\i_peripherals.i_user_peri39._GEN[123] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16627_ (.RESET_B(net971),
    .D(net2980),
    .Q(\i_peripherals.i_user_peri39._GEN[124] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _16628_ (.RESET_B(net958),
    .D(net2934),
    .Q(\i_peripherals.i_user_peri39._GEN[125] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16629_ (.RESET_B(net957),
    .D(net2919),
    .Q(\i_peripherals.i_user_peri39._GEN[126] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _16630_ (.RESET_B(net956),
    .D(net3052),
    .Q(\i_peripherals.i_user_peri39._GEN[127] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16631_ (.RESET_B(net955),
    .D(_00261_),
    .Q(\i_peripherals.i_user_peri39._GEN[32] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _16632_ (.RESET_B(net954),
    .D(net3034),
    .Q(\i_peripherals.i_user_peri39._GEN[33] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _16633_ (.RESET_B(net953),
    .D(net3048),
    .Q(\i_peripherals.i_user_peri39._GEN[34] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _16634_ (.RESET_B(net952),
    .D(net3037),
    .Q(\i_peripherals.i_user_peri39._GEN[35] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _16635_ (.RESET_B(net951),
    .D(net3041),
    .Q(\i_peripherals.i_user_peri39._GEN[36] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _16636_ (.RESET_B(net950),
    .D(_00266_),
    .Q(\i_peripherals.i_user_peri39._GEN[37] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_2 _16637_ (.RESET_B(net949),
    .D(net3153),
    .Q(\i_peripherals.i_user_peri39._GEN[38] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _16638_ (.RESET_B(net948),
    .D(net2905),
    .Q(\i_peripherals.i_user_peri39._GEN[39] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _16639_ (.RESET_B(net947),
    .D(net3610),
    .Q(\i_peripherals.i_user_peri39._GEN[40] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _16640_ (.RESET_B(net946),
    .D(net2971),
    .Q(\i_peripherals.i_user_peri39._GEN[41] ),
    .CLK(clknet_leaf_77_clk_regs));
 sg13g2_dfrbpq_2 _16641_ (.RESET_B(net945),
    .D(net3557),
    .Q(\i_peripherals.i_user_peri39._GEN[42] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _16642_ (.RESET_B(net944),
    .D(net3589),
    .Q(\i_peripherals.i_user_peri39._GEN[43] ),
    .CLK(clknet_leaf_83_clk_regs));
 sg13g2_dfrbpq_2 _16643_ (.RESET_B(net943),
    .D(net3669),
    .Q(\i_peripherals.i_user_peri39._GEN[44] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_1 _16644_ (.RESET_B(net942),
    .D(net3029),
    .Q(\i_peripherals.i_user_peri39._GEN[45] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _16645_ (.RESET_B(net941),
    .D(net2965),
    .Q(\i_peripherals.i_user_peri39._GEN[46] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _16646_ (.RESET_B(net940),
    .D(net3067),
    .Q(\i_peripherals.i_user_peri39._GEN[47] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16647_ (.RESET_B(net939),
    .D(net2823),
    .Q(\i_peripherals.i_user_peri39._GEN[48] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_2 _16648_ (.RESET_B(net938),
    .D(net2866),
    .Q(\i_peripherals.i_user_peri39._GEN[49] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _16649_ (.RESET_B(net937),
    .D(net2961),
    .Q(\i_peripherals.i_user_peri39._GEN[50] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_1 _16650_ (.RESET_B(net936),
    .D(net2982),
    .Q(\i_peripherals.i_user_peri39._GEN[51] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _16651_ (.RESET_B(net935),
    .D(net3736),
    .Q(\i_peripherals.i_user_peri39._GEN[52] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _16652_ (.RESET_B(net934),
    .D(net2912),
    .Q(\i_peripherals.i_user_peri39._GEN[53] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _16653_ (.RESET_B(net933),
    .D(net2984),
    .Q(\i_peripherals.i_user_peri39._GEN[54] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _16654_ (.RESET_B(net932),
    .D(net3014),
    .Q(\i_peripherals.i_user_peri39._GEN[55] ),
    .CLK(clknet_leaf_73_clk_regs));
 sg13g2_dfrbpq_2 _16655_ (.RESET_B(net931),
    .D(net2850),
    .Q(\i_peripherals.i_user_peri39._GEN[56] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _16656_ (.RESET_B(net930),
    .D(net2818),
    .Q(\i_peripherals.i_user_peri39._GEN[57] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _16657_ (.RESET_B(net929),
    .D(net2973),
    .Q(\i_peripherals.i_user_peri39._GEN[58] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _16658_ (.RESET_B(net928),
    .D(net2901),
    .Q(\i_peripherals.i_user_peri39._GEN[59] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16659_ (.RESET_B(net927),
    .D(net2956),
    .Q(\i_peripherals.i_user_peri39._GEN[60] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _16660_ (.RESET_B(net926),
    .D(net2988),
    .Q(\i_peripherals.i_user_peri39._GEN[61] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _16661_ (.RESET_B(net902),
    .D(net2854),
    .Q(\i_peripherals.i_user_peri39._GEN[62] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _16662_ (.RESET_B(net901),
    .D(net2899),
    .Q(\i_peripherals.i_user_peri39._GEN[63] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_2 _16663_ (.RESET_B(net896),
    .D(net3023),
    .Q(\i_peripherals.i_user_peri39.busy_counter[0] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _16664_ (.RESET_B(net894),
    .D(net3703),
    .Q(\i_peripherals.i_user_peri39.busy_counter[1] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_1 _16665_ (.RESET_B(net892),
    .D(net3167),
    .Q(\i_tinyqv.cpu.instr_data[3][0] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _16666_ (.RESET_B(net891),
    .D(net2990),
    .Q(\i_tinyqv.cpu.instr_data[3][1] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _16667_ (.RESET_B(net890),
    .D(net3200),
    .Q(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _16668_ (.RESET_B(net888),
    .D(net3293),
    .Q(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _16669_ (.RESET_B(net886),
    .D(net3214),
    .Q(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_2 _16670_ (.RESET_B(net884),
    .D(net3898),
    .Q(\i_peripherals.i_uart.baud_divider[0] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _16671_ (.RESET_B(net882),
    .D(net3939),
    .Q(\i_peripherals.i_uart.baud_divider[1] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _16672_ (.RESET_B(net880),
    .D(net3878),
    .Q(\i_peripherals.i_uart.baud_divider[2] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16673_ (.RESET_B(net878),
    .D(net3935),
    .Q(\i_peripherals.i_uart.baud_divider[3] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16674_ (.RESET_B(net876),
    .D(net3987),
    .Q(\i_peripherals.i_uart.baud_divider[4] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16675_ (.RESET_B(net874),
    .D(_00305_),
    .Q(\i_peripherals.i_uart.baud_divider[5] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16676_ (.RESET_B(net872),
    .D(net4016),
    .Q(\i_peripherals.i_uart.baud_divider[6] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_2 _16677_ (.RESET_B(net870),
    .D(net3922),
    .Q(\i_peripherals.i_uart.baud_divider[7] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _16678_ (.RESET_B(net868),
    .D(_00308_),
    .Q(\i_peripherals.data_ready_r ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16679_ (.RESET_B(net867),
    .D(_00309_),
    .Q(\i_peripherals.i_uart.uart_rx_buffered ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16680_ (.RESET_B(net866),
    .D(net3064),
    .Q(\i_peripherals.i_uart.rxd_select ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16681_ (.RESET_B(net864),
    .D(net3764),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[0] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16682_ (.RESET_B(net862),
    .D(net3450),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[1] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16683_ (.RESET_B(net860),
    .D(net3300),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[2] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16684_ (.RESET_B(net858),
    .D(net3548),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[3] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16685_ (.RESET_B(net856),
    .D(_00315_),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[4] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16686_ (.RESET_B(net854),
    .D(net3390),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[5] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16687_ (.RESET_B(net852),
    .D(net3401),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[6] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16688_ (.RESET_B(net850),
    .D(net3459),
    .Q(\i_peripherals.i_uart.i_uart_tx.data_to_send[7] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16689_ (.RESET_B(net848),
    .D(net3218),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[0] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _16690_ (.RESET_B(net846),
    .D(_00320_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[1] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _16691_ (.RESET_B(net844),
    .D(_00321_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[2] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _16692_ (.RESET_B(net842),
    .D(net3070),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[3] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _16693_ (.RESET_B(net840),
    .D(_00323_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[4] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _16694_ (.RESET_B(net838),
    .D(net3251),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[5] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_1 _16695_ (.RESET_B(net836),
    .D(_00325_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[6] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16696_ (.RESET_B(net834),
    .D(net3290),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[7] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _16697_ (.RESET_B(net832),
    .D(_00327_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[8] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _16698_ (.RESET_B(net830),
    .D(net3274),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[9] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _16699_ (.RESET_B(net828),
    .D(_00329_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[10] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _16700_ (.RESET_B(net826),
    .D(_00330_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[11] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _16701_ (.RESET_B(net824),
    .D(_00331_),
    .Q(\i_peripherals.i_uart.i_uart_tx.cycle_counter[12] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _16702_ (.RESET_B(net822),
    .D(_00332_),
    .Q(\i_peripherals.i_uart.i_uart_tx.fsm_state[0] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _16703_ (.RESET_B(net820),
    .D(net2885),
    .Q(\i_peripherals.i_uart.i_uart_tx.fsm_state[1] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _16704_ (.RESET_B(net818),
    .D(_00334_),
    .Q(\i_peripherals.i_uart.i_uart_tx.fsm_state[2] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_2 _16705_ (.RESET_B(net816),
    .D(_00335_),
    .Q(\i_peripherals.i_uart.i_uart_tx.fsm_state[3] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _16706_ (.RESET_B(net814),
    .D(_00336_),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[0] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _16707_ (.RESET_B(net813),
    .D(_00337_),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[1] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _16708_ (.RESET_B(net812),
    .D(net3360),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[2] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16709_ (.RESET_B(net811),
    .D(_00339_),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[3] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16710_ (.RESET_B(net810),
    .D(net3427),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[4] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16711_ (.RESET_B(net809),
    .D(_00341_),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[5] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _16712_ (.RESET_B(net808),
    .D(_00342_),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[6] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _16713_ (.RESET_B(net807),
    .D(_00343_),
    .Q(\i_peripherals.i_uart.i_uart_rx.recieved_data[7] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16714_ (.RESET_B(net806),
    .D(net2897),
    .Q(\i_peripherals.i_uart.i_uart_rx.bit_sample ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _16715_ (.RESET_B(net804),
    .D(_00345_),
    .Q(\i_peripherals.i_uart.i_uart_rx.uart_rts ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _16716_ (.RESET_B(net803),
    .D(_00346_),
    .Q(\i_peripherals.i_uart.i_uart_rx.fsm_state[0] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_2 _16717_ (.RESET_B(net801),
    .D(_00347_),
    .Q(\i_peripherals.i_uart.i_uart_rx.fsm_state[1] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _16718_ (.RESET_B(net799),
    .D(net3837),
    .Q(\i_peripherals.i_uart.i_uart_rx.fsm_state[2] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _16719_ (.RESET_B(net797),
    .D(_00349_),
    .Q(\i_peripherals.i_uart.i_uart_rx.fsm_state[3] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _16720_ (.RESET_B(net795),
    .D(net3105),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[0] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16721_ (.RESET_B(net794),
    .D(_00351_),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[1] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _16722_ (.RESET_B(net793),
    .D(net3253),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[2] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16723_ (.RESET_B(net792),
    .D(net3298),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[3] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16724_ (.RESET_B(net791),
    .D(net3248),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[4] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16725_ (.RESET_B(net790),
    .D(net3179),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[5] ),
    .CLK(clknet_leaf_49_clk_regs));
 sg13g2_dfrbpq_1 _16726_ (.RESET_B(net789),
    .D(_00356_),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[6] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_1 _16727_ (.RESET_B(net788),
    .D(_00357_),
    .Q(\i_peripherals.i_uart.uart_rx_buf_data[7] ),
    .CLK(clknet_leaf_48_clk_regs));
 sg13g2_dfrbpq_2 _16728_ (.RESET_B(net787),
    .D(_00358_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[0] ),
    .CLK(clknet_leaf_50_clk_regs));
 sg13g2_dfrbpq_2 _16729_ (.RESET_B(net786),
    .D(_00359_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16730_ (.RESET_B(net785),
    .D(net2976),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[2] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16731_ (.RESET_B(net784),
    .D(_00361_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[3] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16732_ (.RESET_B(net783),
    .D(net3520),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[4] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16733_ (.RESET_B(net782),
    .D(_00363_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16734_ (.RESET_B(net781),
    .D(net3193),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[6] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16735_ (.RESET_B(net780),
    .D(_00365_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[7] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16736_ (.RESET_B(net779),
    .D(_00366_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[8] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _16737_ (.RESET_B(net778),
    .D(_00367_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[9] ),
    .CLK(clknet_leaf_75_clk_regs));
 sg13g2_dfrbpq_2 _16738_ (.RESET_B(net777),
    .D(net3017),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[10] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _16739_ (.RESET_B(net776),
    .D(_00369_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[11] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_1 _16740_ (.RESET_B(net775),
    .D(_00370_),
    .Q(\i_peripherals.i_uart.i_uart_rx.cycle_counter[12] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _16741_ (.RESET_B(net774),
    .D(net3055),
    .Q(\i_peripherals.gpio_out[0] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _16742_ (.RESET_B(net772),
    .D(net2967),
    .Q(\i_peripherals.gpio_out[1] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _16743_ (.RESET_B(net770),
    .D(net3094),
    .Q(\i_peripherals.gpio_out[2] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _16744_ (.RESET_B(net768),
    .D(net3267),
    .Q(\i_peripherals.gpio_out[3] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _16745_ (.RESET_B(net766),
    .D(net3137),
    .Q(\i_peripherals.gpio_out[4] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_2 _16746_ (.RESET_B(net764),
    .D(net3265),
    .Q(\i_peripherals.gpio_out[5] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_2 _16747_ (.RESET_B(net762),
    .D(net3188),
    .Q(\i_peripherals.gpio_out[6] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16748_ (.RESET_B(net760),
    .D(net2947),
    .Q(\i_peripherals.gpio_out[7] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16749_ (.RESET_B(net758),
    .D(net2942),
    .Q(\i_peripherals.func_sel[0] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16750_ (.RESET_B(net756),
    .D(net3418),
    .Q(\i_peripherals.func_sel[1] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16751_ (.RESET_B(net754),
    .D(net3092),
    .Q(\i_peripherals.func_sel[2] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16752_ (.RESET_B(net752),
    .D(net2770),
    .Q(\i_peripherals.func_sel[3] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _16753_ (.RESET_B(net750),
    .D(net2893),
    .Q(\i_peripherals.func_sel[4] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _16754_ (.RESET_B(net748),
    .D(net2774),
    .Q(\i_peripherals.func_sel[5] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _16755_ (.RESET_B(net746),
    .D(net3626),
    .Q(\i_peripherals.data_out[0] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _16756_ (.RESET_B(net744),
    .D(_00386_),
    .Q(\i_peripherals.data_out[1] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _16757_ (.RESET_B(net742),
    .D(net3478),
    .Q(\i_peripherals.data_out[2] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_2 _16758_ (.RESET_B(net740),
    .D(_00388_),
    .Q(\i_peripherals.data_out[3] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _16759_ (.RESET_B(net738),
    .D(_00389_),
    .Q(\i_peripherals.data_out[4] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _16760_ (.RESET_B(net736),
    .D(_00390_),
    .Q(\i_peripherals.data_out[5] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _16761_ (.RESET_B(net734),
    .D(net3475),
    .Q(\i_peripherals.data_out[6] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16762_ (.RESET_B(net732),
    .D(_00392_),
    .Q(\i_peripherals.data_out[7] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16763_ (.RESET_B(net730),
    .D(net3353),
    .Q(\i_peripherals.data_out[8] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _16764_ (.RESET_B(net728),
    .D(net3739),
    .Q(\i_peripherals.data_out[9] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _16765_ (.RESET_B(net726),
    .D(net3606),
    .Q(\i_peripherals.data_out[10] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _16766_ (.RESET_B(net724),
    .D(net3823),
    .Q(\i_peripherals.data_out[11] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16767_ (.RESET_B(net722),
    .D(_00397_),
    .Q(\i_peripherals.data_out[12] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _16768_ (.RESET_B(net720),
    .D(_00398_),
    .Q(\i_peripherals.data_out[13] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16769_ (.RESET_B(net718),
    .D(_00399_),
    .Q(\i_peripherals.data_out[14] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16770_ (.RESET_B(net716),
    .D(_00400_),
    .Q(\i_peripherals.data_out[15] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16771_ (.RESET_B(net714),
    .D(_00401_),
    .Q(\i_peripherals.data_out[16] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _16772_ (.RESET_B(net712),
    .D(_00402_),
    .Q(\i_peripherals.data_out[17] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _16773_ (.RESET_B(net710),
    .D(_00403_),
    .Q(\i_peripherals.data_out[18] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _16774_ (.RESET_B(net708),
    .D(_00404_),
    .Q(\i_peripherals.data_out[19] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _16775_ (.RESET_B(net706),
    .D(_00405_),
    .Q(\i_peripherals.data_out[20] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _16776_ (.RESET_B(net704),
    .D(_00406_),
    .Q(\i_peripherals.data_out[21] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _16777_ (.RESET_B(net702),
    .D(_00407_),
    .Q(\i_peripherals.data_out[22] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_1 _16778_ (.RESET_B(net700),
    .D(_00408_),
    .Q(\i_peripherals.data_out[23] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _16779_ (.RESET_B(net698),
    .D(_00409_),
    .Q(\i_peripherals.data_out[24] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16780_ (.RESET_B(net696),
    .D(_00410_),
    .Q(\i_peripherals.data_out[25] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_1 _16781_ (.RESET_B(net694),
    .D(_00411_),
    .Q(\i_peripherals.data_out[26] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _16782_ (.RESET_B(net692),
    .D(_00412_),
    .Q(\i_peripherals.data_out[27] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16783_ (.RESET_B(net690),
    .D(_00413_),
    .Q(\i_peripherals.data_out[28] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_1 _16784_ (.RESET_B(net688),
    .D(_00414_),
    .Q(\i_peripherals.data_out[29] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_1 _16785_ (.RESET_B(net686),
    .D(_00415_),
    .Q(\i_peripherals.data_out[30] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_1 _16786_ (.RESET_B(net684),
    .D(_00416_),
    .Q(\i_peripherals.data_out[31] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _16787_ (.RESET_B(net682),
    .D(_00417_),
    .Q(\i_peripherals.data_out_hold ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_1 _16788_ (.RESET_B(net680),
    .D(net3696),
    .Q(debug_uart_txd),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _16789_ (.RESET_B(net679),
    .D(net3296),
    .Q(\i_debug_uart_tx.data_to_send[0] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _16790_ (.RESET_B(net677),
    .D(net3546),
    .Q(\i_debug_uart_tx.data_to_send[1] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _16791_ (.RESET_B(net675),
    .D(_00421_),
    .Q(\i_debug_uart_tx.data_to_send[2] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _16792_ (.RESET_B(net673),
    .D(_00422_),
    .Q(\i_debug_uart_tx.data_to_send[3] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _16793_ (.RESET_B(net671),
    .D(net3797),
    .Q(\i_debug_uart_tx.data_to_send[4] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _16794_ (.RESET_B(net669),
    .D(_00424_),
    .Q(\i_debug_uart_tx.data_to_send[5] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _16795_ (.RESET_B(net667),
    .D(net4083),
    .Q(\i_debug_uart_tx.data_to_send[6] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _16796_ (.RESET_B(net665),
    .D(net2795),
    .Q(\i_debug_uart_tx.data_to_send[7] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _16797_ (.RESET_B(net663),
    .D(_00427_),
    .Q(\i_debug_uart_tx.cycle_counter[0] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _16798_ (.RESET_B(net661),
    .D(_00428_),
    .Q(\i_debug_uart_tx.cycle_counter[1] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _16799_ (.RESET_B(net659),
    .D(_00429_),
    .Q(\i_debug_uart_tx.cycle_counter[2] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _16800_ (.RESET_B(net657),
    .D(_00430_),
    .Q(\i_debug_uart_tx.cycle_counter[3] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _16801_ (.RESET_B(net655),
    .D(net2745),
    .Q(\i_debug_uart_tx.cycle_counter[4] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_2 _16802_ (.RESET_B(net653),
    .D(net3989),
    .Q(\i_debug_uart_tx.fsm_state[0] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _16803_ (.RESET_B(net651),
    .D(net3184),
    .Q(\i_debug_uart_tx.fsm_state[1] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _16804_ (.RESET_B(net649),
    .D(net3958),
    .Q(\i_debug_uart_tx.fsm_state[2] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_2 _16805_ (.RESET_B(net647),
    .D(net3367),
    .Q(\i_debug_uart_tx.fsm_state[3] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _16806_ (.RESET_B(net645),
    .D(_00436_),
    .Q(\i_tinyqv.cpu.i_core.mie[11] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _16807_ (.RESET_B(net643),
    .D(net2856),
    .Q(\i_tinyqv.cpu.i_core.mie[10] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _16808_ (.RESET_B(net641),
    .D(net2895),
    .Q(\i_tinyqv.cpu.i_core.mie[9] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16809_ (.RESET_B(net639),
    .D(_00439_),
    .Q(\i_tinyqv.cpu.i_core.mie[8] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _16810_ (.RESET_B(net637),
    .D(_00440_),
    .Q(\i_tinyqv.cpu.i_core.mie[7] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16811_ (.RESET_B(net635),
    .D(_00441_),
    .Q(\i_tinyqv.cpu.i_core.mie[6] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _16812_ (.RESET_B(net633),
    .D(_00442_),
    .Q(\i_tinyqv.cpu.i_core.mie[5] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16813_ (.RESET_B(net631),
    .D(_00443_),
    .Q(\i_tinyqv.cpu.i_core.mie[4] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_2 _16814_ (.RESET_B(net629),
    .D(_00444_),
    .Q(\i_tinyqv.cpu.i_core.mie[3] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16815_ (.RESET_B(net627),
    .D(_00445_),
    .Q(\i_tinyqv.cpu.i_core.mie[2] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16816_ (.RESET_B(net625),
    .D(_00446_),
    .Q(\i_tinyqv.cpu.i_core.mie[1] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_2 _16817_ (.RESET_B(net623),
    .D(_00447_),
    .Q(\i_tinyqv.cpu.i_core.mie[0] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_2 _16818_ (.RESET_B(net621),
    .D(_00448_),
    .Q(\i_tinyqv.cpu.i_core.mie[16] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_2 _16819_ (.RESET_B(net619),
    .D(_00449_),
    .Q(\i_tinyqv.cpu.i_core.mip[1] ),
    .CLK(clknet_leaf_171_clk_regs));
 sg13g2_dfrbpq_2 _16820_ (.RESET_B(net617),
    .D(_00450_),
    .Q(\i_tinyqv.cpu.i_core.mip[0] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _16821_ (.RESET_B(net615),
    .D(_00451_),
    .Q(\i_tinyqv.cpu.i_core.mie[15] ),
    .CLK(clknet_leaf_169_clk_regs));
 sg13g2_dfrbpq_1 _16822_ (.RESET_B(net613),
    .D(_00452_),
    .Q(\i_tinyqv.cpu.i_core.mie[14] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _16823_ (.RESET_B(net611),
    .D(_00453_),
    .Q(\i_tinyqv.cpu.i_core.mie[13] ),
    .CLK(clknet_leaf_170_clk_regs));
 sg13g2_dfrbpq_1 _16824_ (.RESET_B(net898),
    .D(_00454_),
    .Q(\i_tinyqv.cpu.i_core.mie[12] ),
    .CLK(clknet_leaf_174_clk_regs));
 sg13g2_dfrbpq_1 _16825_ (.RESET_B(net899),
    .D(\debug_rd[0] ),
    .Q(\debug_rd_r[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _16826_ (.RESET_B(net900),
    .D(\debug_rd[1] ),
    .Q(\debug_rd_r[1] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _16827_ (.RESET_B(net903),
    .D(\debug_rd[2] ),
    .Q(\debug_rd_r[2] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _16828_ (.RESET_B(net609),
    .D(\debug_rd[3] ),
    .Q(\debug_rd_r[3] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_1 _16829_ (.RESET_B(net607),
    .D(_00455_),
    .Q(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _16830_ (.RESET_B(net904),
    .D(net3864),
    .Q(debug_register_data),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_2 _16831_ (.RESET_B(net905),
    .D(net3880),
    .Q(\gpio_out_sel[6] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_2 _16832_ (.RESET_B(net906),
    .D(net4131),
    .Q(\gpio_out_sel[7] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _16833_ (.RESET_B(net907),
    .D(net4120),
    .Q(\time_limit[2] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _16834_ (.RESET_B(net908),
    .D(net4103),
    .Q(\time_limit[3] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _16835_ (.RESET_B(net909),
    .D(net4123),
    .Q(\time_limit[4] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _16836_ (.RESET_B(net910),
    .D(net4092),
    .Q(\time_limit[5] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _16837_ (.RESET_B(net911),
    .D(net3783),
    .Q(\time_limit[6] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16838_ (.RESET_B(net912),
    .D(net2),
    .Q(\ui_in_sync0[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _16839_ (.RESET_B(net913),
    .D(net3),
    .Q(\ui_in_sync0[1] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _16840_ (.RESET_B(net914),
    .D(net4),
    .Q(\ui_in_sync0[2] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16841_ (.RESET_B(net915),
    .D(net5),
    .Q(\ui_in_sync0[3] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16842_ (.RESET_B(net916),
    .D(net6),
    .Q(\ui_in_sync0[4] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _16843_ (.RESET_B(net917),
    .D(net7),
    .Q(\ui_in_sync0[5] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _16844_ (.RESET_B(net918),
    .D(net8),
    .Q(\ui_in_sync0[6] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _16845_ (.RESET_B(net919),
    .D(net9),
    .Q(\ui_in_sync0[7] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_2 _16846_ (.RESET_B(net920),
    .D(net2633),
    .Q(\i_peripherals.i_uart.ui_in[0] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_2 _16847_ (.RESET_B(net921),
    .D(net1599),
    .Q(\i_peripherals.i_uart.ui_in[1] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _16848_ (.RESET_B(net922),
    .D(net2668),
    .Q(\i_peripherals.i_uart.ui_in[2] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _16849_ (.RESET_B(net923),
    .D(net1600),
    .Q(\i_peripherals.i_uart.ui_in[3] ),
    .CLK(clknet_leaf_47_clk_regs));
 sg13g2_dfrbpq_1 _16850_ (.RESET_B(net924),
    .D(net1539),
    .Q(\i_peripherals.i_uart.ui_in[4] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _16851_ (.RESET_B(net925),
    .D(net1571),
    .Q(\i_peripherals.i_uart.ui_in[5] ),
    .CLK(clknet_leaf_44_clk_regs));
 sg13g2_dfrbpq_1 _16852_ (.RESET_B(net959),
    .D(net2553),
    .Q(\i_peripherals.i_uart.ui_in[6] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _16853_ (.RESET_B(net606),
    .D(net1564),
    .Q(\i_peripherals.i_uart.ui_in[7] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _16854_ (.RESET_B(net605),
    .D(net1),
    .Q(\i_debug_uart_tx.resetn ),
    .CLK(net1434));
 sg13g2_dfrbpq_1 _16855_ (.RESET_B(net604),
    .D(net3466),
    .Q(\i_tinyqv.cpu.instr_data[0][2] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _16856_ (.RESET_B(net603),
    .D(net3491),
    .Q(\i_tinyqv.cpu.instr_data[0][3] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _16857_ (.RESET_B(net602),
    .D(_00459_),
    .Q(\i_tinyqv.cpu.instr_data[0][4] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _16858_ (.RESET_B(net601),
    .D(net3462),
    .Q(\i_tinyqv.cpu.instr_data[0][5] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16859_ (.RESET_B(net600),
    .D(net3364),
    .Q(\i_tinyqv.cpu.instr_data[0][6] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _16860_ (.RESET_B(net599),
    .D(net3084),
    .Q(\i_tinyqv.cpu.instr_data[0][7] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _16861_ (.RESET_B(net598),
    .D(net3233),
    .Q(\i_tinyqv.cpu.instr_data[0][8] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _16862_ (.RESET_B(net597),
    .D(net3146),
    .Q(\i_tinyqv.cpu.instr_data[0][9] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16863_ (.RESET_B(net596),
    .D(net3082),
    .Q(\i_tinyqv.cpu.instr_data[0][10] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _16864_ (.RESET_B(net595),
    .D(net3118),
    .Q(\i_tinyqv.cpu.instr_data[0][11] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16865_ (.RESET_B(net594),
    .D(net3598),
    .Q(\i_tinyqv.cpu.instr_data[0][12] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _16866_ (.RESET_B(net593),
    .D(net3148),
    .Q(\i_tinyqv.cpu.instr_data[0][13] ),
    .CLK(clknet_leaf_95_clk_regs));
 sg13g2_dfrbpq_1 _16867_ (.RESET_B(net592),
    .D(net3162),
    .Q(\i_tinyqv.cpu.instr_data[0][14] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _16868_ (.RESET_B(net591),
    .D(net3413),
    .Q(\i_tinyqv.cpu.instr_data[0][15] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _16869_ (.RESET_B(net590),
    .D(net3408),
    .Q(\i_tinyqv.cpu.instr_data[3][2] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _16870_ (.RESET_B(net589),
    .D(net3572),
    .Q(\i_tinyqv.cpu.instr_data[3][3] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _16871_ (.RESET_B(net588),
    .D(net2814),
    .Q(\i_tinyqv.cpu.instr_data[3][4] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _16872_ (.RESET_B(net587),
    .D(net3654),
    .Q(\i_tinyqv.cpu.instr_data[3][5] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16873_ (.RESET_B(net586),
    .D(net3362),
    .Q(\i_tinyqv.cpu.instr_data[3][6] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _16874_ (.RESET_B(net585),
    .D(net2831),
    .Q(\i_tinyqv.cpu.instr_data[3][7] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _16875_ (.RESET_B(net584),
    .D(net3526),
    .Q(\i_tinyqv.cpu.instr_data[3][8] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16876_ (.RESET_B(net554),
    .D(net2864),
    .Q(\i_tinyqv.cpu.instr_data[3][9] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _16877_ (.RESET_B(net553),
    .D(net2799),
    .Q(\i_tinyqv.cpu.instr_data[3][10] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _16878_ (.RESET_B(net552),
    .D(net2786),
    .Q(\i_tinyqv.cpu.instr_data[3][11] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _16879_ (.RESET_B(net551),
    .D(net3392),
    .Q(\i_tinyqv.cpu.instr_data[3][12] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _16880_ (.RESET_B(net550),
    .D(net2793),
    .Q(\i_tinyqv.cpu.instr_data[3][13] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _16881_ (.RESET_B(net549),
    .D(net2844),
    .Q(\i_tinyqv.cpu.instr_data[3][14] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _16882_ (.RESET_B(net548),
    .D(net3496),
    .Q(\i_tinyqv.cpu.instr_data[3][15] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _16883_ (.RESET_B(net547),
    .D(_00485_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _16884_ (.RESET_B(net546),
    .D(_00486_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _16885_ (.RESET_B(net545),
    .D(_00487_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _16886_ (.RESET_B(net960),
    .D(net3312),
    .Q(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_1 _16887_ (.RESET_B(net961),
    .D(_00007_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _16888_ (.RESET_B(net962),
    .D(_00010_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[1] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _16889_ (.RESET_B(net963),
    .D(_00011_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[2] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _16890_ (.RESET_B(net964),
    .D(_00012_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[3] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _16891_ (.RESET_B(net965),
    .D(_00013_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[4] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _16892_ (.RESET_B(net966),
    .D(_00014_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[5] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_1 _16893_ (.RESET_B(net967),
    .D(_00015_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[6] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16894_ (.RESET_B(net968),
    .D(_00016_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[7] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16895_ (.RESET_B(net969),
    .D(_00017_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[8] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16896_ (.RESET_B(net970),
    .D(_00018_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[9] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16897_ (.RESET_B(net1147),
    .D(_00008_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[10] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_1 _16898_ (.RESET_B(net544),
    .D(_00009_),
    .Q(\i_tinyqv.cpu.i_core.multiplier.accum[11] ),
    .CLK(clknet_leaf_176_clk_regs));
 sg13g2_dfrbpq_2 _16899_ (.RESET_B(net543),
    .D(net3580),
    .Q(\i_tinyqv.cpu.i_core.mepc[0] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16900_ (.RESET_B(net510),
    .D(net3766),
    .Q(\i_tinyqv.cpu.i_core.mepc[1] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16901_ (.RESET_B(net509),
    .D(net3326),
    .Q(\i_tinyqv.cpu.i_core.mepc[2] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _16902_ (.RESET_B(net508),
    .D(_00492_),
    .Q(\i_tinyqv.cpu.i_core.mepc[3] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16903_ (.RESET_B(net507),
    .D(_00493_),
    .Q(\i_tinyqv.cpu.i_core.mepc[4] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _16904_ (.RESET_B(net506),
    .D(net3566),
    .Q(\i_tinyqv.cpu.i_core.mepc[5] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _16905_ (.RESET_B(net505),
    .D(_00495_),
    .Q(\i_tinyqv.cpu.i_core.mepc[6] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _16906_ (.RESET_B(net504),
    .D(net3358),
    .Q(\i_tinyqv.cpu.i_core.mepc[7] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_1 _16907_ (.RESET_B(net502),
    .D(net3388),
    .Q(\i_tinyqv.cpu.i_core.mepc[8] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16908_ (.RESET_B(net501),
    .D(net3276),
    .Q(\i_tinyqv.cpu.i_core.mepc[9] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16909_ (.RESET_B(net500),
    .D(net3345),
    .Q(\i_tinyqv.cpu.i_core.mepc[10] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _16910_ (.RESET_B(net499),
    .D(_00500_),
    .Q(\i_tinyqv.cpu.i_core.mepc[11] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_1 _16911_ (.RESET_B(net498),
    .D(net3340),
    .Q(\i_tinyqv.cpu.i_core.mepc[12] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _16912_ (.RESET_B(net497),
    .D(_00502_),
    .Q(\i_tinyqv.cpu.i_core.mepc[13] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16913_ (.RESET_B(net496),
    .D(_00503_),
    .Q(\i_tinyqv.cpu.i_core.mepc[14] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _16914_ (.RESET_B(net495),
    .D(_00504_),
    .Q(\i_tinyqv.cpu.i_core.mepc[15] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _16915_ (.RESET_B(net494),
    .D(_00505_),
    .Q(\i_tinyqv.cpu.i_core.mepc[16] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_1 _16916_ (.RESET_B(net493),
    .D(_00506_),
    .Q(\i_tinyqv.cpu.i_core.mepc[17] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_1 _16917_ (.RESET_B(net492),
    .D(_00507_),
    .Q(\i_tinyqv.cpu.i_core.mepc[18] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_1 _16918_ (.RESET_B(net491),
    .D(_00508_),
    .Q(\i_tinyqv.cpu.i_core.mepc[19] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_1 _16919_ (.RESET_B(net490),
    .D(net3541),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_1 _16920_ (.RESET_B(net488),
    .D(net4105),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _16921_ (.RESET_B(net487),
    .D(net3994),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .CLK(clknet_leaf_175_clk_regs));
 sg13g2_dfrbpq_2 _16922_ (.RESET_B(net486),
    .D(net3720),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[3] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_2 _16923_ (.RESET_B(net485),
    .D(_00513_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_2 _16924_ (.RESET_B(net484),
    .D(_00514_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_1 _16925_ (.RESET_B(net483),
    .D(_00515_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16926_ (.RESET_B(net482),
    .D(_00516_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .CLK(clknet_leaf_177_clk_regs));
 sg13g2_dfrbpq_2 _16927_ (.RESET_B(net68),
    .D(_00517_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16928_ (.RESET_B(net67),
    .D(_00518_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16929_ (.RESET_B(net66),
    .D(_00519_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _16930_ (.RESET_B(net65),
    .D(_00520_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16931_ (.RESET_B(net64),
    .D(net3539),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16932_ (.RESET_B(net63),
    .D(net3687),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .CLK(clknet_leaf_1_clk_regs));
 sg13g2_dfrbpq_2 _16933_ (.RESET_B(net34),
    .D(net3616),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16934_ (.RESET_B(net33),
    .D(net3639),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16935_ (.RESET_B(net32),
    .D(net3722),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16936_ (.RESET_B(net31),
    .D(net3833),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16937_ (.RESET_B(net30),
    .D(net3849),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16938_ (.RESET_B(net1421),
    .D(net3787),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16939_ (.RESET_B(net1420),
    .D(_00529_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16940_ (.RESET_B(net1419),
    .D(net3930),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _16941_ (.RESET_B(net1418),
    .D(net3951),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .CLK(clknet_leaf_4_clk_regs));
 sg13g2_dfrbpq_2 _16942_ (.RESET_B(net1417),
    .D(net3942),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16943_ (.RESET_B(net1416),
    .D(net3399),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .CLK(clknet_leaf_0_clk_regs));
 sg13g2_dfrbpq_2 _16944_ (.RESET_B(net1415),
    .D(_00534_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16945_ (.RESET_B(net1414),
    .D(net4019),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .CLK(clknet_leaf_7_clk_regs));
 sg13g2_dfrbpq_2 _16946_ (.RESET_B(net1413),
    .D(net3981),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .CLK(clknet_leaf_3_clk_regs));
 sg13g2_dfrbpq_2 _16947_ (.RESET_B(net1412),
    .D(net3000),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[30] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _16948_ (.RESET_B(net1411),
    .D(_00538_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _16949_ (.RESET_B(net1410),
    .D(net2871),
    .Q(\i_tinyqv.cpu.instr_data[1][0] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _16950_ (.RESET_B(net1408),
    .D(net2908),
    .Q(\i_tinyqv.cpu.instr_data[1][1] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _16951_ (.RESET_B(net1406),
    .D(net3103),
    .Q(\i_peripherals.func_sel[42] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _16952_ (.RESET_B(net1404),
    .D(net3552),
    .Q(\i_peripherals.func_sel[43] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _16953_ (.RESET_B(net1402),
    .D(net3777),
    .Q(\i_peripherals.func_sel[44] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _16954_ (.RESET_B(net1400),
    .D(net3379),
    .Q(\i_peripherals.func_sel[45] ),
    .CLK(clknet_leaf_42_clk_regs));
 sg13g2_dfrbpq_1 _16955_ (.RESET_B(net1398),
    .D(net3724),
    .Q(\i_peripherals.func_sel[46] ),
    .CLK(clknet_leaf_41_clk_regs));
 sg13g2_dfrbpq_1 _16956_ (.RESET_B(net1396),
    .D(_00546_),
    .Q(\i_peripherals.func_sel[47] ),
    .CLK(clknet_leaf_43_clk_regs));
 sg13g2_dfrbpq_1 _16957_ (.RESET_B(net1394),
    .D(_00547_),
    .Q(\i_peripherals.func_sel[36] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16958_ (.RESET_B(net1392),
    .D(net2758),
    .Q(\i_peripherals.func_sel[37] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16959_ (.RESET_B(net1390),
    .D(_00549_),
    .Q(\i_peripherals.func_sel[38] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16960_ (.RESET_B(net1388),
    .D(net3349),
    .Q(\i_peripherals.func_sel[39] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16961_ (.RESET_B(net1386),
    .D(net2825),
    .Q(\i_peripherals.func_sel[40] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _16962_ (.RESET_B(net1384),
    .D(_00552_),
    .Q(\i_peripherals.func_sel[41] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16963_ (.RESET_B(net1382),
    .D(_00553_),
    .Q(\i_peripherals.func_sel[30] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16964_ (.RESET_B(net1380),
    .D(net2778),
    .Q(\i_peripherals.func_sel[31] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16965_ (.RESET_B(net1378),
    .D(_00555_),
    .Q(\i_peripherals.func_sel[32] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16966_ (.RESET_B(net1376),
    .D(net2791),
    .Q(\i_peripherals.func_sel[33] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16967_ (.RESET_B(net1374),
    .D(net2889),
    .Q(\i_peripherals.func_sel[34] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16968_ (.RESET_B(net1372),
    .D(net2766),
    .Q(\i_peripherals.func_sel[35] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16969_ (.RESET_B(net1370),
    .D(_00559_),
    .Q(\i_peripherals.func_sel[24] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16970_ (.RESET_B(net1368),
    .D(net2749),
    .Q(\i_peripherals.func_sel[25] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16971_ (.RESET_B(net1366),
    .D(net2816),
    .Q(\i_peripherals.func_sel[26] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16972_ (.RESET_B(net1364),
    .D(_00562_),
    .Q(\i_peripherals.func_sel[27] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16973_ (.RESET_B(net1362),
    .D(net3025),
    .Q(\i_peripherals.func_sel[28] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16974_ (.RESET_B(net1360),
    .D(net2768),
    .Q(\i_peripherals.func_sel[29] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16975_ (.RESET_B(net1358),
    .D(_00565_),
    .Q(\i_peripherals.func_sel[18] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _16976_ (.RESET_B(net1356),
    .D(net2760),
    .Q(\i_peripherals.func_sel[19] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _16977_ (.RESET_B(net1354),
    .D(_00567_),
    .Q(\i_peripherals.func_sel[20] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16978_ (.RESET_B(net1352),
    .D(net2762),
    .Q(\i_peripherals.func_sel[21] ),
    .CLK(clknet_leaf_34_clk_regs));
 sg13g2_dfrbpq_1 _16979_ (.RESET_B(net1350),
    .D(net2804),
    .Q(\i_peripherals.func_sel[22] ),
    .CLK(clknet_leaf_32_clk_regs));
 sg13g2_dfrbpq_1 _16980_ (.RESET_B(net1348),
    .D(net2756),
    .Q(\i_peripherals.func_sel[23] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _16981_ (.RESET_B(net1346),
    .D(net3618),
    .Q(\i_peripherals.func_sel[12] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16982_ (.RESET_B(net1344),
    .D(net2754),
    .Q(\i_peripherals.func_sel[13] ),
    .CLK(clknet_leaf_37_clk_regs));
 sg13g2_dfrbpq_1 _16983_ (.RESET_B(net1342),
    .D(_00573_),
    .Q(\i_peripherals.func_sel[14] ),
    .CLK(clknet_leaf_35_clk_regs));
 sg13g2_dfrbpq_1 _16984_ (.RESET_B(net1340),
    .D(_00574_),
    .Q(\i_peripherals.func_sel[15] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16985_ (.RESET_B(net1338),
    .D(net2891),
    .Q(\i_peripherals.func_sel[16] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16986_ (.RESET_B(net1336),
    .D(net2764),
    .Q(\i_peripherals.func_sel[17] ),
    .CLK(clknet_leaf_36_clk_regs));
 sg13g2_dfrbpq_1 _16987_ (.RESET_B(net1334),
    .D(net3075),
    .Q(\i_peripherals.func_sel[6] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _16988_ (.RESET_B(net1332),
    .D(net3278),
    .Q(\i_peripherals.func_sel[7] ),
    .CLK(clknet_leaf_39_clk_regs));
 sg13g2_dfrbpq_1 _16989_ (.RESET_B(net1330),
    .D(_00579_),
    .Q(\i_peripherals.func_sel[8] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _16990_ (.RESET_B(net1327),
    .D(net2797),
    .Q(\i_peripherals.func_sel[9] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_1 _16991_ (.RESET_B(net1325),
    .D(net2921),
    .Q(\i_peripherals.func_sel[10] ),
    .CLK(clknet_leaf_40_clk_regs));
 sg13g2_dfrbpq_1 _16992_ (.RESET_B(net1323),
    .D(net2784),
    .Q(\i_peripherals.func_sel[11] ),
    .CLK(clknet_leaf_38_clk_regs));
 sg13g2_dfrbpq_2 _16993_ (.RESET_B(net1321),
    .D(net3691),
    .Q(\i_peripherals.i_uart.baud_divider[8] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16994_ (.RESET_B(net1319),
    .D(net3925),
    .Q(\i_peripherals.i_uart.baud_divider[9] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _16995_ (.RESET_B(net1317),
    .D(net3728),
    .Q(\i_peripherals.i_uart.baud_divider[10] ),
    .CLK(clknet_leaf_51_clk_regs));
 sg13g2_dfrbpq_2 _16996_ (.RESET_B(net1315),
    .D(net3893),
    .Q(\i_peripherals.i_uart.baud_divider[11] ),
    .CLK(clknet_leaf_74_clk_regs));
 sg13g2_dfrbpq_2 _16997_ (.RESET_B(net1313),
    .D(net3785),
    .Q(\i_peripherals.i_uart.baud_divider[12] ),
    .CLK(clknet_leaf_52_clk_regs));
 sg13g2_dfrbpq_2 _16998_ (.RESET_B(net1311),
    .D(_00588_),
    .Q(\i_peripherals.i_user_peri39.busy_counter[2] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _16999_ (.RESET_B(net1309),
    .D(_00589_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[22] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_2 _17000_ (.RESET_B(net1308),
    .D(_00590_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[23] ),
    .CLK(clknet_leaf_87_clk_regs));
 sg13g2_dfrbpq_1 _17001_ (.RESET_B(net1307),
    .D(_00591_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[24] ),
    .CLK(clknet_leaf_85_clk_regs));
 sg13g2_dfrbpq_2 _17002_ (.RESET_B(net1306),
    .D(_00592_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[25] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _17003_ (.RESET_B(net1305),
    .D(_00593_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[26] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _17004_ (.RESET_B(net1304),
    .D(net3706),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[27] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _17005_ (.RESET_B(net1303),
    .D(_00595_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[28] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _17006_ (.RESET_B(net1302),
    .D(_00596_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[29] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _17007_ (.RESET_B(net1301),
    .D(_00597_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[30] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_2 _17008_ (.RESET_B(net1300),
    .D(_00598_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[31] ),
    .CLK(clknet_leaf_88_clk_regs));
 sg13g2_dfrbpq_1 _17009_ (.RESET_B(net1299),
    .D(_00599_),
    .Q(\i_peripherals.i_user_peri39.stage1_math_rec[32] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _17010_ (.RESET_B(net1298),
    .D(_00600_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _17011_ (.RESET_B(net1297),
    .D(_00601_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17012_ (.RESET_B(net1296),
    .D(_00602_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _17013_ (.RESET_B(net1295),
    .D(_00603_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_2 _17014_ (.RESET_B(net1294),
    .D(_00604_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _17015_ (.RESET_B(net1293),
    .D(_00605_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _17016_ (.RESET_B(net1292),
    .D(_00606_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _17017_ (.RESET_B(net1291),
    .D(_00607_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _17018_ (.RESET_B(net1290),
    .D(_00608_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _17019_ (.RESET_B(net1289),
    .D(_00609_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _17020_ (.RESET_B(net1288),
    .D(_00610_),
    .Q(\i_tinyqv.cpu.imm[12] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _17021_ (.RESET_B(net1287),
    .D(_00611_),
    .Q(\i_tinyqv.cpu.imm[13] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_2 _17022_ (.RESET_B(net1286),
    .D(_00612_),
    .Q(\i_tinyqv.cpu.imm[14] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _17023_ (.RESET_B(net1285),
    .D(_00613_),
    .Q(\i_tinyqv.cpu.imm[15] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17024_ (.RESET_B(net1284),
    .D(_00614_),
    .Q(\i_tinyqv.cpu.imm[16] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _17025_ (.RESET_B(net1283),
    .D(_00615_),
    .Q(\i_tinyqv.cpu.imm[17] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17026_ (.RESET_B(net1282),
    .D(_00616_),
    .Q(\i_tinyqv.cpu.imm[18] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_2 _17027_ (.RESET_B(net1281),
    .D(_00617_),
    .Q(\i_tinyqv.cpu.imm[19] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _17028_ (.RESET_B(net1280),
    .D(_00618_),
    .Q(\i_tinyqv.cpu.imm[20] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _17029_ (.RESET_B(net1279),
    .D(_00619_),
    .Q(\i_tinyqv.cpu.imm[21] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _17030_ (.RESET_B(net1278),
    .D(_00620_),
    .Q(\i_tinyqv.cpu.imm[22] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_2 _17031_ (.RESET_B(net1277),
    .D(_00621_),
    .Q(\i_tinyqv.cpu.imm[23] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _17032_ (.RESET_B(net1276),
    .D(_00622_),
    .Q(\i_tinyqv.cpu.imm[24] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _17033_ (.RESET_B(net1275),
    .D(_00623_),
    .Q(\i_tinyqv.cpu.imm[25] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_1 _17034_ (.RESET_B(net1274),
    .D(_00624_),
    .Q(\i_tinyqv.cpu.imm[26] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _17035_ (.RESET_B(net1273),
    .D(_00625_),
    .Q(\i_tinyqv.cpu.imm[27] ),
    .CLK(clknet_leaf_13_clk_regs));
 sg13g2_dfrbpq_1 _17036_ (.RESET_B(net1272),
    .D(_00626_),
    .Q(\i_tinyqv.cpu.imm[28] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _17037_ (.RESET_B(net1271),
    .D(_00627_),
    .Q(\i_tinyqv.cpu.imm[29] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_1 _17038_ (.RESET_B(net1270),
    .D(_00628_),
    .Q(\i_tinyqv.cpu.imm[30] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_1 _17039_ (.RESET_B(net1269),
    .D(_00629_),
    .Q(\i_tinyqv.cpu.imm[31] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _17040_ (.RESET_B(net1268),
    .D(_00630_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _17041_ (.RESET_B(net1266),
    .D(_00631_),
    .Q(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _17042_ (.RESET_B(net1264),
    .D(_00632_),
    .Q(\i_tinyqv.cpu.instr_write_offset[1] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _17043_ (.RESET_B(net1263),
    .D(_00633_),
    .Q(\i_tinyqv.cpu.instr_write_offset[2] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _17044_ (.RESET_B(net1262),
    .D(_00634_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17045_ (.RESET_B(net1261),
    .D(net3165),
    .Q(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _17046_ (.RESET_B(net1260),
    .D(net3562),
    .Q(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _17047_ (.RESET_B(net1259),
    .D(net3175),
    .Q(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_1 _17048_ (.RESET_B(net1258),
    .D(net3600),
    .Q(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17049_ (.RESET_B(net1257),
    .D(net3209),
    .Q(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17050_ (.RESET_B(net1229),
    .D(_00640_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17051_ (.RESET_B(net1227),
    .D(net3657),
    .Q(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17052_ (.RESET_B(net1224),
    .D(_00642_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17053_ (.RESET_B(net1222),
    .D(net2810),
    .Q(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17054_ (.RESET_B(net1220),
    .D(net3524),
    .Q(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _17055_ (.RESET_B(net1218),
    .D(_00645_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _17056_ (.RESET_B(net1216),
    .D(net3537),
    .Q(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_1 _17057_ (.RESET_B(net1214),
    .D(net2917),
    .Q(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_1 _17058_ (.RESET_B(net1212),
    .D(_00648_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _17059_ (.RESET_B(net1210),
    .D(net3544),
    .Q(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_1 _17060_ (.RESET_B(net1208),
    .D(_00650_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17061_ (.RESET_B(net1207),
    .D(_00651_),
    .Q(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17062_ (.RESET_B(net1206),
    .D(net3304),
    .Q(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17063_ (.RESET_B(net1204),
    .D(net3320),
    .Q(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_1 _17064_ (.RESET_B(net1202),
    .D(net2930),
    .Q(\i_tinyqv.cpu.instr_data[0][0] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17065_ (.RESET_B(net1198),
    .D(net2944),
    .Q(\i_tinyqv.cpu.instr_data[0][1] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _17066_ (.RESET_B(net1192),
    .D(net3224),
    .Q(\i_tinyqv.cpu.instr_data[2][0] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _17067_ (.RESET_B(net1172),
    .D(net3114),
    .Q(\i_tinyqv.cpu.instr_data[2][1] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_1 _17068_ (.RESET_B(net1168),
    .D(_00658_),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[28] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _17069_ (.RESET_B(net1166),
    .D(_00659_),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[29] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17070_ (.RESET_B(net1164),
    .D(_00660_),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[30] ),
    .CLK(clknet_leaf_96_clk_regs));
 sg13g2_dfrbpq_1 _17071_ (.RESET_B(net1162),
    .D(_00661_),
    .Q(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[31] ),
    .CLK(clknet_leaf_161_clk_regs));
 sg13g2_dfrbpq_2 _17072_ (.RESET_B(net1160),
    .D(net2959),
    .Q(\i_tinyqv.mem.data_stall ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _17073_ (.RESET_B(net1156),
    .D(net3947),
    .Q(\i_tinyqv.mem.data_txn_len[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _17074_ (.RESET_B(net1329),
    .D(net3884),
    .Q(\i_tinyqv.mem.data_txn_len[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _17075_ (.RESET_B(net1152),
    .D(net3424),
    .Q(\i_tinyqv.mem.qspi_write_done ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _17076_ (.RESET_B(net1148),
    .D(net3647),
    .Q(\i_tinyqv.mem.continue_txn ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _17077_ (.RESET_B(net1145),
    .D(net4029),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _17078_ (.RESET_B(net1141),
    .D(_00667_),
    .Q(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _17079_ (.RESET_B(net1137),
    .D(net3246),
    .Q(\i_tinyqv.cpu.instr_data_in[0] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _17080_ (.RESET_B(net1135),
    .D(net3555),
    .Q(\i_tinyqv.cpu.instr_data_in[1] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17081_ (.RESET_B(net1133),
    .D(net3845),
    .Q(\i_tinyqv.cpu.instr_data_in[2] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _17082_ (.RESET_B(net1131),
    .D(net3637),
    .Q(\i_tinyqv.cpu.instr_data_in[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_2 _17083_ (.RESET_B(net1129),
    .D(net3046),
    .Q(\i_tinyqv.cpu.instr_data_in[4] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17084_ (.RESET_B(net1127),
    .D(net4087),
    .Q(\i_tinyqv.cpu.instr_data_in[5] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17085_ (.RESET_B(net1125),
    .D(net4056),
    .Q(\i_tinyqv.cpu.instr_data_in[6] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17086_ (.RESET_B(net1123),
    .D(net3933),
    .Q(\i_tinyqv.cpu.instr_data_in[7] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17087_ (.RESET_B(net1121),
    .D(net2950),
    .Q(\i_tinyqv.mem.qspi_data_buf[8] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17088_ (.RESET_B(net1119),
    .D(net3019),
    .Q(\i_tinyqv.mem.qspi_data_buf[9] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _17089_ (.RESET_B(net1117),
    .D(net2932),
    .Q(\i_tinyqv.mem.qspi_data_buf[10] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17090_ (.RESET_B(net1115),
    .D(net2788),
    .Q(\i_tinyqv.mem.qspi_data_buf[11] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17091_ (.RESET_B(net1113),
    .D(net2883),
    .Q(\i_tinyqv.mem.qspi_data_buf[12] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17092_ (.RESET_B(net1111),
    .D(net3088),
    .Q(\i_tinyqv.mem.qspi_data_buf[13] ),
    .CLK(clknet_leaf_56_clk_regs));
 sg13g2_dfrbpq_1 _17093_ (.RESET_B(net1109),
    .D(net3630),
    .Q(\i_tinyqv.mem.qspi_data_buf[14] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _17094_ (.RESET_B(net1107),
    .D(_00683_),
    .Q(\i_tinyqv.mem.qspi_data_buf[15] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17095_ (.RESET_B(net1105),
    .D(net2852),
    .Q(\i_tinyqv.mem.data_from_read[16] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _17096_ (.RESET_B(net1103),
    .D(net2840),
    .Q(\i_tinyqv.mem.data_from_read[17] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17097_ (.RESET_B(net1101),
    .D(net2868),
    .Q(\i_tinyqv.mem.data_from_read[18] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17098_ (.RESET_B(net1099),
    .D(net2833),
    .Q(\i_tinyqv.mem.data_from_read[19] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _17099_ (.RESET_B(net1097),
    .D(net3010),
    .Q(\i_tinyqv.mem.data_from_read[20] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17100_ (.RESET_B(net1095),
    .D(net3614),
    .Q(\i_tinyqv.mem.data_from_read[21] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_1 _17101_ (.RESET_B(net1093),
    .D(net3594),
    .Q(\i_tinyqv.mem.data_from_read[22] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _17102_ (.RESET_B(net1091),
    .D(net3494),
    .Q(\i_tinyqv.mem.data_from_read[23] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _17103_ (.RESET_B(net1089),
    .D(net3343),
    .Q(\i_tinyqv.mem.qspi_data_buf[24] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17104_ (.RESET_B(net1087),
    .D(net3434),
    .Q(\i_tinyqv.mem.qspi_data_buf[25] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_2 _17105_ (.RESET_B(net1085),
    .D(_00694_),
    .Q(\i_tinyqv.mem.qspi_data_buf[26] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17106_ (.RESET_B(net1083),
    .D(net3455),
    .Q(\i_tinyqv.mem.qspi_data_buf[27] ),
    .CLK(clknet_leaf_66_clk_regs));
 sg13g2_dfrbpq_2 _17107_ (.RESET_B(net1081),
    .D(net3322),
    .Q(\i_tinyqv.mem.qspi_data_buf[28] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17108_ (.RESET_B(net1079),
    .D(net3612),
    .Q(\i_tinyqv.mem.qspi_data_buf[29] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17109_ (.RESET_B(net1077),
    .D(net3660),
    .Q(\i_tinyqv.mem.qspi_data_buf[30] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_1 _17110_ (.RESET_B(net1075),
    .D(_00699_),
    .Q(\i_tinyqv.mem.qspi_data_buf[31] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_1 _17111_ (.RESET_B(net1073),
    .D(_00700_),
    .Q(\i_tinyqv.cpu.instr_fetch_started ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _17112_ (.RESET_B(net1071),
    .D(net4116),
    .Q(\i_tinyqv.mem.instr_active ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _17113_ (.RESET_B(net1067),
    .D(_00702_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _17114_ (.RESET_B(net1065),
    .D(_00703_),
    .Q(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _17115_ (.RESET_B(net1063),
    .D(net4072),
    .Q(\i_tinyqv.mem.q_ctrl.data_req ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _17116_ (.RESET_B(net1061),
    .D(net3793),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _17117_ (.RESET_B(net1057),
    .D(net3709),
    .Q(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _17118_ (.RESET_B(net1053),
    .D(net3754),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .CLK(clknet_leaf_30_clk_regs));
 sg13g2_dfrbpq_2 _17119_ (.RESET_B(net1049),
    .D(net3483),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _17120_ (.RESET_B(net1045),
    .D(net3815),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _17121_ (.RESET_B(net1041),
    .D(net3240),
    .Q(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _17122_ (.RESET_B(net1037),
    .D(_00711_),
    .Q(\i_tinyqv.mem.q_ctrl.is_writing ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_2 _17123_ (.RESET_B(net1033),
    .D(net3968),
    .Q(\i_tinyqv.mem.q_ctrl.data_ready ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_2 _17124_ (.RESET_B(net1031),
    .D(_00713_),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _17125_ (.RESET_B(net1027),
    .D(net3280),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _17126_ (.RESET_B(net1023),
    .D(net4094),
    .Q(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_1 _17127_ (.RESET_B(net1019),
    .D(_00716_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17128_ (.RESET_B(net1015),
    .D(_00717_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17129_ (.RESET_B(net1011),
    .D(_00718_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .CLK(clknet_leaf_29_clk_regs));
 sg13g2_dfrbpq_1 _17130_ (.RESET_B(net1007),
    .D(net3510),
    .Q(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .CLK(clknet_leaf_33_clk_regs));
 sg13g2_dfrbpq_2 _17131_ (.RESET_B(net1003),
    .D(_00720_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .CLK(clknet_leaf_173_clk_regs));
 sg13g2_dfrbpq_2 _17132_ (.RESET_B(net895),
    .D(_00721_),
    .Q(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _17133_ (.RESET_B(net889),
    .D(net3156),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _17134_ (.RESET_B(net887),
    .D(net3132),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _17135_ (.RESET_B(net885),
    .D(net3139),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_1 _17136_ (.RESET_B(net883),
    .D(net3171),
    .Q(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _17137_ (.RESET_B(net881),
    .D(_00726_),
    .Q(\i_tinyqv.cpu.instr_data_in[8] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _17138_ (.RESET_B(net879),
    .D(net3992),
    .Q(\i_tinyqv.cpu.instr_data_in[9] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _17139_ (.RESET_B(net877),
    .D(_00728_),
    .Q(\i_tinyqv.cpu.instr_data_in[10] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _17140_ (.RESET_B(net875),
    .D(net3955),
    .Q(\i_tinyqv.cpu.instr_data_in[11] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_1 _17141_ (.RESET_B(net873),
    .D(_00730_),
    .Q(\i_tinyqv.cpu.instr_data_in[12] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _17142_ (.RESET_B(net871),
    .D(_00731_),
    .Q(\i_tinyqv.cpu.instr_data_in[13] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _17143_ (.RESET_B(net869),
    .D(net3997),
    .Q(\i_tinyqv.cpu.instr_data_in[14] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_2 _17144_ (.RESET_B(net865),
    .D(_00733_),
    .Q(\i_tinyqv.cpu.instr_data_in[15] ),
    .CLK(clknet_leaf_58_clk_regs));
 sg13g2_dfrbpq_1 _17145_ (.RESET_B(net863),
    .D(_00734_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17146_ (.RESET_B(net861),
    .D(_00735_),
    .Q(\i_tinyqv.mem.q_ctrl.last_ram_a_sel ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_1 _17147_ (.RESET_B(net859),
    .D(_00736_),
    .Q(\i_tinyqv.cpu.instr_fetch_stopped ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _17148_ (.RESET_B(net857),
    .D(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_neg ),
    .CLK(net1435));
 sg13g2_dfrbpq_1 _17149_ (.RESET_B(net855),
    .D(_00737_),
    .Q(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ),
    .CLK(clknet_leaf_31_clk_regs));
 sg13g2_dfrbpq_1 _17150_ (.RESET_B(net853),
    .D(net3453),
    .Q(\i_tinyqv.cpu.instr_data[2][2] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17151_ (.RESET_B(net851),
    .D(net3441),
    .Q(\i_tinyqv.cpu.instr_data[2][3] ),
    .CLK(clknet_leaf_14_clk_regs));
 sg13g2_dfrbpq_1 _17152_ (.RESET_B(net849),
    .D(_00740_),
    .Q(\i_tinyqv.cpu.instr_data[2][4] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _17153_ (.RESET_B(net847),
    .D(net3522),
    .Q(\i_tinyqv.cpu.instr_data[2][5] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_1 _17154_ (.RESET_B(net845),
    .D(net3422),
    .Q(\i_tinyqv.cpu.instr_data[2][6] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _17155_ (.RESET_B(net843),
    .D(net3116),
    .Q(\i_tinyqv.cpu.instr_data[2][7] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _17156_ (.RESET_B(net841),
    .D(net3439),
    .Q(\i_tinyqv.cpu.instr_data[2][8] ),
    .CLK(clknet_leaf_154_clk_regs));
 sg13g2_dfrbpq_1 _17157_ (.RESET_B(net839),
    .D(net3211),
    .Q(\i_tinyqv.cpu.instr_data[2][9] ),
    .CLK(clknet_leaf_152_clk_regs));
 sg13g2_dfrbpq_1 _17158_ (.RESET_B(net837),
    .D(net3231),
    .Q(\i_tinyqv.cpu.instr_data[2][10] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_1 _17159_ (.RESET_B(net835),
    .D(net3080),
    .Q(\i_tinyqv.cpu.instr_data[2][11] ),
    .CLK(clknet_leaf_153_clk_regs));
 sg13g2_dfrbpq_1 _17160_ (.RESET_B(net833),
    .D(net3429),
    .Q(\i_tinyqv.cpu.instr_data[2][12] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _17161_ (.RESET_B(net831),
    .D(net3107),
    .Q(\i_tinyqv.cpu.instr_data[2][13] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_1 _17162_ (.RESET_B(net829),
    .D(net3078),
    .Q(\i_tinyqv.cpu.instr_data[2][14] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _17163_ (.RESET_B(net827),
    .D(net3712),
    .Q(\i_tinyqv.cpu.instr_data[2][15] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _17164_ (.RESET_B(net825),
    .D(net3008),
    .Q(\i_tinyqv.cpu.i_core.load_top_bit ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _17165_ (.RESET_B(net821),
    .D(_00753_),
    .Q(\i_tinyqv.cpu.pc[1] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17166_ (.RESET_B(net817),
    .D(_00754_),
    .Q(\i_tinyqv.cpu.pc[2] ),
    .CLK(clknet_leaf_12_clk_regs));
 sg13g2_dfrbpq_2 _17167_ (.RESET_B(net805),
    .D(net3112),
    .Q(\i_peripherals.i_user_peri39._GEN[64] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17168_ (.RESET_B(net802),
    .D(net2986),
    .Q(\i_peripherals.i_user_peri39._GEN[65] ),
    .CLK(clknet_leaf_80_clk_regs));
 sg13g2_dfrbpq_2 _17169_ (.RESET_B(net800),
    .D(net3181),
    .Q(\i_peripherals.i_user_peri39._GEN[66] ),
    .CLK(clknet_leaf_79_clk_regs));
 sg13g2_dfrbpq_2 _17170_ (.RESET_B(net798),
    .D(net3263),
    .Q(\i_peripherals.i_user_peri39._GEN[67] ),
    .CLK(clknet_leaf_84_clk_regs));
 sg13g2_dfrbpq_2 _17171_ (.RESET_B(net796),
    .D(net3159),
    .Q(\i_peripherals.i_user_peri39._GEN[68] ),
    .CLK(clknet_leaf_76_clk_regs));
 sg13g2_dfrbpq_2 _17172_ (.RESET_B(net773),
    .D(_00760_),
    .Q(\i_peripherals.i_user_peri39._GEN[69] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_2 _17173_ (.RESET_B(net771),
    .D(net3101),
    .Q(\i_peripherals.i_user_peri39._GEN[70] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17174_ (.RESET_B(net769),
    .D(net3242),
    .Q(\i_peripherals.i_user_peri39._GEN[71] ),
    .CLK(clknet_leaf_78_clk_regs));
 sg13g2_dfrbpq_2 _17175_ (.RESET_B(net767),
    .D(net3531),
    .Q(\i_peripherals.i_user_peri39._GEN[72] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17176_ (.RESET_B(net765),
    .D(net3583),
    .Q(\i_peripherals.i_user_peri39._GEN[73] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _17177_ (.RESET_B(net763),
    .D(net3673),
    .Q(\i_peripherals.i_user_peri39._GEN[74] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17178_ (.RESET_B(net761),
    .D(net3501),
    .Q(\i_peripherals.i_user_peri39._GEN[75] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_2 _17179_ (.RESET_B(net759),
    .D(net3489),
    .Q(\i_peripherals.i_user_peri39._GEN[76] ),
    .CLK(clknet_leaf_81_clk_regs));
 sg13g2_dfrbpq_2 _17180_ (.RESET_B(net757),
    .D(net3021),
    .Q(\i_peripherals.i_user_peri39._GEN[77] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_1 _17181_ (.RESET_B(net755),
    .D(net2936),
    .Q(\i_peripherals.i_user_peri39._GEN[78] ),
    .CLK(clknet_leaf_90_clk_regs));
 sg13g2_dfrbpq_1 _17182_ (.RESET_B(net753),
    .D(net2879),
    .Q(\i_peripherals.i_user_peri39._GEN[79] ),
    .CLK(clknet_leaf_67_clk_regs));
 sg13g2_dfrbpq_2 _17183_ (.RESET_B(net751),
    .D(net2903),
    .Q(\i_peripherals.i_user_peri39._GEN[80] ),
    .CLK(clknet_leaf_91_clk_regs));
 sg13g2_dfrbpq_2 _17184_ (.RESET_B(net749),
    .D(net2848),
    .Q(\i_peripherals.i_user_peri39._GEN[81] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_2 _17185_ (.RESET_B(net747),
    .D(net2954),
    .Q(\i_peripherals.i_user_peri39._GEN[82] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_2 _17186_ (.RESET_B(net745),
    .D(net2881),
    .Q(\i_peripherals.i_user_peri39._GEN[83] ),
    .CLK(clknet_leaf_92_clk_regs));
 sg13g2_dfrbpq_2 _17187_ (.RESET_B(net743),
    .D(net3515),
    .Q(\i_peripherals.i_user_peri39._GEN[84] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17188_ (.RESET_B(net741),
    .D(net2842),
    .Q(\i_peripherals.i_user_peri39._GEN[85] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_2 _17189_ (.RESET_B(net739),
    .D(net2914),
    .Q(\i_peripherals.i_user_peri39._GEN[86] ),
    .CLK(clknet_leaf_93_clk_regs));
 sg13g2_dfrbpq_1 _17190_ (.RESET_B(net737),
    .D(net3050),
    .Q(\i_peripherals.i_user_peri39._GEN[87] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_2 _17191_ (.RESET_B(net735),
    .D(net2877),
    .Q(\i_peripherals.i_user_peri39._GEN[88] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_1 _17192_ (.RESET_B(net733),
    .D(net2808),
    .Q(\i_peripherals.i_user_peri39._GEN[89] ),
    .CLK(clknet_leaf_70_clk_regs));
 sg13g2_dfrbpq_2 _17193_ (.RESET_B(net731),
    .D(net2827),
    .Q(\i_peripherals.i_user_peri39._GEN[90] ),
    .CLK(clknet_leaf_68_clk_regs));
 sg13g2_dfrbpq_1 _17194_ (.RESET_B(net729),
    .D(net2812),
    .Q(\i_peripherals.i_user_peri39._GEN[91] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_1 _17195_ (.RESET_B(net727),
    .D(net2875),
    .Q(\i_peripherals.i_user_peri39._GEN[92] ),
    .CLK(clknet_leaf_71_clk_regs));
 sg13g2_dfrbpq_1 _17196_ (.RESET_B(net725),
    .D(net2820),
    .Q(\i_peripherals.i_user_peri39._GEN[93] ),
    .CLK(clknet_leaf_82_clk_regs));
 sg13g2_dfrbpq_1 _17197_ (.RESET_B(net723),
    .D(net3135),
    .Q(\i_peripherals.i_user_peri39._GEN[94] ),
    .CLK(clknet_leaf_89_clk_regs));
 sg13g2_dfrbpq_1 _17198_ (.RESET_B(net721),
    .D(net3006),
    .Q(\i_peripherals.i_user_peri39._GEN[95] ),
    .CLK(clknet_leaf_69_clk_regs));
 sg13g2_dfrbpq_2 _17199_ (.RESET_B(net719),
    .D(_00787_),
    .Q(\i_tinyqv.cpu.instr_data_start[3] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17200_ (.RESET_B(net715),
    .D(_00788_),
    .Q(\i_tinyqv.cpu.instr_data_start[4] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _17201_ (.RESET_B(net711),
    .D(_00789_),
    .Q(\i_tinyqv.cpu.instr_data_start[5] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _17202_ (.RESET_B(net707),
    .D(_00790_),
    .Q(\i_tinyqv.cpu.instr_data_start[6] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _17203_ (.RESET_B(net703),
    .D(_00791_),
    .Q(\i_tinyqv.cpu.instr_data_start[7] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _17204_ (.RESET_B(net699),
    .D(_00792_),
    .Q(\i_tinyqv.cpu.instr_data_start[8] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _17205_ (.RESET_B(net695),
    .D(_00793_),
    .Q(\i_tinyqv.cpu.instr_data_start[9] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _17206_ (.RESET_B(net691),
    .D(_00794_),
    .Q(\i_tinyqv.cpu.instr_data_start[10] ),
    .CLK(clknet_leaf_2_clk_regs));
 sg13g2_dfrbpq_2 _17207_ (.RESET_B(net687),
    .D(_00795_),
    .Q(\i_tinyqv.cpu.instr_data_start[11] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _17208_ (.RESET_B(net683),
    .D(_00796_),
    .Q(\i_tinyqv.cpu.instr_data_start[12] ),
    .CLK(clknet_leaf_6_clk_regs));
 sg13g2_dfrbpq_2 _17209_ (.RESET_B(net678),
    .D(_00797_),
    .Q(\i_tinyqv.cpu.instr_data_start[13] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_1 _17210_ (.RESET_B(net674),
    .D(_00798_),
    .Q(\i_tinyqv.cpu.instr_data_start[14] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _17211_ (.RESET_B(net670),
    .D(_00799_),
    .Q(\i_tinyqv.cpu.instr_data_start[15] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _17212_ (.RESET_B(net666),
    .D(_00800_),
    .Q(\i_tinyqv.cpu.instr_data_start[16] ),
    .CLK(clknet_leaf_5_clk_regs));
 sg13g2_dfrbpq_2 _17213_ (.RESET_B(net662),
    .D(_00801_),
    .Q(\i_tinyqv.cpu.instr_data_start[17] ),
    .CLK(clknet_leaf_8_clk_regs));
 sg13g2_dfrbpq_2 _17214_ (.RESET_B(net658),
    .D(_00802_),
    .Q(\i_tinyqv.cpu.instr_data_start[18] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _17215_ (.RESET_B(net654),
    .D(_00803_),
    .Q(\i_tinyqv.cpu.instr_data_start[19] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _17216_ (.RESET_B(net650),
    .D(_00804_),
    .Q(\i_tinyqv.cpu.instr_data_start[20] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _17217_ (.RESET_B(net646),
    .D(_00805_),
    .Q(\i_tinyqv.cpu.instr_data_start[21] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _17218_ (.RESET_B(net642),
    .D(_00806_),
    .Q(\i_tinyqv.cpu.instr_data_start[22] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _17219_ (.RESET_B(net638),
    .D(_00807_),
    .Q(\i_tinyqv.cpu.instr_data_start[23] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _17220_ (.RESET_B(net634),
    .D(_00808_),
    .Q(\i_tinyqv.cpu.instr_fetch_running ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _17221_ (.RESET_B(net630),
    .D(_00809_),
    .Q(\i_tinyqv.cpu.was_early_branch ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _17222_ (.RESET_B(net626),
    .D(_00810_),
    .Q(\data_to_write[0] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _17223_ (.RESET_B(net622),
    .D(_00811_),
    .Q(\data_to_write[1] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _17224_ (.RESET_B(net618),
    .D(_00812_),
    .Q(\data_to_write[2] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_1 _17225_ (.RESET_B(net614),
    .D(_00813_),
    .Q(\data_to_write[3] ),
    .CLK(clknet_leaf_15_clk_regs));
 sg13g2_dfrbpq_1 _17226_ (.RESET_B(net610),
    .D(_00814_),
    .Q(\data_to_write[4] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_1 _17227_ (.RESET_B(net1409),
    .D(_00815_),
    .Q(\data_to_write[5] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _17228_ (.RESET_B(net1405),
    .D(_00816_),
    .Q(\data_to_write[6] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _17229_ (.RESET_B(net1401),
    .D(_00817_),
    .Q(\data_to_write[7] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _17230_ (.RESET_B(net1397),
    .D(_00818_),
    .Q(\data_to_write[8] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17231_ (.RESET_B(net1393),
    .D(_00819_),
    .Q(\data_to_write[9] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17232_ (.RESET_B(net1389),
    .D(_00820_),
    .Q(\data_to_write[10] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _17233_ (.RESET_B(net1385),
    .D(_00821_),
    .Q(\data_to_write[11] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17234_ (.RESET_B(net1381),
    .D(_00822_),
    .Q(\data_to_write[12] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17235_ (.RESET_B(net1377),
    .D(_00823_),
    .Q(\data_to_write[13] ),
    .CLK(clknet_leaf_62_clk_regs));
 sg13g2_dfrbpq_2 _17236_ (.RESET_B(net1373),
    .D(_00824_),
    .Q(\data_to_write[14] ),
    .CLK(clknet_leaf_61_clk_regs));
 sg13g2_dfrbpq_2 _17237_ (.RESET_B(net1369),
    .D(_00825_),
    .Q(\data_to_write[15] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17238_ (.RESET_B(net1365),
    .D(_00826_),
    .Q(\data_to_write[16] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _17239_ (.RESET_B(net1361),
    .D(_00827_),
    .Q(\data_to_write[17] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _17240_ (.RESET_B(net1357),
    .D(_00828_),
    .Q(\data_to_write[18] ),
    .CLK(clknet_leaf_94_clk_regs));
 sg13g2_dfrbpq_2 _17241_ (.RESET_B(net1353),
    .D(_00829_),
    .Q(\data_to_write[19] ),
    .CLK(clknet_leaf_63_clk_regs));
 sg13g2_dfrbpq_2 _17242_ (.RESET_B(net1349),
    .D(_00830_),
    .Q(\data_to_write[20] ),
    .CLK(clknet_leaf_53_clk_regs));
 sg13g2_dfrbpq_2 _17243_ (.RESET_B(net1345),
    .D(_00831_),
    .Q(\data_to_write[21] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17244_ (.RESET_B(net1341),
    .D(_00832_),
    .Q(\data_to_write[22] ),
    .CLK(clknet_leaf_55_clk_regs));
 sg13g2_dfrbpq_2 _17245_ (.RESET_B(net1337),
    .D(_00833_),
    .Q(\data_to_write[23] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17246_ (.RESET_B(net1333),
    .D(_00834_),
    .Q(\data_to_write[24] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17247_ (.RESET_B(net1328),
    .D(_00835_),
    .Q(\data_to_write[25] ),
    .CLK(clknet_leaf_59_clk_regs));
 sg13g2_dfrbpq_2 _17248_ (.RESET_B(net1324),
    .D(_00836_),
    .Q(\data_to_write[26] ),
    .CLK(clknet_leaf_54_clk_regs));
 sg13g2_dfrbpq_2 _17249_ (.RESET_B(net1320),
    .D(_00837_),
    .Q(\data_to_write[27] ),
    .CLK(clknet_leaf_72_clk_regs));
 sg13g2_dfrbpq_2 _17250_ (.RESET_B(net1316),
    .D(_00838_),
    .Q(\data_to_write[28] ),
    .CLK(clknet_leaf_64_clk_regs));
 sg13g2_dfrbpq_2 _17251_ (.RESET_B(net1312),
    .D(_00839_),
    .Q(\data_to_write[29] ),
    .CLK(clknet_leaf_65_clk_regs));
 sg13g2_dfrbpq_2 _17252_ (.RESET_B(net1267),
    .D(_00840_),
    .Q(\data_to_write[30] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17253_ (.RESET_B(net1200),
    .D(_00841_),
    .Q(\data_to_write[31] ),
    .CLK(clknet_leaf_60_clk_regs));
 sg13g2_dfrbpq_2 _17254_ (.RESET_B(net1186),
    .D(net4052),
    .Q(\i_tinyqv.cpu.data_write_n[0] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _17255_ (.RESET_B(net1158),
    .D(net4050),
    .Q(\i_tinyqv.cpu.data_write_n[1] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _17256_ (.RESET_B(net1150),
    .D(net3799),
    .Q(\i_tinyqv.cpu.data_read_n[0] ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _17257_ (.RESET_B(net644),
    .D(net3801),
    .Q(\i_tinyqv.cpu.data_read_n[1] ),
    .CLK(clknet_leaf_18_clk_regs));
 sg13g2_dfrbpq_2 _17258_ (.RESET_B(net1139),
    .D(net4004),
    .Q(debug_data_continue),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _17259_ (.RESET_B(net1059),
    .D(_00846_),
    .Q(\i_tinyqv.cpu.no_write_in_progress ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_1 _17260_ (.RESET_B(net1051),
    .D(net2776),
    .Q(\i_tinyqv.cpu.load_started ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _17261_ (.RESET_B(net1043),
    .D(net3853),
    .Q(\addr[0] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_1 _17262_ (.RESET_B(net1035),
    .D(_00849_),
    .Q(\addr[1] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _17263_ (.RESET_B(net1025),
    .D(_00850_),
    .Q(\addr[2] ),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17264_ (.RESET_B(net1017),
    .D(_00851_),
    .Q(\addr[3] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _17265_ (.RESET_B(net1009),
    .D(_00852_),
    .Q(\addr[4] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_2 _17266_ (.RESET_B(net1001),
    .D(net4062),
    .Q(\addr[5] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _17267_ (.RESET_B(net823),
    .D(net3667),
    .Q(\addr[6] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_2 _17268_ (.RESET_B(net815),
    .D(net3828),
    .Q(\addr[7] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_2 _17269_ (.RESET_B(net713),
    .D(_00856_),
    .Q(\addr[8] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _17270_ (.RESET_B(net705),
    .D(_00857_),
    .Q(\addr[9] ),
    .CLK(clknet_leaf_20_clk_regs));
 sg13g2_dfrbpq_2 _17271_ (.RESET_B(net697),
    .D(net3377),
    .Q(\addr[10] ),
    .CLK(clknet_leaf_22_clk_regs));
 sg13g2_dfrbpq_2 _17272_ (.RESET_B(net689),
    .D(_00859_),
    .Q(\addr[11] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _17273_ (.RESET_B(net681),
    .D(net2992),
    .Q(\addr[12] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _17274_ (.RESET_B(net672),
    .D(net3177),
    .Q(\addr[13] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _17275_ (.RESET_B(net664),
    .D(net3173),
    .Q(\addr[14] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _17276_ (.RESET_B(net656),
    .D(net3238),
    .Q(\addr[15] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _17277_ (.RESET_B(net648),
    .D(net3096),
    .Q(\addr[16] ),
    .CLK(clknet_leaf_25_clk_regs));
 sg13g2_dfrbpq_2 _17278_ (.RESET_B(net640),
    .D(net3220),
    .Q(\addr[17] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _17279_ (.RESET_B(net632),
    .D(net3169),
    .Q(\addr[18] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _17280_ (.RESET_B(net624),
    .D(net3198),
    .Q(\addr[19] ),
    .CLK(clknet_leaf_26_clk_regs));
 sg13g2_dfrbpq_2 _17281_ (.RESET_B(net616),
    .D(_00868_),
    .Q(\addr[20] ),
    .CLK(clknet_leaf_27_clk_regs));
 sg13g2_dfrbpq_2 _17282_ (.RESET_B(net608),
    .D(_00869_),
    .Q(\addr[21] ),
    .CLK(clknet_leaf_28_clk_regs));
 sg13g2_dfrbpq_2 _17283_ (.RESET_B(net1403),
    .D(net3044),
    .Q(\addr[22] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _17284_ (.RESET_B(net1395),
    .D(net3445),
    .Q(\addr[23] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _17285_ (.RESET_B(net1387),
    .D(_00872_),
    .Q(\addr[24] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_2 _17286_ (.RESET_B(net1379),
    .D(_00873_),
    .Q(\addr[25] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _17287_ (.RESET_B(net1371),
    .D(_00874_),
    .Q(\addr[26] ),
    .CLK(clknet_leaf_23_clk_regs));
 sg13g2_dfrbpq_2 _17288_ (.RESET_B(net1363),
    .D(_00875_),
    .Q(\addr[27] ),
    .CLK(clknet_leaf_24_clk_regs));
 sg13g2_dfrbpq_1 _17289_ (.RESET_B(net1355),
    .D(_00876_),
    .Q(\i_tinyqv.cpu.counter[2] ),
    .CLK(clknet_leaf_19_clk_regs));
 sg13g2_dfrbpq_1 _17290_ (.RESET_B(net1351),
    .D(_00877_),
    .Q(\i_tinyqv.cpu.counter[3] ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_1 _17291_ (.RESET_B(net1347),
    .D(_00878_),
    .Q(\i_tinyqv.cpu.counter[4] ),
    .CLK(clknet_leaf_16_clk_regs));
 sg13g2_dfrbpq_1 _17292_ (.RESET_B(net1343),
    .D(_00879_),
    .Q(\i_tinyqv.cpu.data_ready_sync ),
    .CLK(clknet_leaf_17_clk_regs));
 sg13g2_dfrbpq_2 _17293_ (.RESET_B(net1335),
    .D(_00880_),
    .Q(\i_tinyqv.cpu.is_load ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _17294_ (.RESET_B(net1326),
    .D(_00881_),
    .Q(\i_tinyqv.cpu.is_alu_imm ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _17295_ (.RESET_B(net1318),
    .D(_00882_),
    .Q(\i_tinyqv.cpu.is_auipc ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _17296_ (.RESET_B(net1310),
    .D(_00883_),
    .Q(\i_tinyqv.cpu.is_store ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_2 _17297_ (.RESET_B(net1194),
    .D(_00884_),
    .Q(\i_tinyqv.cpu.is_alu_reg ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_2 _17298_ (.RESET_B(net1154),
    .D(_00885_),
    .Q(\i_tinyqv.cpu.is_lui ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _17299_ (.RESET_B(net1069),
    .D(_00886_),
    .Q(\i_tinyqv.cpu.is_branch ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _17300_ (.RESET_B(net1047),
    .D(_00887_),
    .Q(\i_tinyqv.cpu.is_jalr ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _17301_ (.RESET_B(net1029),
    .D(_00888_),
    .Q(\i_tinyqv.cpu.is_jal ),
    .CLK(clknet_leaf_157_clk_regs));
 sg13g2_dfrbpq_2 _17302_ (.RESET_B(net1013),
    .D(_00889_),
    .Q(\i_tinyqv.cpu.is_system ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_2 _17303_ (.RESET_B(net893),
    .D(_00890_),
    .Q(\i_tinyqv.cpu.instr_len[1] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_2 _17304_ (.RESET_B(net717),
    .D(_00891_),
    .Q(\i_tinyqv.cpu.instr_len[2] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_2 _17305_ (.RESET_B(net701),
    .D(_00892_),
    .Q(\i_tinyqv.cpu.alu_op[0] ),
    .CLK(clknet_leaf_158_clk_regs));
 sg13g2_dfrbpq_1 _17306_ (.RESET_B(net685),
    .D(_00893_),
    .Q(\i_tinyqv.cpu.alu_op[1] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_1 _17307_ (.RESET_B(net668),
    .D(_00894_),
    .Q(\i_tinyqv.cpu.alu_op[2] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_2 _17308_ (.RESET_B(net652),
    .D(_00895_),
    .Q(\i_tinyqv.cpu.alu_op[3] ),
    .CLK(clknet_leaf_172_clk_regs));
 sg13g2_dfrbpq_1 _17309_ (.RESET_B(net636),
    .D(_00896_),
    .Q(\i_tinyqv.cpu.data_ready_latch ),
    .CLK(clknet_leaf_21_clk_regs));
 sg13g2_dfrbpq_2 _17310_ (.RESET_B(net628),
    .D(_00897_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .CLK(clknet_leaf_156_clk_regs));
 sg13g2_dfrbpq_2 _17311_ (.RESET_B(net620),
    .D(_00898_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .CLK(clknet_leaf_155_clk_regs));
 sg13g2_dfrbpq_2 _17312_ (.RESET_B(net612),
    .D(_00899_),
    .Q(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .CLK(clknet_leaf_159_clk_regs));
 sg13g2_dfrbpq_2 _17313_ (.RESET_B(net1407),
    .D(_00900_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _17314_ (.RESET_B(net1399),
    .D(_00901_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_2 _17315_ (.RESET_B(net1391),
    .D(_00902_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .CLK(clknet_leaf_147_clk_regs));
 sg13g2_dfrbpq_2 _17316_ (.RESET_B(net1383),
    .D(_00903_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .CLK(clknet_leaf_148_clk_regs));
 sg13g2_dfrbpq_2 _17317_ (.RESET_B(net1375),
    .D(_00904_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .CLK(clknet_leaf_146_clk_regs));
 sg13g2_dfrbpq_2 _17318_ (.RESET_B(net1367),
    .D(_00905_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _17319_ (.RESET_B(net1359),
    .D(_00906_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_2 _17320_ (.RESET_B(net1339),
    .D(_00907_),
    .Q(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .CLK(clknet_leaf_145_clk_regs));
 sg13g2_dfrbpq_2 _17321_ (.RESET_B(net1331),
    .D(_00908_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_2 _17322_ (.RESET_B(net1314),
    .D(net3840),
    .Q(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_1 _17323_ (.RESET_B(net1170),
    .D(_00910_),
    .Q(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .CLK(clknet_leaf_151_clk_regs));
 sg13g2_dfrbpq_2 _17324_ (.RESET_B(net1055),
    .D(_00911_),
    .Q(\i_tinyqv.cpu.addr_offset[2] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_1 _17325_ (.RESET_B(net1021),
    .D(net2802),
    .Q(\i_tinyqv.cpu.addr_offset[3] ),
    .CLK(clknet_leaf_9_clk_regs));
 sg13g2_dfrbpq_2 _17326_ (.RESET_B(net819),
    .D(_00913_),
    .Q(\i_tinyqv.cpu.mem_op_increment_reg ),
    .CLK(clknet_leaf_150_clk_regs));
 sg13g2_dfrbpq_2 _17327_ (.RESET_B(net693),
    .D(_00914_),
    .Q(\i_tinyqv.cpu.i_core.is_interrupt ),
    .CLK(clknet_leaf_10_clk_regs));
 sg13g2_dfrbpq_2 _17328_ (.RESET_B(net660),
    .D(_00915_),
    .Q(debug_instr_valid),
    .CLK(clknet_leaf_11_clk_regs));
 sg13g2_dfrbpq_2 _17329_ (.RESET_B(net1322),
    .D(_00916_),
    .Q(\time_count[0] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17330_ (.RESET_B(net1265),
    .D(_00917_),
    .Q(\time_count[1] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17331_ (.RESET_B(net1143),
    .D(_00918_),
    .Q(\time_count[2] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17332_ (.RESET_B(net1039),
    .D(net4022),
    .Q(\time_count[3] ),
    .CLK(clknet_leaf_46_clk_regs));
 sg13g2_dfrbpq_1 _17333_ (.RESET_B(net1005),
    .D(_00920_),
    .Q(\time_count[4] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_dfrbpq_2 _17334_ (.RESET_B(net709),
    .D(_00921_),
    .Q(\time_count[5] ),
    .CLK(clknet_leaf_45_clk_regs));
 sg13g2_dfrbpq_1 _17335_ (.RESET_B(net676),
    .D(_00922_),
    .Q(\time_count[6] ),
    .CLK(clknet_leaf_57_clk_regs));
 sg13g2_tiehi _15941__15 (.L_HI(net15));
 sg13g2_tiehi _15942__16 (.L_HI(net16));
 sg13g2_tiehi _15943__17 (.L_HI(net17));
 sg13g2_tiehi _15944__18 (.L_HI(net18));
 sg13g2_tiehi _15945__19 (.L_HI(net19));
 sg13g2_tiehi _15946__20 (.L_HI(net20));
 sg13g2_tiehi _15947__21 (.L_HI(net21));
 sg13g2_tiehi _15948__22 (.L_HI(net22));
 sg13g2_tiehi _15949__23 (.L_HI(net23));
 sg13g2_tiehi _15950__24 (.L_HI(net24));
 sg13g2_tiehi _15951__25 (.L_HI(net25));
 sg13g2_tiehi _15952__26 (.L_HI(net26));
 sg13g2_tiehi _15953__27 (.L_HI(net27));
 sg13g2_tiehi _15954__28 (.L_HI(net28));
 sg13g2_tiehi _15955__29 (.L_HI(net29));
 sg13g2_tiehi _16937__30 (.L_HI(net30));
 sg13g2_tiehi _16936__31 (.L_HI(net31));
 sg13g2_tiehi _16935__32 (.L_HI(net32));
 sg13g2_tiehi _16934__33 (.L_HI(net33));
 sg13g2_tiehi _16933__34 (.L_HI(net34));
 sg13g2_tiehi _15956__35 (.L_HI(net35));
 sg13g2_tiehi _15962__36 (.L_HI(net36));
 sg13g2_tiehi _15963__37 (.L_HI(net37));
 sg13g2_tiehi _15964__38 (.L_HI(net38));
 sg13g2_tiehi _15965__39 (.L_HI(net39));
 sg13g2_tiehi _15966__40 (.L_HI(net40));
 sg13g2_tiehi _15967__41 (.L_HI(net41));
 sg13g2_tiehi _15968__42 (.L_HI(net42));
 sg13g2_tiehi _15969__43 (.L_HI(net43));
 sg13g2_tiehi _15970__44 (.L_HI(net44));
 sg13g2_tiehi _15971__45 (.L_HI(net45));
 sg13g2_tiehi _15972__46 (.L_HI(net46));
 sg13g2_tiehi _15973__47 (.L_HI(net47));
 sg13g2_tiehi _15974__48 (.L_HI(net48));
 sg13g2_tiehi _15975__49 (.L_HI(net49));
 sg13g2_tiehi _15976__50 (.L_HI(net50));
 sg13g2_tiehi _15977__51 (.L_HI(net51));
 sg13g2_tiehi _15978__52 (.L_HI(net52));
 sg13g2_tiehi _15979__53 (.L_HI(net53));
 sg13g2_tiehi _15980__54 (.L_HI(net54));
 sg13g2_tiehi _15981__55 (.L_HI(net55));
 sg13g2_tiehi _15982__56 (.L_HI(net56));
 sg13g2_tiehi _15983__57 (.L_HI(net57));
 sg13g2_tiehi _15984__58 (.L_HI(net58));
 sg13g2_tiehi _15985__59 (.L_HI(net59));
 sg13g2_tiehi _15986__60 (.L_HI(net60));
 sg13g2_tiehi _15987__61 (.L_HI(net61));
 sg13g2_tiehi _15988__62 (.L_HI(net62));
 sg13g2_tiehi _16932__63 (.L_HI(net63));
 sg13g2_tiehi _16931__64 (.L_HI(net64));
 sg13g2_tiehi _16930__65 (.L_HI(net65));
 sg13g2_tiehi _16929__66 (.L_HI(net66));
 sg13g2_tiehi _16928__67 (.L_HI(net67));
 sg13g2_tiehi _16927__68 (.L_HI(net68));
 sg13g2_tiehi _15989__69 (.L_HI(net69));
 sg13g2_tiehi _15996__70 (.L_HI(net70));
 sg13g2_tiehi _15997__71 (.L_HI(net71));
 sg13g2_tiehi _15998__72 (.L_HI(net72));
 sg13g2_tiehi _15999__73 (.L_HI(net73));
 sg13g2_tiehi _16000__74 (.L_HI(net74));
 sg13g2_tiehi _16001__75 (.L_HI(net75));
 sg13g2_tiehi _16002__76 (.L_HI(net76));
 sg13g2_tiehi _16003__77 (.L_HI(net77));
 sg13g2_tiehi _16004__78 (.L_HI(net78));
 sg13g2_tiehi _16005__79 (.L_HI(net79));
 sg13g2_tiehi _16006__80 (.L_HI(net80));
 sg13g2_tiehi _16007__81 (.L_HI(net81));
 sg13g2_tiehi _16008__82 (.L_HI(net82));
 sg13g2_tiehi _16009__83 (.L_HI(net83));
 sg13g2_tiehi _16010__84 (.L_HI(net84));
 sg13g2_tiehi _16011__85 (.L_HI(net85));
 sg13g2_tiehi _16012__86 (.L_HI(net86));
 sg13g2_tiehi _16013__87 (.L_HI(net87));
 sg13g2_tiehi _16014__88 (.L_HI(net88));
 sg13g2_tiehi _16015__89 (.L_HI(net89));
 sg13g2_tiehi _16016__90 (.L_HI(net90));
 sg13g2_tiehi _16017__91 (.L_HI(net91));
 sg13g2_tiehi _16018__92 (.L_HI(net92));
 sg13g2_tiehi _16019__93 (.L_HI(net93));
 sg13g2_tiehi _16020__94 (.L_HI(net94));
 sg13g2_tiehi _16021__95 (.L_HI(net95));
 sg13g2_tiehi _16022__96 (.L_HI(net96));
 sg13g2_tiehi _16023__97 (.L_HI(net97));
 sg13g2_tiehi _16024__98 (.L_HI(net98));
 sg13g2_tiehi _16025__99 (.L_HI(net99));
 sg13g2_tiehi _16026__100 (.L_HI(net100));
 sg13g2_tiehi _16027__101 (.L_HI(net101));
 sg13g2_tiehi _16028__102 (.L_HI(net102));
 sg13g2_tiehi _16029__103 (.L_HI(net103));
 sg13g2_tiehi _16030__104 (.L_HI(net104));
 sg13g2_tiehi _16031__105 (.L_HI(net105));
 sg13g2_tiehi _16032__106 (.L_HI(net106));
 sg13g2_tiehi _16033__107 (.L_HI(net107));
 sg13g2_tiehi _16034__108 (.L_HI(net108));
 sg13g2_tiehi _16035__109 (.L_HI(net109));
 sg13g2_tiehi _16036__110 (.L_HI(net110));
 sg13g2_tiehi _16037__111 (.L_HI(net111));
 sg13g2_tiehi _16038__112 (.L_HI(net112));
 sg13g2_tiehi _16039__113 (.L_HI(net113));
 sg13g2_tiehi _16040__114 (.L_HI(net114));
 sg13g2_tiehi _16041__115 (.L_HI(net115));
 sg13g2_tiehi _16042__116 (.L_HI(net116));
 sg13g2_tiehi _16043__117 (.L_HI(net117));
 sg13g2_tiehi _16044__118 (.L_HI(net118));
 sg13g2_tiehi _16045__119 (.L_HI(net119));
 sg13g2_tiehi _16046__120 (.L_HI(net120));
 sg13g2_tiehi _16047__121 (.L_HI(net121));
 sg13g2_tiehi _16048__122 (.L_HI(net122));
 sg13g2_tiehi _16049__123 (.L_HI(net123));
 sg13g2_tiehi _16050__124 (.L_HI(net124));
 sg13g2_tiehi _16051__125 (.L_HI(net125));
 sg13g2_tiehi _16052__126 (.L_HI(net126));
 sg13g2_tiehi _16053__127 (.L_HI(net127));
 sg13g2_tiehi _16054__128 (.L_HI(net128));
 sg13g2_tiehi _16055__129 (.L_HI(net129));
 sg13g2_tiehi _16056__130 (.L_HI(net130));
 sg13g2_tiehi _16057__131 (.L_HI(net131));
 sg13g2_tiehi _16058__132 (.L_HI(net132));
 sg13g2_tiehi _16059__133 (.L_HI(net133));
 sg13g2_tiehi _16060__134 (.L_HI(net134));
 sg13g2_tiehi _16061__135 (.L_HI(net135));
 sg13g2_tiehi _16062__136 (.L_HI(net136));
 sg13g2_tiehi _16063__137 (.L_HI(net137));
 sg13g2_tiehi _16064__138 (.L_HI(net138));
 sg13g2_tiehi _16065__139 (.L_HI(net139));
 sg13g2_tiehi _16066__140 (.L_HI(net140));
 sg13g2_tiehi _16067__141 (.L_HI(net141));
 sg13g2_tiehi _16068__142 (.L_HI(net142));
 sg13g2_tiehi _16069__143 (.L_HI(net143));
 sg13g2_tiehi _16070__144 (.L_HI(net144));
 sg13g2_tiehi _16071__145 (.L_HI(net145));
 sg13g2_tiehi _16072__146 (.L_HI(net146));
 sg13g2_tiehi _16073__147 (.L_HI(net147));
 sg13g2_tiehi _16074__148 (.L_HI(net148));
 sg13g2_tiehi _16075__149 (.L_HI(net149));
 sg13g2_tiehi _16076__150 (.L_HI(net150));
 sg13g2_tiehi _16077__151 (.L_HI(net151));
 sg13g2_tiehi _16078__152 (.L_HI(net152));
 sg13g2_tiehi _16079__153 (.L_HI(net153));
 sg13g2_tiehi _16080__154 (.L_HI(net154));
 sg13g2_tiehi _16081__155 (.L_HI(net155));
 sg13g2_tiehi _16082__156 (.L_HI(net156));
 sg13g2_tiehi _16083__157 (.L_HI(net157));
 sg13g2_tiehi _16084__158 (.L_HI(net158));
 sg13g2_tiehi _16085__159 (.L_HI(net159));
 sg13g2_tiehi _16086__160 (.L_HI(net160));
 sg13g2_tiehi _16087__161 (.L_HI(net161));
 sg13g2_tiehi _16088__162 (.L_HI(net162));
 sg13g2_tiehi _16089__163 (.L_HI(net163));
 sg13g2_tiehi _16090__164 (.L_HI(net164));
 sg13g2_tiehi _16091__165 (.L_HI(net165));
 sg13g2_tiehi _16092__166 (.L_HI(net166));
 sg13g2_tiehi _16093__167 (.L_HI(net167));
 sg13g2_tiehi _16094__168 (.L_HI(net168));
 sg13g2_tiehi _16095__169 (.L_HI(net169));
 sg13g2_tiehi _16096__170 (.L_HI(net170));
 sg13g2_tiehi _16097__171 (.L_HI(net171));
 sg13g2_tiehi _16098__172 (.L_HI(net172));
 sg13g2_tiehi _16099__173 (.L_HI(net173));
 sg13g2_tiehi _16100__174 (.L_HI(net174));
 sg13g2_tiehi _16101__175 (.L_HI(net175));
 sg13g2_tiehi _16102__176 (.L_HI(net176));
 sg13g2_tiehi _16103__177 (.L_HI(net177));
 sg13g2_tiehi _16104__178 (.L_HI(net178));
 sg13g2_tiehi _16105__179 (.L_HI(net179));
 sg13g2_tiehi _16106__180 (.L_HI(net180));
 sg13g2_tiehi _16107__181 (.L_HI(net181));
 sg13g2_tiehi _16108__182 (.L_HI(net182));
 sg13g2_tiehi _16109__183 (.L_HI(net183));
 sg13g2_tiehi _16110__184 (.L_HI(net184));
 sg13g2_tiehi _16111__185 (.L_HI(net185));
 sg13g2_tiehi _16112__186 (.L_HI(net186));
 sg13g2_tiehi _16113__187 (.L_HI(net187));
 sg13g2_tiehi _16114__188 (.L_HI(net188));
 sg13g2_tiehi _16115__189 (.L_HI(net189));
 sg13g2_tiehi _16116__190 (.L_HI(net190));
 sg13g2_tiehi _16117__191 (.L_HI(net191));
 sg13g2_tiehi _16118__192 (.L_HI(net192));
 sg13g2_tiehi _16119__193 (.L_HI(net193));
 sg13g2_tiehi _16120__194 (.L_HI(net194));
 sg13g2_tiehi _16121__195 (.L_HI(net195));
 sg13g2_tiehi _16122__196 (.L_HI(net196));
 sg13g2_tiehi _16123__197 (.L_HI(net197));
 sg13g2_tiehi _16124__198 (.L_HI(net198));
 sg13g2_tiehi _16125__199 (.L_HI(net199));
 sg13g2_tiehi _16126__200 (.L_HI(net200));
 sg13g2_tiehi _16127__201 (.L_HI(net201));
 sg13g2_tiehi _16128__202 (.L_HI(net202));
 sg13g2_tiehi _16129__203 (.L_HI(net203));
 sg13g2_tiehi _16130__204 (.L_HI(net204));
 sg13g2_tiehi _16131__205 (.L_HI(net205));
 sg13g2_tiehi _16132__206 (.L_HI(net206));
 sg13g2_tiehi _16133__207 (.L_HI(net207));
 sg13g2_tiehi _16134__208 (.L_HI(net208));
 sg13g2_tiehi _16135__209 (.L_HI(net209));
 sg13g2_tiehi _16136__210 (.L_HI(net210));
 sg13g2_tiehi _16137__211 (.L_HI(net211));
 sg13g2_tiehi _16138__212 (.L_HI(net212));
 sg13g2_tiehi _16139__213 (.L_HI(net213));
 sg13g2_tiehi _16140__214 (.L_HI(net214));
 sg13g2_tiehi _16141__215 (.L_HI(net215));
 sg13g2_tiehi _16142__216 (.L_HI(net216));
 sg13g2_tiehi _16143__217 (.L_HI(net217));
 sg13g2_tiehi _16144__218 (.L_HI(net218));
 sg13g2_tiehi _16145__219 (.L_HI(net219));
 sg13g2_tiehi _16146__220 (.L_HI(net220));
 sg13g2_tiehi _16147__221 (.L_HI(net221));
 sg13g2_tiehi _16148__222 (.L_HI(net222));
 sg13g2_tiehi _16149__223 (.L_HI(net223));
 sg13g2_tiehi _16150__224 (.L_HI(net224));
 sg13g2_tiehi _16151__225 (.L_HI(net225));
 sg13g2_tiehi _16152__226 (.L_HI(net226));
 sg13g2_tiehi _16153__227 (.L_HI(net227));
 sg13g2_tiehi _16154__228 (.L_HI(net228));
 sg13g2_tiehi _16155__229 (.L_HI(net229));
 sg13g2_tiehi _16156__230 (.L_HI(net230));
 sg13g2_tiehi _16157__231 (.L_HI(net231));
 sg13g2_tiehi _16158__232 (.L_HI(net232));
 sg13g2_tiehi _16159__233 (.L_HI(net233));
 sg13g2_tiehi _16160__234 (.L_HI(net234));
 sg13g2_tiehi _16161__235 (.L_HI(net235));
 sg13g2_tiehi _16162__236 (.L_HI(net236));
 sg13g2_tiehi _16163__237 (.L_HI(net237));
 sg13g2_tiehi _16164__238 (.L_HI(net238));
 sg13g2_tiehi _16165__239 (.L_HI(net239));
 sg13g2_tiehi _16166__240 (.L_HI(net240));
 sg13g2_tiehi _16167__241 (.L_HI(net241));
 sg13g2_tiehi _16168__242 (.L_HI(net242));
 sg13g2_tiehi _16169__243 (.L_HI(net243));
 sg13g2_tiehi _16170__244 (.L_HI(net244));
 sg13g2_tiehi _16171__245 (.L_HI(net245));
 sg13g2_tiehi _16172__246 (.L_HI(net246));
 sg13g2_tiehi _16173__247 (.L_HI(net247));
 sg13g2_tiehi _16174__248 (.L_HI(net248));
 sg13g2_tiehi _16175__249 (.L_HI(net249));
 sg13g2_tiehi _16176__250 (.L_HI(net250));
 sg13g2_tiehi _16177__251 (.L_HI(net251));
 sg13g2_tiehi _16178__252 (.L_HI(net252));
 sg13g2_tiehi _16179__253 (.L_HI(net253));
 sg13g2_tiehi _16180__254 (.L_HI(net254));
 sg13g2_tiehi _16181__255 (.L_HI(net255));
 sg13g2_tiehi _16182__256 (.L_HI(net256));
 sg13g2_tiehi _16183__257 (.L_HI(net257));
 sg13g2_tiehi _16184__258 (.L_HI(net258));
 sg13g2_tiehi _16185__259 (.L_HI(net259));
 sg13g2_tiehi _16186__260 (.L_HI(net260));
 sg13g2_tiehi _16187__261 (.L_HI(net261));
 sg13g2_tiehi _16188__262 (.L_HI(net262));
 sg13g2_tiehi _16189__263 (.L_HI(net263));
 sg13g2_tiehi _16190__264 (.L_HI(net264));
 sg13g2_tiehi _16191__265 (.L_HI(net265));
 sg13g2_tiehi _16192__266 (.L_HI(net266));
 sg13g2_tiehi _16193__267 (.L_HI(net267));
 sg13g2_tiehi _16194__268 (.L_HI(net268));
 sg13g2_tiehi _16195__269 (.L_HI(net269));
 sg13g2_tiehi _16196__270 (.L_HI(net270));
 sg13g2_tiehi _16197__271 (.L_HI(net271));
 sg13g2_tiehi _16198__272 (.L_HI(net272));
 sg13g2_tiehi _16199__273 (.L_HI(net273));
 sg13g2_tiehi _16200__274 (.L_HI(net274));
 sg13g2_tiehi _16201__275 (.L_HI(net275));
 sg13g2_tiehi _16202__276 (.L_HI(net276));
 sg13g2_tiehi _16203__277 (.L_HI(net277));
 sg13g2_tiehi _16204__278 (.L_HI(net278));
 sg13g2_tiehi _16205__279 (.L_HI(net279));
 sg13g2_tiehi _16206__280 (.L_HI(net280));
 sg13g2_tiehi _16207__281 (.L_HI(net281));
 sg13g2_tiehi _16208__282 (.L_HI(net282));
 sg13g2_tiehi _16209__283 (.L_HI(net283));
 sg13g2_tiehi _16210__284 (.L_HI(net284));
 sg13g2_tiehi _16211__285 (.L_HI(net285));
 sg13g2_tiehi _16212__286 (.L_HI(net286));
 sg13g2_tiehi _16213__287 (.L_HI(net287));
 sg13g2_tiehi _16214__288 (.L_HI(net288));
 sg13g2_tiehi _16215__289 (.L_HI(net289));
 sg13g2_tiehi _16216__290 (.L_HI(net290));
 sg13g2_tiehi _16217__291 (.L_HI(net291));
 sg13g2_tiehi _16218__292 (.L_HI(net292));
 sg13g2_tiehi _16219__293 (.L_HI(net293));
 sg13g2_tiehi _16220__294 (.L_HI(net294));
 sg13g2_tiehi _16221__295 (.L_HI(net295));
 sg13g2_tiehi _16222__296 (.L_HI(net296));
 sg13g2_tiehi _16223__297 (.L_HI(net297));
 sg13g2_tiehi _16224__298 (.L_HI(net298));
 sg13g2_tiehi _16225__299 (.L_HI(net299));
 sg13g2_tiehi _16226__300 (.L_HI(net300));
 sg13g2_tiehi _16227__301 (.L_HI(net301));
 sg13g2_tiehi _16228__302 (.L_HI(net302));
 sg13g2_tiehi _16229__303 (.L_HI(net303));
 sg13g2_tiehi _16230__304 (.L_HI(net304));
 sg13g2_tiehi _16231__305 (.L_HI(net305));
 sg13g2_tiehi _16232__306 (.L_HI(net306));
 sg13g2_tiehi _16233__307 (.L_HI(net307));
 sg13g2_tiehi _16234__308 (.L_HI(net308));
 sg13g2_tiehi _16235__309 (.L_HI(net309));
 sg13g2_tiehi _16236__310 (.L_HI(net310));
 sg13g2_tiehi _16237__311 (.L_HI(net311));
 sg13g2_tiehi _16238__312 (.L_HI(net312));
 sg13g2_tiehi _16239__313 (.L_HI(net313));
 sg13g2_tiehi _16240__314 (.L_HI(net314));
 sg13g2_tiehi _16241__315 (.L_HI(net315));
 sg13g2_tiehi _16242__316 (.L_HI(net316));
 sg13g2_tiehi _16243__317 (.L_HI(net317));
 sg13g2_tiehi _16244__318 (.L_HI(net318));
 sg13g2_tiehi _16245__319 (.L_HI(net319));
 sg13g2_tiehi _16246__320 (.L_HI(net320));
 sg13g2_tiehi _16247__321 (.L_HI(net321));
 sg13g2_tiehi _16248__322 (.L_HI(net322));
 sg13g2_tiehi _16249__323 (.L_HI(net323));
 sg13g2_tiehi _16250__324 (.L_HI(net324));
 sg13g2_tiehi _16251__325 (.L_HI(net325));
 sg13g2_tiehi _16252__326 (.L_HI(net326));
 sg13g2_tiehi _16253__327 (.L_HI(net327));
 sg13g2_tiehi _16254__328 (.L_HI(net328));
 sg13g2_tiehi _16255__329 (.L_HI(net329));
 sg13g2_tiehi _16256__330 (.L_HI(net330));
 sg13g2_tiehi _16257__331 (.L_HI(net331));
 sg13g2_tiehi _16258__332 (.L_HI(net332));
 sg13g2_tiehi _16259__333 (.L_HI(net333));
 sg13g2_tiehi _16260__334 (.L_HI(net334));
 sg13g2_tiehi _16261__335 (.L_HI(net335));
 sg13g2_tiehi _16262__336 (.L_HI(net336));
 sg13g2_tiehi _16263__337 (.L_HI(net337));
 sg13g2_tiehi _16264__338 (.L_HI(net338));
 sg13g2_tiehi _16265__339 (.L_HI(net339));
 sg13g2_tiehi _16266__340 (.L_HI(net340));
 sg13g2_tiehi _16267__341 (.L_HI(net341));
 sg13g2_tiehi _16268__342 (.L_HI(net342));
 sg13g2_tiehi _16269__343 (.L_HI(net343));
 sg13g2_tiehi _16270__344 (.L_HI(net344));
 sg13g2_tiehi _16271__345 (.L_HI(net345));
 sg13g2_tiehi _16272__346 (.L_HI(net346));
 sg13g2_tiehi _16273__347 (.L_HI(net347));
 sg13g2_tiehi _16274__348 (.L_HI(net348));
 sg13g2_tiehi _16275__349 (.L_HI(net349));
 sg13g2_tiehi _16276__350 (.L_HI(net350));
 sg13g2_tiehi _16277__351 (.L_HI(net351));
 sg13g2_tiehi _16278__352 (.L_HI(net352));
 sg13g2_tiehi _16279__353 (.L_HI(net353));
 sg13g2_tiehi _16280__354 (.L_HI(net354));
 sg13g2_tiehi _16281__355 (.L_HI(net355));
 sg13g2_tiehi _16282__356 (.L_HI(net356));
 sg13g2_tiehi _16283__357 (.L_HI(net357));
 sg13g2_tiehi _16284__358 (.L_HI(net358));
 sg13g2_tiehi _16285__359 (.L_HI(net359));
 sg13g2_tiehi _16286__360 (.L_HI(net360));
 sg13g2_tiehi _16287__361 (.L_HI(net361));
 sg13g2_tiehi _16288__362 (.L_HI(net362));
 sg13g2_tiehi _16289__363 (.L_HI(net363));
 sg13g2_tiehi _16290__364 (.L_HI(net364));
 sg13g2_tiehi _16291__365 (.L_HI(net365));
 sg13g2_tiehi _16292__366 (.L_HI(net366));
 sg13g2_tiehi _16293__367 (.L_HI(net367));
 sg13g2_tiehi _16294__368 (.L_HI(net368));
 sg13g2_tiehi _16295__369 (.L_HI(net369));
 sg13g2_tiehi _16296__370 (.L_HI(net370));
 sg13g2_tiehi _16297__371 (.L_HI(net371));
 sg13g2_tiehi _16298__372 (.L_HI(net372));
 sg13g2_tiehi _16299__373 (.L_HI(net373));
 sg13g2_tiehi _16300__374 (.L_HI(net374));
 sg13g2_tiehi _16301__375 (.L_HI(net375));
 sg13g2_tiehi _16302__376 (.L_HI(net376));
 sg13g2_tiehi _16303__377 (.L_HI(net377));
 sg13g2_tiehi _16304__378 (.L_HI(net378));
 sg13g2_tiehi _16305__379 (.L_HI(net379));
 sg13g2_tiehi _16306__380 (.L_HI(net380));
 sg13g2_tiehi _16307__381 (.L_HI(net381));
 sg13g2_tiehi _16308__382 (.L_HI(net382));
 sg13g2_tiehi _16309__383 (.L_HI(net383));
 sg13g2_tiehi _16310__384 (.L_HI(net384));
 sg13g2_tiehi _16311__385 (.L_HI(net385));
 sg13g2_tiehi _16312__386 (.L_HI(net386));
 sg13g2_tiehi _16313__387 (.L_HI(net387));
 sg13g2_tiehi _16314__388 (.L_HI(net388));
 sg13g2_tiehi _16315__389 (.L_HI(net389));
 sg13g2_tiehi _16316__390 (.L_HI(net390));
 sg13g2_tiehi _16317__391 (.L_HI(net391));
 sg13g2_tiehi _16318__392 (.L_HI(net392));
 sg13g2_tiehi _16319__393 (.L_HI(net393));
 sg13g2_tiehi _16320__394 (.L_HI(net394));
 sg13g2_tiehi _16321__395 (.L_HI(net395));
 sg13g2_tiehi _16322__396 (.L_HI(net396));
 sg13g2_tiehi _16323__397 (.L_HI(net397));
 sg13g2_tiehi _16324__398 (.L_HI(net398));
 sg13g2_tiehi _16325__399 (.L_HI(net399));
 sg13g2_tiehi _16326__400 (.L_HI(net400));
 sg13g2_tiehi _16327__401 (.L_HI(net401));
 sg13g2_tiehi _16328__402 (.L_HI(net402));
 sg13g2_tiehi _16329__403 (.L_HI(net403));
 sg13g2_tiehi _16330__404 (.L_HI(net404));
 sg13g2_tiehi _16331__405 (.L_HI(net405));
 sg13g2_tiehi _16332__406 (.L_HI(net406));
 sg13g2_tiehi _16333__407 (.L_HI(net407));
 sg13g2_tiehi _16334__408 (.L_HI(net408));
 sg13g2_tiehi _16335__409 (.L_HI(net409));
 sg13g2_tiehi _16336__410 (.L_HI(net410));
 sg13g2_tiehi _16337__411 (.L_HI(net411));
 sg13g2_tiehi _16338__412 (.L_HI(net412));
 sg13g2_tiehi _16339__413 (.L_HI(net413));
 sg13g2_tiehi _16340__414 (.L_HI(net414));
 sg13g2_tiehi _16341__415 (.L_HI(net415));
 sg13g2_tiehi _16342__416 (.L_HI(net416));
 sg13g2_tiehi _16343__417 (.L_HI(net417));
 sg13g2_tiehi _16344__418 (.L_HI(net418));
 sg13g2_tiehi _16345__419 (.L_HI(net419));
 sg13g2_tiehi _16346__420 (.L_HI(net420));
 sg13g2_tiehi _16347__421 (.L_HI(net421));
 sg13g2_tiehi _16348__422 (.L_HI(net422));
 sg13g2_tiehi _16349__423 (.L_HI(net423));
 sg13g2_tiehi _16350__424 (.L_HI(net424));
 sg13g2_tiehi _16351__425 (.L_HI(net425));
 sg13g2_tiehi _16352__426 (.L_HI(net426));
 sg13g2_tiehi _16353__427 (.L_HI(net427));
 sg13g2_tiehi _16354__428 (.L_HI(net428));
 sg13g2_tiehi _16355__429 (.L_HI(net429));
 sg13g2_tiehi _16356__430 (.L_HI(net430));
 sg13g2_tiehi _16357__431 (.L_HI(net431));
 sg13g2_tiehi _16358__432 (.L_HI(net432));
 sg13g2_tiehi _16359__433 (.L_HI(net433));
 sg13g2_tiehi _16360__434 (.L_HI(net434));
 sg13g2_tiehi _16361__435 (.L_HI(net435));
 sg13g2_tiehi _16362__436 (.L_HI(net436));
 sg13g2_tiehi _16363__437 (.L_HI(net437));
 sg13g2_tiehi _16364__438 (.L_HI(net438));
 sg13g2_tiehi _16365__439 (.L_HI(net439));
 sg13g2_tiehi _16366__440 (.L_HI(net440));
 sg13g2_tiehi _16367__441 (.L_HI(net441));
 sg13g2_tiehi _16368__442 (.L_HI(net442));
 sg13g2_tiehi _16369__443 (.L_HI(net443));
 sg13g2_tiehi _16370__444 (.L_HI(net444));
 sg13g2_tiehi _16371__445 (.L_HI(net445));
 sg13g2_tiehi _16372__446 (.L_HI(net446));
 sg13g2_tiehi _16373__447 (.L_HI(net447));
 sg13g2_tiehi _16374__448 (.L_HI(net448));
 sg13g2_tiehi _16375__449 (.L_HI(net449));
 sg13g2_tiehi _16376__450 (.L_HI(net450));
 sg13g2_tiehi _16377__451 (.L_HI(net451));
 sg13g2_tiehi _16378__452 (.L_HI(net452));
 sg13g2_tiehi _16379__453 (.L_HI(net453));
 sg13g2_tiehi _16380__454 (.L_HI(net454));
 sg13g2_tiehi _16381__455 (.L_HI(net455));
 sg13g2_tiehi _16382__456 (.L_HI(net456));
 sg13g2_tiehi _16383__457 (.L_HI(net457));
 sg13g2_tiehi _16384__458 (.L_HI(net458));
 sg13g2_tiehi _16385__459 (.L_HI(net459));
 sg13g2_tiehi _16386__460 (.L_HI(net460));
 sg13g2_tiehi _16387__461 (.L_HI(net461));
 sg13g2_tiehi _16388__462 (.L_HI(net462));
 sg13g2_tiehi _16389__463 (.L_HI(net463));
 sg13g2_tiehi _16390__464 (.L_HI(net464));
 sg13g2_tiehi _16391__465 (.L_HI(net465));
 sg13g2_tiehi _16392__466 (.L_HI(net466));
 sg13g2_tiehi _16393__467 (.L_HI(net467));
 sg13g2_tiehi _16394__468 (.L_HI(net468));
 sg13g2_tiehi _16395__469 (.L_HI(net469));
 sg13g2_tiehi _16396__470 (.L_HI(net470));
 sg13g2_tiehi _16397__471 (.L_HI(net471));
 sg13g2_tiehi _16398__472 (.L_HI(net472));
 sg13g2_tiehi _16399__473 (.L_HI(net473));
 sg13g2_tiehi _16400__474 (.L_HI(net474));
 sg13g2_tiehi _16401__475 (.L_HI(net475));
 sg13g2_tiehi _16402__476 (.L_HI(net476));
 sg13g2_tiehi _16403__477 (.L_HI(net477));
 sg13g2_tiehi _16404__478 (.L_HI(net478));
 sg13g2_tiehi _16405__479 (.L_HI(net479));
 sg13g2_tiehi _16406__480 (.L_HI(net480));
 sg13g2_tiehi _16407__481 (.L_HI(net481));
 sg13g2_tiehi _16926__482 (.L_HI(net482));
 sg13g2_tiehi _16925__483 (.L_HI(net483));
 sg13g2_tiehi _16924__484 (.L_HI(net484));
 sg13g2_tiehi _16923__485 (.L_HI(net485));
 sg13g2_tiehi _16922__486 (.L_HI(net486));
 sg13g2_tiehi _16921__487 (.L_HI(net487));
 sg13g2_tiehi _16920__488 (.L_HI(net488));
 sg13g2_tiehi _16408__489 (.L_HI(net489));
 sg13g2_tiehi _16919__490 (.L_HI(net490));
 sg13g2_tiehi _16918__491 (.L_HI(net491));
 sg13g2_tiehi _16917__492 (.L_HI(net492));
 sg13g2_tiehi _16916__493 (.L_HI(net493));
 sg13g2_tiehi _16915__494 (.L_HI(net494));
 sg13g2_tiehi _16914__495 (.L_HI(net495));
 sg13g2_tiehi _16913__496 (.L_HI(net496));
 sg13g2_tiehi _16912__497 (.L_HI(net497));
 sg13g2_tiehi _16911__498 (.L_HI(net498));
 sg13g2_tiehi _16910__499 (.L_HI(net499));
 sg13g2_tiehi _16909__500 (.L_HI(net500));
 sg13g2_tiehi _16908__501 (.L_HI(net501));
 sg13g2_tiehi _16907__502 (.L_HI(net502));
 sg13g2_tiehi _16416__503 (.L_HI(net503));
 sg13g2_tiehi _16906__504 (.L_HI(net504));
 sg13g2_tiehi _16905__505 (.L_HI(net505));
 sg13g2_tiehi _16904__506 (.L_HI(net506));
 sg13g2_tiehi _16903__507 (.L_HI(net507));
 sg13g2_tiehi _16902__508 (.L_HI(net508));
 sg13g2_tiehi _16901__509 (.L_HI(net509));
 sg13g2_tiehi _16900__510 (.L_HI(net510));
 sg13g2_tiehi _16430__511 (.L_HI(net511));
 sg13g2_tiehi _16438__512 (.L_HI(net512));
 sg13g2_tiehi _16439__513 (.L_HI(net513));
 sg13g2_tiehi _16440__514 (.L_HI(net514));
 sg13g2_tiehi _16441__515 (.L_HI(net515));
 sg13g2_tiehi _16442__516 (.L_HI(net516));
 sg13g2_tiehi _16443__517 (.L_HI(net517));
 sg13g2_tiehi _16444__518 (.L_HI(net518));
 sg13g2_tiehi _16445__519 (.L_HI(net519));
 sg13g2_tiehi _16446__520 (.L_HI(net520));
 sg13g2_tiehi _16447__521 (.L_HI(net521));
 sg13g2_tiehi _16448__522 (.L_HI(net522));
 sg13g2_tiehi _16449__523 (.L_HI(net523));
 sg13g2_tiehi _16450__524 (.L_HI(net524));
 sg13g2_tiehi _16451__525 (.L_HI(net525));
 sg13g2_tiehi _16452__526 (.L_HI(net526));
 sg13g2_tiehi _16453__527 (.L_HI(net527));
 sg13g2_tiehi _16454__528 (.L_HI(net528));
 sg13g2_tiehi _16455__529 (.L_HI(net529));
 sg13g2_tiehi _16456__530 (.L_HI(net530));
 sg13g2_tiehi _16457__531 (.L_HI(net531));
 sg13g2_tiehi _16458__532 (.L_HI(net532));
 sg13g2_tiehi _16459__533 (.L_HI(net533));
 sg13g2_tiehi _16460__534 (.L_HI(net534));
 sg13g2_tiehi _16461__535 (.L_HI(net535));
 sg13g2_tiehi _16462__536 (.L_HI(net536));
 sg13g2_tiehi _16463__537 (.L_HI(net537));
 sg13g2_tiehi _16464__538 (.L_HI(net538));
 sg13g2_tiehi _16465__539 (.L_HI(net539));
 sg13g2_tiehi _16466__540 (.L_HI(net540));
 sg13g2_tiehi _16467__541 (.L_HI(net541));
 sg13g2_tiehi _16468__542 (.L_HI(net542));
 sg13g2_tiehi _16899__543 (.L_HI(net543));
 sg13g2_tiehi _16898__544 (.L_HI(net544));
 sg13g2_tiehi _16885__545 (.L_HI(net545));
 sg13g2_tiehi _16884__546 (.L_HI(net546));
 sg13g2_tiehi _16883__547 (.L_HI(net547));
 sg13g2_tiehi _16882__548 (.L_HI(net548));
 sg13g2_tiehi _16881__549 (.L_HI(net549));
 sg13g2_tiehi _16880__550 (.L_HI(net550));
 sg13g2_tiehi _16879__551 (.L_HI(net551));
 sg13g2_tiehi _16878__552 (.L_HI(net552));
 sg13g2_tiehi _16877__553 (.L_HI(net553));
 sg13g2_tiehi _16876__554 (.L_HI(net554));
 sg13g2_tiehi _16469__555 (.L_HI(net555));
 sg13g2_tiehi _16482__556 (.L_HI(net556));
 sg13g2_tiehi _16483__557 (.L_HI(net557));
 sg13g2_tiehi _16484__558 (.L_HI(net558));
 sg13g2_tiehi _16485__559 (.L_HI(net559));
 sg13g2_tiehi _16486__560 (.L_HI(net560));
 sg13g2_tiehi _16487__561 (.L_HI(net561));
 sg13g2_tiehi _16488__562 (.L_HI(net562));
 sg13g2_tiehi _16489__563 (.L_HI(net563));
 sg13g2_tiehi _16490__564 (.L_HI(net564));
 sg13g2_tiehi _16491__565 (.L_HI(net565));
 sg13g2_tiehi _16492__566 (.L_HI(net566));
 sg13g2_tiehi _16493__567 (.L_HI(net567));
 sg13g2_tiehi _16494__568 (.L_HI(net568));
 sg13g2_tiehi _16495__569 (.L_HI(net569));
 sg13g2_tiehi _16496__570 (.L_HI(net570));
 sg13g2_tiehi _16497__571 (.L_HI(net571));
 sg13g2_tiehi _16498__572 (.L_HI(net572));
 sg13g2_tiehi _16499__573 (.L_HI(net573));
 sg13g2_tiehi _16500__574 (.L_HI(net574));
 sg13g2_tiehi _16501__575 (.L_HI(net575));
 sg13g2_tiehi _16502__576 (.L_HI(net576));
 sg13g2_tiehi _16503__577 (.L_HI(net577));
 sg13g2_tiehi _16504__578 (.L_HI(net578));
 sg13g2_tiehi _16505__579 (.L_HI(net579));
 sg13g2_tiehi _16506__580 (.L_HI(net580));
 sg13g2_tiehi _16507__581 (.L_HI(net581));
 sg13g2_tiehi _16508__582 (.L_HI(net582));
 sg13g2_tiehi _16509__583 (.L_HI(net583));
 sg13g2_tiehi _16875__584 (.L_HI(net584));
 sg13g2_tiehi _16874__585 (.L_HI(net585));
 sg13g2_tiehi _16873__586 (.L_HI(net586));
 sg13g2_tiehi _16872__587 (.L_HI(net587));
 sg13g2_tiehi _16871__588 (.L_HI(net588));
 sg13g2_tiehi _16870__589 (.L_HI(net589));
 sg13g2_tiehi _16869__590 (.L_HI(net590));
 sg13g2_tiehi _16868__591 (.L_HI(net591));
 sg13g2_tiehi _16867__592 (.L_HI(net592));
 sg13g2_tiehi _16866__593 (.L_HI(net593));
 sg13g2_tiehi _16865__594 (.L_HI(net594));
 sg13g2_tiehi _16864__595 (.L_HI(net595));
 sg13g2_tiehi _16863__596 (.L_HI(net596));
 sg13g2_tiehi _16862__597 (.L_HI(net597));
 sg13g2_tiehi _16861__598 (.L_HI(net598));
 sg13g2_tiehi _16860__599 (.L_HI(net599));
 sg13g2_tiehi _16859__600 (.L_HI(net600));
 sg13g2_tiehi _16858__601 (.L_HI(net601));
 sg13g2_tiehi _16857__602 (.L_HI(net602));
 sg13g2_tiehi _16856__603 (.L_HI(net603));
 sg13g2_tiehi _16855__604 (.L_HI(net604));
 sg13g2_tiehi _16854__605 (.L_HI(net605));
 sg13g2_tiehi _16853__606 (.L_HI(net606));
 sg13g2_tiehi _16829__607 (.L_HI(net607));
 sg13g2_tiehi _17282__608 (.L_HI(net608));
 sg13g2_tiehi _16828__609 (.L_HI(net609));
 sg13g2_tiehi _17226__610 (.L_HI(net610));
 sg13g2_tiehi _16823__611 (.L_HI(net611));
 sg13g2_tiehi _17312__612 (.L_HI(net612));
 sg13g2_tiehi _16822__613 (.L_HI(net613));
 sg13g2_tiehi _17225__614 (.L_HI(net614));
 sg13g2_tiehi _16821__615 (.L_HI(net615));
 sg13g2_tiehi _17281__616 (.L_HI(net616));
 sg13g2_tiehi _16820__617 (.L_HI(net617));
 sg13g2_tiehi _17224__618 (.L_HI(net618));
 sg13g2_tiehi _16819__619 (.L_HI(net619));
 sg13g2_tiehi _17311__620 (.L_HI(net620));
 sg13g2_tiehi _16818__621 (.L_HI(net621));
 sg13g2_tiehi _17223__622 (.L_HI(net622));
 sg13g2_tiehi _16817__623 (.L_HI(net623));
 sg13g2_tiehi _17280__624 (.L_HI(net624));
 sg13g2_tiehi _16816__625 (.L_HI(net625));
 sg13g2_tiehi _17222__626 (.L_HI(net626));
 sg13g2_tiehi _16815__627 (.L_HI(net627));
 sg13g2_tiehi _17310__628 (.L_HI(net628));
 sg13g2_tiehi _16814__629 (.L_HI(net629));
 sg13g2_tiehi _17221__630 (.L_HI(net630));
 sg13g2_tiehi _16813__631 (.L_HI(net631));
 sg13g2_tiehi _17279__632 (.L_HI(net632));
 sg13g2_tiehi _16812__633 (.L_HI(net633));
 sg13g2_tiehi _17220__634 (.L_HI(net634));
 sg13g2_tiehi _16811__635 (.L_HI(net635));
 sg13g2_tiehi _17309__636 (.L_HI(net636));
 sg13g2_tiehi _16810__637 (.L_HI(net637));
 sg13g2_tiehi _17219__638 (.L_HI(net638));
 sg13g2_tiehi _16809__639 (.L_HI(net639));
 sg13g2_tiehi _17278__640 (.L_HI(net640));
 sg13g2_tiehi _16808__641 (.L_HI(net641));
 sg13g2_tiehi _17218__642 (.L_HI(net642));
 sg13g2_tiehi _16807__643 (.L_HI(net643));
 sg13g2_tiehi _17257__644 (.L_HI(net644));
 sg13g2_tiehi _16806__645 (.L_HI(net645));
 sg13g2_tiehi _17217__646 (.L_HI(net646));
 sg13g2_tiehi _16805__647 (.L_HI(net647));
 sg13g2_tiehi _17277__648 (.L_HI(net648));
 sg13g2_tiehi _16804__649 (.L_HI(net649));
 sg13g2_tiehi _17216__650 (.L_HI(net650));
 sg13g2_tiehi _16803__651 (.L_HI(net651));
 sg13g2_tiehi _17308__652 (.L_HI(net652));
 sg13g2_tiehi _16802__653 (.L_HI(net653));
 sg13g2_tiehi _17215__654 (.L_HI(net654));
 sg13g2_tiehi _16801__655 (.L_HI(net655));
 sg13g2_tiehi _17276__656 (.L_HI(net656));
 sg13g2_tiehi _16800__657 (.L_HI(net657));
 sg13g2_tiehi _17214__658 (.L_HI(net658));
 sg13g2_tiehi _16799__659 (.L_HI(net659));
 sg13g2_tiehi _17328__660 (.L_HI(net660));
 sg13g2_tiehi _16798__661 (.L_HI(net661));
 sg13g2_tiehi _17213__662 (.L_HI(net662));
 sg13g2_tiehi _16797__663 (.L_HI(net663));
 sg13g2_tiehi _17275__664 (.L_HI(net664));
 sg13g2_tiehi _16796__665 (.L_HI(net665));
 sg13g2_tiehi _17212__666 (.L_HI(net666));
 sg13g2_tiehi _16795__667 (.L_HI(net667));
 sg13g2_tiehi _17307__668 (.L_HI(net668));
 sg13g2_tiehi _16794__669 (.L_HI(net669));
 sg13g2_tiehi _17211__670 (.L_HI(net670));
 sg13g2_tiehi _16793__671 (.L_HI(net671));
 sg13g2_tiehi _17274__672 (.L_HI(net672));
 sg13g2_tiehi _16792__673 (.L_HI(net673));
 sg13g2_tiehi _17210__674 (.L_HI(net674));
 sg13g2_tiehi _16791__675 (.L_HI(net675));
 sg13g2_tiehi _17335__676 (.L_HI(net676));
 sg13g2_tiehi _16790__677 (.L_HI(net677));
 sg13g2_tiehi _17209__678 (.L_HI(net678));
 sg13g2_tiehi _16789__679 (.L_HI(net679));
 sg13g2_tiehi _16788__680 (.L_HI(net680));
 sg13g2_tiehi _17273__681 (.L_HI(net681));
 sg13g2_tiehi _16787__682 (.L_HI(net682));
 sg13g2_tiehi _17208__683 (.L_HI(net683));
 sg13g2_tiehi _16786__684 (.L_HI(net684));
 sg13g2_tiehi _17306__685 (.L_HI(net685));
 sg13g2_tiehi _16785__686 (.L_HI(net686));
 sg13g2_tiehi _17207__687 (.L_HI(net687));
 sg13g2_tiehi _16784__688 (.L_HI(net688));
 sg13g2_tiehi _17272__689 (.L_HI(net689));
 sg13g2_tiehi _16783__690 (.L_HI(net690));
 sg13g2_tiehi _17206__691 (.L_HI(net691));
 sg13g2_tiehi _16782__692 (.L_HI(net692));
 sg13g2_tiehi _17327__693 (.L_HI(net693));
 sg13g2_tiehi _16781__694 (.L_HI(net694));
 sg13g2_tiehi _17205__695 (.L_HI(net695));
 sg13g2_tiehi _16780__696 (.L_HI(net696));
 sg13g2_tiehi _17271__697 (.L_HI(net697));
 sg13g2_tiehi _16779__698 (.L_HI(net698));
 sg13g2_tiehi _17204__699 (.L_HI(net699));
 sg13g2_tiehi _16778__700 (.L_HI(net700));
 sg13g2_tiehi _17305__701 (.L_HI(net701));
 sg13g2_tiehi _16777__702 (.L_HI(net702));
 sg13g2_tiehi _17203__703 (.L_HI(net703));
 sg13g2_tiehi _16776__704 (.L_HI(net704));
 sg13g2_tiehi _17270__705 (.L_HI(net705));
 sg13g2_tiehi _16775__706 (.L_HI(net706));
 sg13g2_tiehi _17202__707 (.L_HI(net707));
 sg13g2_tiehi _16774__708 (.L_HI(net708));
 sg13g2_tiehi _17334__709 (.L_HI(net709));
 sg13g2_tiehi _16773__710 (.L_HI(net710));
 sg13g2_tiehi _17201__711 (.L_HI(net711));
 sg13g2_tiehi _16772__712 (.L_HI(net712));
 sg13g2_tiehi _17269__713 (.L_HI(net713));
 sg13g2_tiehi _16771__714 (.L_HI(net714));
 sg13g2_tiehi _17200__715 (.L_HI(net715));
 sg13g2_tiehi _16770__716 (.L_HI(net716));
 sg13g2_tiehi _17304__717 (.L_HI(net717));
 sg13g2_tiehi _16769__718 (.L_HI(net718));
 sg13g2_tiehi _17199__719 (.L_HI(net719));
 sg13g2_tiehi _16768__720 (.L_HI(net720));
 sg13g2_tiehi _17198__721 (.L_HI(net721));
 sg13g2_tiehi _16767__722 (.L_HI(net722));
 sg13g2_tiehi _17197__723 (.L_HI(net723));
 sg13g2_tiehi _16766__724 (.L_HI(net724));
 sg13g2_tiehi _17196__725 (.L_HI(net725));
 sg13g2_tiehi _16765__726 (.L_HI(net726));
 sg13g2_tiehi _17195__727 (.L_HI(net727));
 sg13g2_tiehi _16764__728 (.L_HI(net728));
 sg13g2_tiehi _17194__729 (.L_HI(net729));
 sg13g2_tiehi _16763__730 (.L_HI(net730));
 sg13g2_tiehi _17193__731 (.L_HI(net731));
 sg13g2_tiehi _16762__732 (.L_HI(net732));
 sg13g2_tiehi _17192__733 (.L_HI(net733));
 sg13g2_tiehi _16761__734 (.L_HI(net734));
 sg13g2_tiehi _17191__735 (.L_HI(net735));
 sg13g2_tiehi _16760__736 (.L_HI(net736));
 sg13g2_tiehi _17190__737 (.L_HI(net737));
 sg13g2_tiehi _16759__738 (.L_HI(net738));
 sg13g2_tiehi _17189__739 (.L_HI(net739));
 sg13g2_tiehi _16758__740 (.L_HI(net740));
 sg13g2_tiehi _17188__741 (.L_HI(net741));
 sg13g2_tiehi _16757__742 (.L_HI(net742));
 sg13g2_tiehi _17187__743 (.L_HI(net743));
 sg13g2_tiehi _16756__744 (.L_HI(net744));
 sg13g2_tiehi _17186__745 (.L_HI(net745));
 sg13g2_tiehi _16755__746 (.L_HI(net746));
 sg13g2_tiehi _17185__747 (.L_HI(net747));
 sg13g2_tiehi _16754__748 (.L_HI(net748));
 sg13g2_tiehi _17184__749 (.L_HI(net749));
 sg13g2_tiehi _16753__750 (.L_HI(net750));
 sg13g2_tiehi _17183__751 (.L_HI(net751));
 sg13g2_tiehi _16752__752 (.L_HI(net752));
 sg13g2_tiehi _17182__753 (.L_HI(net753));
 sg13g2_tiehi _16751__754 (.L_HI(net754));
 sg13g2_tiehi _17181__755 (.L_HI(net755));
 sg13g2_tiehi _16750__756 (.L_HI(net756));
 sg13g2_tiehi _17180__757 (.L_HI(net757));
 sg13g2_tiehi _16749__758 (.L_HI(net758));
 sg13g2_tiehi _17179__759 (.L_HI(net759));
 sg13g2_tiehi _16748__760 (.L_HI(net760));
 sg13g2_tiehi _17178__761 (.L_HI(net761));
 sg13g2_tiehi _16747__762 (.L_HI(net762));
 sg13g2_tiehi _17177__763 (.L_HI(net763));
 sg13g2_tiehi _16746__764 (.L_HI(net764));
 sg13g2_tiehi _17176__765 (.L_HI(net765));
 sg13g2_tiehi _16745__766 (.L_HI(net766));
 sg13g2_tiehi _17175__767 (.L_HI(net767));
 sg13g2_tiehi _16744__768 (.L_HI(net768));
 sg13g2_tiehi _17174__769 (.L_HI(net769));
 sg13g2_tiehi _16743__770 (.L_HI(net770));
 sg13g2_tiehi _17173__771 (.L_HI(net771));
 sg13g2_tiehi _16742__772 (.L_HI(net772));
 sg13g2_tiehi _17172__773 (.L_HI(net773));
 sg13g2_tiehi _16741__774 (.L_HI(net774));
 sg13g2_tiehi _16740__775 (.L_HI(net775));
 sg13g2_tiehi _16739__776 (.L_HI(net776));
 sg13g2_tiehi _16738__777 (.L_HI(net777));
 sg13g2_tiehi _16737__778 (.L_HI(net778));
 sg13g2_tiehi _16736__779 (.L_HI(net779));
 sg13g2_tiehi _16735__780 (.L_HI(net780));
 sg13g2_tiehi _16734__781 (.L_HI(net781));
 sg13g2_tiehi _16733__782 (.L_HI(net782));
 sg13g2_tiehi _16732__783 (.L_HI(net783));
 sg13g2_tiehi _16731__784 (.L_HI(net784));
 sg13g2_tiehi _16730__785 (.L_HI(net785));
 sg13g2_tiehi _16729__786 (.L_HI(net786));
 sg13g2_tiehi _16728__787 (.L_HI(net787));
 sg13g2_tiehi _16727__788 (.L_HI(net788));
 sg13g2_tiehi _16726__789 (.L_HI(net789));
 sg13g2_tiehi _16725__790 (.L_HI(net790));
 sg13g2_tiehi _16724__791 (.L_HI(net791));
 sg13g2_tiehi _16723__792 (.L_HI(net792));
 sg13g2_tiehi _16722__793 (.L_HI(net793));
 sg13g2_tiehi _16721__794 (.L_HI(net794));
 sg13g2_tiehi _16720__795 (.L_HI(net795));
 sg13g2_tiehi _17171__796 (.L_HI(net796));
 sg13g2_tiehi _16719__797 (.L_HI(net797));
 sg13g2_tiehi _17170__798 (.L_HI(net798));
 sg13g2_tiehi _16718__799 (.L_HI(net799));
 sg13g2_tiehi _17169__800 (.L_HI(net800));
 sg13g2_tiehi _16717__801 (.L_HI(net801));
 sg13g2_tiehi _17168__802 (.L_HI(net802));
 sg13g2_tiehi _16716__803 (.L_HI(net803));
 sg13g2_tiehi _16715__804 (.L_HI(net804));
 sg13g2_tiehi _17167__805 (.L_HI(net805));
 sg13g2_tiehi _16714__806 (.L_HI(net806));
 sg13g2_tiehi _16713__807 (.L_HI(net807));
 sg13g2_tiehi _16712__808 (.L_HI(net808));
 sg13g2_tiehi _16711__809 (.L_HI(net809));
 sg13g2_tiehi _16710__810 (.L_HI(net810));
 sg13g2_tiehi _16709__811 (.L_HI(net811));
 sg13g2_tiehi _16708__812 (.L_HI(net812));
 sg13g2_tiehi _16707__813 (.L_HI(net813));
 sg13g2_tiehi _16706__814 (.L_HI(net814));
 sg13g2_tiehi _17268__815 (.L_HI(net815));
 sg13g2_tiehi _16705__816 (.L_HI(net816));
 sg13g2_tiehi _17166__817 (.L_HI(net817));
 sg13g2_tiehi _16704__818 (.L_HI(net818));
 sg13g2_tiehi _17326__819 (.L_HI(net819));
 sg13g2_tiehi _16703__820 (.L_HI(net820));
 sg13g2_tiehi _17165__821 (.L_HI(net821));
 sg13g2_tiehi _16702__822 (.L_HI(net822));
 sg13g2_tiehi _17267__823 (.L_HI(net823));
 sg13g2_tiehi _16701__824 (.L_HI(net824));
 sg13g2_tiehi _17164__825 (.L_HI(net825));
 sg13g2_tiehi _16700__826 (.L_HI(net826));
 sg13g2_tiehi _17163__827 (.L_HI(net827));
 sg13g2_tiehi _16699__828 (.L_HI(net828));
 sg13g2_tiehi _17162__829 (.L_HI(net829));
 sg13g2_tiehi _16698__830 (.L_HI(net830));
 sg13g2_tiehi _17161__831 (.L_HI(net831));
 sg13g2_tiehi _16697__832 (.L_HI(net832));
 sg13g2_tiehi _17160__833 (.L_HI(net833));
 sg13g2_tiehi _16696__834 (.L_HI(net834));
 sg13g2_tiehi _17159__835 (.L_HI(net835));
 sg13g2_tiehi _16695__836 (.L_HI(net836));
 sg13g2_tiehi _17158__837 (.L_HI(net837));
 sg13g2_tiehi _16694__838 (.L_HI(net838));
 sg13g2_tiehi _17157__839 (.L_HI(net839));
 sg13g2_tiehi _16693__840 (.L_HI(net840));
 sg13g2_tiehi _17156__841 (.L_HI(net841));
 sg13g2_tiehi _16692__842 (.L_HI(net842));
 sg13g2_tiehi _17155__843 (.L_HI(net843));
 sg13g2_tiehi _16691__844 (.L_HI(net844));
 sg13g2_tiehi _17154__845 (.L_HI(net845));
 sg13g2_tiehi _16690__846 (.L_HI(net846));
 sg13g2_tiehi _17153__847 (.L_HI(net847));
 sg13g2_tiehi _16689__848 (.L_HI(net848));
 sg13g2_tiehi _17152__849 (.L_HI(net849));
 sg13g2_tiehi _16688__850 (.L_HI(net850));
 sg13g2_tiehi _17151__851 (.L_HI(net851));
 sg13g2_tiehi _16687__852 (.L_HI(net852));
 sg13g2_tiehi _17150__853 (.L_HI(net853));
 sg13g2_tiehi _16686__854 (.L_HI(net854));
 sg13g2_tiehi _17149__855 (.L_HI(net855));
 sg13g2_tiehi _16685__856 (.L_HI(net856));
 sg13g2_tiehi _17148__857 (.L_HI(net857));
 sg13g2_tiehi _16684__858 (.L_HI(net858));
 sg13g2_tiehi _17147__859 (.L_HI(net859));
 sg13g2_tiehi _16683__860 (.L_HI(net860));
 sg13g2_tiehi _17146__861 (.L_HI(net861));
 sg13g2_tiehi _16682__862 (.L_HI(net862));
 sg13g2_tiehi _17145__863 (.L_HI(net863));
 sg13g2_tiehi _16681__864 (.L_HI(net864));
 sg13g2_tiehi _17144__865 (.L_HI(net865));
 sg13g2_tiehi _16680__866 (.L_HI(net866));
 sg13g2_tiehi _16679__867 (.L_HI(net867));
 sg13g2_tiehi _16678__868 (.L_HI(net868));
 sg13g2_tiehi _17143__869 (.L_HI(net869));
 sg13g2_tiehi _16677__870 (.L_HI(net870));
 sg13g2_tiehi _17142__871 (.L_HI(net871));
 sg13g2_tiehi _16676__872 (.L_HI(net872));
 sg13g2_tiehi _17141__873 (.L_HI(net873));
 sg13g2_tiehi _16675__874 (.L_HI(net874));
 sg13g2_tiehi _17140__875 (.L_HI(net875));
 sg13g2_tiehi _16674__876 (.L_HI(net876));
 sg13g2_tiehi _17139__877 (.L_HI(net877));
 sg13g2_tiehi _16673__878 (.L_HI(net878));
 sg13g2_tiehi _17138__879 (.L_HI(net879));
 sg13g2_tiehi _16672__880 (.L_HI(net880));
 sg13g2_tiehi _17137__881 (.L_HI(net881));
 sg13g2_tiehi _16671__882 (.L_HI(net882));
 sg13g2_tiehi _17136__883 (.L_HI(net883));
 sg13g2_tiehi _16670__884 (.L_HI(net884));
 sg13g2_tiehi _17135__885 (.L_HI(net885));
 sg13g2_tiehi _16669__886 (.L_HI(net886));
 sg13g2_tiehi _17134__887 (.L_HI(net887));
 sg13g2_tiehi _16668__888 (.L_HI(net888));
 sg13g2_tiehi _17133__889 (.L_HI(net889));
 sg13g2_tiehi _16667__890 (.L_HI(net890));
 sg13g2_tiehi _16666__891 (.L_HI(net891));
 sg13g2_tiehi _16665__892 (.L_HI(net892));
 sg13g2_tiehi _17303__893 (.L_HI(net893));
 sg13g2_tiehi _16664__894 (.L_HI(net894));
 sg13g2_tiehi _17132__895 (.L_HI(net895));
 sg13g2_tiehi _16663__896 (.L_HI(net896));
 sg13g2_tiehi _16510__897 (.L_HI(net897));
 sg13g2_tiehi _16824__898 (.L_HI(net898));
 sg13g2_tiehi _16825__899 (.L_HI(net899));
 sg13g2_tiehi _16826__900 (.L_HI(net900));
 sg13g2_tiehi _16662__901 (.L_HI(net901));
 sg13g2_tiehi _16661__902 (.L_HI(net902));
 sg13g2_tiehi _16827__903 (.L_HI(net903));
 sg13g2_tiehi _16830__904 (.L_HI(net904));
 sg13g2_tiehi _16831__905 (.L_HI(net905));
 sg13g2_tiehi _16832__906 (.L_HI(net906));
 sg13g2_tiehi _16833__907 (.L_HI(net907));
 sg13g2_tiehi _16834__908 (.L_HI(net908));
 sg13g2_tiehi _16835__909 (.L_HI(net909));
 sg13g2_tiehi _16836__910 (.L_HI(net910));
 sg13g2_tiehi _16837__911 (.L_HI(net911));
 sg13g2_tiehi _16838__912 (.L_HI(net912));
 sg13g2_tiehi _16839__913 (.L_HI(net913));
 sg13g2_tiehi _16840__914 (.L_HI(net914));
 sg13g2_tiehi _16841__915 (.L_HI(net915));
 sg13g2_tiehi _16842__916 (.L_HI(net916));
 sg13g2_tiehi _16843__917 (.L_HI(net917));
 sg13g2_tiehi _16844__918 (.L_HI(net918));
 sg13g2_tiehi _16845__919 (.L_HI(net919));
 sg13g2_tiehi _16846__920 (.L_HI(net920));
 sg13g2_tiehi _16847__921 (.L_HI(net921));
 sg13g2_tiehi _16848__922 (.L_HI(net922));
 sg13g2_tiehi _16849__923 (.L_HI(net923));
 sg13g2_tiehi _16850__924 (.L_HI(net924));
 sg13g2_tiehi _16851__925 (.L_HI(net925));
 sg13g2_tiehi _16660__926 (.L_HI(net926));
 sg13g2_tiehi _16659__927 (.L_HI(net927));
 sg13g2_tiehi _16658__928 (.L_HI(net928));
 sg13g2_tiehi _16657__929 (.L_HI(net929));
 sg13g2_tiehi _16656__930 (.L_HI(net930));
 sg13g2_tiehi _16655__931 (.L_HI(net931));
 sg13g2_tiehi _16654__932 (.L_HI(net932));
 sg13g2_tiehi _16653__933 (.L_HI(net933));
 sg13g2_tiehi _16652__934 (.L_HI(net934));
 sg13g2_tiehi _16651__935 (.L_HI(net935));
 sg13g2_tiehi _16650__936 (.L_HI(net936));
 sg13g2_tiehi _16649__937 (.L_HI(net937));
 sg13g2_tiehi _16648__938 (.L_HI(net938));
 sg13g2_tiehi _16647__939 (.L_HI(net939));
 sg13g2_tiehi _16646__940 (.L_HI(net940));
 sg13g2_tiehi _16645__941 (.L_HI(net941));
 sg13g2_tiehi _16644__942 (.L_HI(net942));
 sg13g2_tiehi _16643__943 (.L_HI(net943));
 sg13g2_tiehi _16642__944 (.L_HI(net944));
 sg13g2_tiehi _16641__945 (.L_HI(net945));
 sg13g2_tiehi _16640__946 (.L_HI(net946));
 sg13g2_tiehi _16639__947 (.L_HI(net947));
 sg13g2_tiehi _16638__948 (.L_HI(net948));
 sg13g2_tiehi _16637__949 (.L_HI(net949));
 sg13g2_tiehi _16636__950 (.L_HI(net950));
 sg13g2_tiehi _16635__951 (.L_HI(net951));
 sg13g2_tiehi _16634__952 (.L_HI(net952));
 sg13g2_tiehi _16633__953 (.L_HI(net953));
 sg13g2_tiehi _16632__954 (.L_HI(net954));
 sg13g2_tiehi _16631__955 (.L_HI(net955));
 sg13g2_tiehi _16630__956 (.L_HI(net956));
 sg13g2_tiehi _16629__957 (.L_HI(net957));
 sg13g2_tiehi _16628__958 (.L_HI(net958));
 sg13g2_tiehi _16852__959 (.L_HI(net959));
 sg13g2_tiehi _16886__960 (.L_HI(net960));
 sg13g2_tiehi _16887__961 (.L_HI(net961));
 sg13g2_tiehi _16888__962 (.L_HI(net962));
 sg13g2_tiehi _16889__963 (.L_HI(net963));
 sg13g2_tiehi _16890__964 (.L_HI(net964));
 sg13g2_tiehi _16891__965 (.L_HI(net965));
 sg13g2_tiehi _16892__966 (.L_HI(net966));
 sg13g2_tiehi _16893__967 (.L_HI(net967));
 sg13g2_tiehi _16894__968 (.L_HI(net968));
 sg13g2_tiehi _16895__969 (.L_HI(net969));
 sg13g2_tiehi _16896__970 (.L_HI(net970));
 sg13g2_tiehi _16627__971 (.L_HI(net971));
 sg13g2_tiehi _16626__972 (.L_HI(net972));
 sg13g2_tiehi _16625__973 (.L_HI(net973));
 sg13g2_tiehi _16624__974 (.L_HI(net974));
 sg13g2_tiehi _16623__975 (.L_HI(net975));
 sg13g2_tiehi _16622__976 (.L_HI(net976));
 sg13g2_tiehi _16621__977 (.L_HI(net977));
 sg13g2_tiehi _16620__978 (.L_HI(net978));
 sg13g2_tiehi _16619__979 (.L_HI(net979));
 sg13g2_tiehi _16618__980 (.L_HI(net980));
 sg13g2_tiehi _16617__981 (.L_HI(net981));
 sg13g2_tiehi _16616__982 (.L_HI(net982));
 sg13g2_tiehi _16615__983 (.L_HI(net983));
 sg13g2_tiehi _16614__984 (.L_HI(net984));
 sg13g2_tiehi _16613__985 (.L_HI(net985));
 sg13g2_tiehi _16612__986 (.L_HI(net986));
 sg13g2_tiehi _16611__987 (.L_HI(net987));
 sg13g2_tiehi _16610__988 (.L_HI(net988));
 sg13g2_tiehi _16609__989 (.L_HI(net989));
 sg13g2_tiehi _16608__990 (.L_HI(net990));
 sg13g2_tiehi _16607__991 (.L_HI(net991));
 sg13g2_tiehi _16606__992 (.L_HI(net992));
 sg13g2_tiehi _16605__993 (.L_HI(net993));
 sg13g2_tiehi _16604__994 (.L_HI(net994));
 sg13g2_tiehi _16603__995 (.L_HI(net995));
 sg13g2_tiehi _16602__996 (.L_HI(net996));
 sg13g2_tiehi _16601__997 (.L_HI(net997));
 sg13g2_tiehi _16600__998 (.L_HI(net998));
 sg13g2_tiehi _16599__999 (.L_HI(net999));
 sg13g2_tiehi _16598__1000 (.L_HI(net1000));
 sg13g2_tiehi _17266__1001 (.L_HI(net1001));
 sg13g2_tiehi _16597__1002 (.L_HI(net1002));
 sg13g2_tiehi _17131__1003 (.L_HI(net1003));
 sg13g2_tiehi _16596__1004 (.L_HI(net1004));
 sg13g2_tiehi _17333__1005 (.L_HI(net1005));
 sg13g2_tiehi _16595__1006 (.L_HI(net1006));
 sg13g2_tiehi _17130__1007 (.L_HI(net1007));
 sg13g2_tiehi _16594__1008 (.L_HI(net1008));
 sg13g2_tiehi _17265__1009 (.L_HI(net1009));
 sg13g2_tiehi _16593__1010 (.L_HI(net1010));
 sg13g2_tiehi _17129__1011 (.L_HI(net1011));
 sg13g2_tiehi _16592__1012 (.L_HI(net1012));
 sg13g2_tiehi _17302__1013 (.L_HI(net1013));
 sg13g2_tiehi _16591__1014 (.L_HI(net1014));
 sg13g2_tiehi _17128__1015 (.L_HI(net1015));
 sg13g2_tiehi _16590__1016 (.L_HI(net1016));
 sg13g2_tiehi _17264__1017 (.L_HI(net1017));
 sg13g2_tiehi _16589__1018 (.L_HI(net1018));
 sg13g2_tiehi _17127__1019 (.L_HI(net1019));
 sg13g2_tiehi _16588__1020 (.L_HI(net1020));
 sg13g2_tiehi _17325__1021 (.L_HI(net1021));
 sg13g2_tiehi _16587__1022 (.L_HI(net1022));
 sg13g2_tiehi _17126__1023 (.L_HI(net1023));
 sg13g2_tiehi _16586__1024 (.L_HI(net1024));
 sg13g2_tiehi _17263__1025 (.L_HI(net1025));
 sg13g2_tiehi _16585__1026 (.L_HI(net1026));
 sg13g2_tiehi _17125__1027 (.L_HI(net1027));
 sg13g2_tiehi _16584__1028 (.L_HI(net1028));
 sg13g2_tiehi _17301__1029 (.L_HI(net1029));
 sg13g2_tiehi _16583__1030 (.L_HI(net1030));
 sg13g2_tiehi _17124__1031 (.L_HI(net1031));
 sg13g2_tiehi _16582__1032 (.L_HI(net1032));
 sg13g2_tiehi _17123__1033 (.L_HI(net1033));
 sg13g2_tiehi _16581__1034 (.L_HI(net1034));
 sg13g2_tiehi _17262__1035 (.L_HI(net1035));
 sg13g2_tiehi _16580__1036 (.L_HI(net1036));
 sg13g2_tiehi _17122__1037 (.L_HI(net1037));
 sg13g2_tiehi _16579__1038 (.L_HI(net1038));
 sg13g2_tiehi _17332__1039 (.L_HI(net1039));
 sg13g2_tiehi _16578__1040 (.L_HI(net1040));
 sg13g2_tiehi _17121__1041 (.L_HI(net1041));
 sg13g2_tiehi _16577__1042 (.L_HI(net1042));
 sg13g2_tiehi _17261__1043 (.L_HI(net1043));
 sg13g2_tiehi _16576__1044 (.L_HI(net1044));
 sg13g2_tiehi _17120__1045 (.L_HI(net1045));
 sg13g2_tiehi _16575__1046 (.L_HI(net1046));
 sg13g2_tiehi _17300__1047 (.L_HI(net1047));
 sg13g2_tiehi _16574__1048 (.L_HI(net1048));
 sg13g2_tiehi _17119__1049 (.L_HI(net1049));
 sg13g2_tiehi _16573__1050 (.L_HI(net1050));
 sg13g2_tiehi _17260__1051 (.L_HI(net1051));
 sg13g2_tiehi _16572__1052 (.L_HI(net1052));
 sg13g2_tiehi _17118__1053 (.L_HI(net1053));
 sg13g2_tiehi _16571__1054 (.L_HI(net1054));
 sg13g2_tiehi _17324__1055 (.L_HI(net1055));
 sg13g2_tiehi _16570__1056 (.L_HI(net1056));
 sg13g2_tiehi _17117__1057 (.L_HI(net1057));
 sg13g2_tiehi _16569__1058 (.L_HI(net1058));
 sg13g2_tiehi _17259__1059 (.L_HI(net1059));
 sg13g2_tiehi _16568__1060 (.L_HI(net1060));
 sg13g2_tiehi _17116__1061 (.L_HI(net1061));
 sg13g2_tiehi _16567__1062 (.L_HI(net1062));
 sg13g2_tiehi _17115__1063 (.L_HI(net1063));
 sg13g2_tiehi _16566__1064 (.L_HI(net1064));
 sg13g2_tiehi _17114__1065 (.L_HI(net1065));
 sg13g2_tiehi _16565__1066 (.L_HI(net1066));
 sg13g2_tiehi _17113__1067 (.L_HI(net1067));
 sg13g2_tiehi _16564__1068 (.L_HI(net1068));
 sg13g2_tiehi _17299__1069 (.L_HI(net1069));
 sg13g2_tiehi _16563__1070 (.L_HI(net1070));
 sg13g2_tiehi _17112__1071 (.L_HI(net1071));
 sg13g2_tiehi _16562__1072 (.L_HI(net1072));
 sg13g2_tiehi _17111__1073 (.L_HI(net1073));
 sg13g2_tiehi _16561__1074 (.L_HI(net1074));
 sg13g2_tiehi _17110__1075 (.L_HI(net1075));
 sg13g2_tiehi _16560__1076 (.L_HI(net1076));
 sg13g2_tiehi _17109__1077 (.L_HI(net1077));
 sg13g2_tiehi _16559__1078 (.L_HI(net1078));
 sg13g2_tiehi _17108__1079 (.L_HI(net1079));
 sg13g2_tiehi _16558__1080 (.L_HI(net1080));
 sg13g2_tiehi _17107__1081 (.L_HI(net1081));
 sg13g2_tiehi _16557__1082 (.L_HI(net1082));
 sg13g2_tiehi _17106__1083 (.L_HI(net1083));
 sg13g2_tiehi _16556__1084 (.L_HI(net1084));
 sg13g2_tiehi _17105__1085 (.L_HI(net1085));
 sg13g2_tiehi _16555__1086 (.L_HI(net1086));
 sg13g2_tiehi _17104__1087 (.L_HI(net1087));
 sg13g2_tiehi _16554__1088 (.L_HI(net1088));
 sg13g2_tiehi _17103__1089 (.L_HI(net1089));
 sg13g2_tiehi _16553__1090 (.L_HI(net1090));
 sg13g2_tiehi _17102__1091 (.L_HI(net1091));
 sg13g2_tiehi _16552__1092 (.L_HI(net1092));
 sg13g2_tiehi _17101__1093 (.L_HI(net1093));
 sg13g2_tiehi _16551__1094 (.L_HI(net1094));
 sg13g2_tiehi _17100__1095 (.L_HI(net1095));
 sg13g2_tiehi _16550__1096 (.L_HI(net1096));
 sg13g2_tiehi _17099__1097 (.L_HI(net1097));
 sg13g2_tiehi _16549__1098 (.L_HI(net1098));
 sg13g2_tiehi _17098__1099 (.L_HI(net1099));
 sg13g2_tiehi _16548__1100 (.L_HI(net1100));
 sg13g2_tiehi _17097__1101 (.L_HI(net1101));
 sg13g2_tiehi _16547__1102 (.L_HI(net1102));
 sg13g2_tiehi _17096__1103 (.L_HI(net1103));
 sg13g2_tiehi _16546__1104 (.L_HI(net1104));
 sg13g2_tiehi _17095__1105 (.L_HI(net1105));
 sg13g2_tiehi _16545__1106 (.L_HI(net1106));
 sg13g2_tiehi _17094__1107 (.L_HI(net1107));
 sg13g2_tiehi _16544__1108 (.L_HI(net1108));
 sg13g2_tiehi _17093__1109 (.L_HI(net1109));
 sg13g2_tiehi _16543__1110 (.L_HI(net1110));
 sg13g2_tiehi _17092__1111 (.L_HI(net1111));
 sg13g2_tiehi _16542__1112 (.L_HI(net1112));
 sg13g2_tiehi _17091__1113 (.L_HI(net1113));
 sg13g2_tiehi _16541__1114 (.L_HI(net1114));
 sg13g2_tiehi _17090__1115 (.L_HI(net1115));
 sg13g2_tiehi _16540__1116 (.L_HI(net1116));
 sg13g2_tiehi _17089__1117 (.L_HI(net1117));
 sg13g2_tiehi _16539__1118 (.L_HI(net1118));
 sg13g2_tiehi _17088__1119 (.L_HI(net1119));
 sg13g2_tiehi _16538__1120 (.L_HI(net1120));
 sg13g2_tiehi _17087__1121 (.L_HI(net1121));
 sg13g2_tiehi _16537__1122 (.L_HI(net1122));
 sg13g2_tiehi _17086__1123 (.L_HI(net1123));
 sg13g2_tiehi _16536__1124 (.L_HI(net1124));
 sg13g2_tiehi _17085__1125 (.L_HI(net1125));
 sg13g2_tiehi _16535__1126 (.L_HI(net1126));
 sg13g2_tiehi _17084__1127 (.L_HI(net1127));
 sg13g2_tiehi _16534__1128 (.L_HI(net1128));
 sg13g2_tiehi _17083__1129 (.L_HI(net1129));
 sg13g2_tiehi _16533__1130 (.L_HI(net1130));
 sg13g2_tiehi _17082__1131 (.L_HI(net1131));
 sg13g2_tiehi _16532__1132 (.L_HI(net1132));
 sg13g2_tiehi _17081__1133 (.L_HI(net1133));
 sg13g2_tiehi _16531__1134 (.L_HI(net1134));
 sg13g2_tiehi _17080__1135 (.L_HI(net1135));
 sg13g2_tiehi _16530__1136 (.L_HI(net1136));
 sg13g2_tiehi _17079__1137 (.L_HI(net1137));
 sg13g2_tiehi _16529__1138 (.L_HI(net1138));
 sg13g2_tiehi _17258__1139 (.L_HI(net1139));
 sg13g2_tiehi _16528__1140 (.L_HI(net1140));
 sg13g2_tiehi _17078__1141 (.L_HI(net1141));
 sg13g2_tiehi _16527__1142 (.L_HI(net1142));
 sg13g2_tiehi _17331__1143 (.L_HI(net1143));
 sg13g2_tiehi _16526__1144 (.L_HI(net1144));
 sg13g2_tiehi _17077__1145 (.L_HI(net1145));
 sg13g2_tiehi _16525__1146 (.L_HI(net1146));
 sg13g2_tiehi _16897__1147 (.L_HI(net1147));
 sg13g2_tiehi _17076__1148 (.L_HI(net1148));
 sg13g2_tiehi _16524__1149 (.L_HI(net1149));
 sg13g2_tiehi _17256__1150 (.L_HI(net1150));
 sg13g2_tiehi _16523__1151 (.L_HI(net1151));
 sg13g2_tiehi _17075__1152 (.L_HI(net1152));
 sg13g2_tiehi _16522__1153 (.L_HI(net1153));
 sg13g2_tiehi _17298__1154 (.L_HI(net1154));
 sg13g2_tiehi _16521__1155 (.L_HI(net1155));
 sg13g2_tiehi _17073__1156 (.L_HI(net1156));
 sg13g2_tiehi _16520__1157 (.L_HI(net1157));
 sg13g2_tiehi _17255__1158 (.L_HI(net1158));
 sg13g2_tiehi _16519__1159 (.L_HI(net1159));
 sg13g2_tiehi _17072__1160 (.L_HI(net1160));
 sg13g2_tiehi _16518__1161 (.L_HI(net1161));
 sg13g2_tiehi _17071__1162 (.L_HI(net1162));
 sg13g2_tiehi _16517__1163 (.L_HI(net1163));
 sg13g2_tiehi _17070__1164 (.L_HI(net1164));
 sg13g2_tiehi _16516__1165 (.L_HI(net1165));
 sg13g2_tiehi _17069__1166 (.L_HI(net1166));
 sg13g2_tiehi _16515__1167 (.L_HI(net1167));
 sg13g2_tiehi _17068__1168 (.L_HI(net1168));
 sg13g2_tiehi _16514__1169 (.L_HI(net1169));
 sg13g2_tiehi _17323__1170 (.L_HI(net1170));
 sg13g2_tiehi _16513__1171 (.L_HI(net1171));
 sg13g2_tiehi _17067__1172 (.L_HI(net1172));
 sg13g2_tiehi _16512__1173 (.L_HI(net1173));
 sg13g2_tiehi _16511__1174 (.L_HI(net1174));
 sg13g2_tiehi _16481__1175 (.L_HI(net1175));
 sg13g2_tiehi _16480__1176 (.L_HI(net1176));
 sg13g2_tiehi _16479__1177 (.L_HI(net1177));
 sg13g2_tiehi _16478__1178 (.L_HI(net1178));
 sg13g2_tiehi _16477__1179 (.L_HI(net1179));
 sg13g2_tiehi _16476__1180 (.L_HI(net1180));
 sg13g2_tiehi _16475__1181 (.L_HI(net1181));
 sg13g2_tiehi _16474__1182 (.L_HI(net1182));
 sg13g2_tiehi _16473__1183 (.L_HI(net1183));
 sg13g2_tiehi _16472__1184 (.L_HI(net1184));
 sg13g2_tiehi _16471__1185 (.L_HI(net1185));
 sg13g2_tiehi _17254__1186 (.L_HI(net1186));
 sg13g2_tiehi _16470__1187 (.L_HI(net1187));
 sg13g2_tiehi _16437__1188 (.L_HI(net1188));
 sg13g2_tiehi _16436__1189 (.L_HI(net1189));
 sg13g2_tiehi _16435__1190 (.L_HI(net1190));
 sg13g2_tiehi _16434__1191 (.L_HI(net1191));
 sg13g2_tiehi _17066__1192 (.L_HI(net1192));
 sg13g2_tiehi _16433__1193 (.L_HI(net1193));
 sg13g2_tiehi _17297__1194 (.L_HI(net1194));
 sg13g2_tiehi _16432__1195 (.L_HI(net1195));
 sg13g2_tiehi _16431__1196 (.L_HI(net1196));
 sg13g2_tiehi _16429__1197 (.L_HI(net1197));
 sg13g2_tiehi _17065__1198 (.L_HI(net1198));
 sg13g2_tiehi _16428__1199 (.L_HI(net1199));
 sg13g2_tiehi _17253__1200 (.L_HI(net1200));
 sg13g2_tiehi _16427__1201 (.L_HI(net1201));
 sg13g2_tiehi _17064__1202 (.L_HI(net1202));
 sg13g2_tiehi _16426__1203 (.L_HI(net1203));
 sg13g2_tiehi _17063__1204 (.L_HI(net1204));
 sg13g2_tiehi _16425__1205 (.L_HI(net1205));
 sg13g2_tiehi _17062__1206 (.L_HI(net1206));
 sg13g2_tiehi _17061__1207 (.L_HI(net1207));
 sg13g2_tiehi _17060__1208 (.L_HI(net1208));
 sg13g2_tiehi _16423__1209 (.L_HI(net1209));
 sg13g2_tiehi _17059__1210 (.L_HI(net1210));
 sg13g2_tiehi _16422__1211 (.L_HI(net1211));
 sg13g2_tiehi _17058__1212 (.L_HI(net1212));
 sg13g2_tiehi _16421__1213 (.L_HI(net1213));
 sg13g2_tiehi _17057__1214 (.L_HI(net1214));
 sg13g2_tiehi _16420__1215 (.L_HI(net1215));
 sg13g2_tiehi _17056__1216 (.L_HI(net1216));
 sg13g2_tiehi _16419__1217 (.L_HI(net1217));
 sg13g2_tiehi _17055__1218 (.L_HI(net1218));
 sg13g2_tiehi _16418__1219 (.L_HI(net1219));
 sg13g2_tiehi _17054__1220 (.L_HI(net1220));
 sg13g2_tiehi _16417__1221 (.L_HI(net1221));
 sg13g2_tiehi _17053__1222 (.L_HI(net1222));
 sg13g2_tiehi _16415__1223 (.L_HI(net1223));
 sg13g2_tiehi _17052__1224 (.L_HI(net1224));
 sg13g2_tiehi _16414__1225 (.L_HI(net1225));
 sg13g2_tiehi _16413__1226 (.L_HI(net1226));
 sg13g2_tiehi _17051__1227 (.L_HI(net1227));
 sg13g2_tiehi _16412__1228 (.L_HI(net1228));
 sg13g2_tiehi _17050__1229 (.L_HI(net1229));
 sg13g2_tiehi _16411__1230 (.L_HI(net1230));
 sg13g2_tiehi _16410__1231 (.L_HI(net1231));
 sg13g2_tiehi _16409__1232 (.L_HI(net1232));
 sg13g2_tiehi _15995__1233 (.L_HI(net1233));
 sg13g2_tiehi _15994__1234 (.L_HI(net1234));
 sg13g2_tiehi _15993__1235 (.L_HI(net1235));
 sg13g2_tiehi _15992__1236 (.L_HI(net1236));
 sg13g2_tiehi _15991__1237 (.L_HI(net1237));
 sg13g2_tiehi _15990__1238 (.L_HI(net1238));
 sg13g2_tiehi _15961__1239 (.L_HI(net1239));
 sg13g2_tiehi _15960__1240 (.L_HI(net1240));
 sg13g2_tiehi _15959__1241 (.L_HI(net1241));
 sg13g2_tiehi _15958__1242 (.L_HI(net1242));
 sg13g2_tiehi _15957__1243 (.L_HI(net1243));
 sg13g2_tiehi _15928__1244 (.L_HI(net1244));
 sg13g2_tiehi _15927__1245 (.L_HI(net1245));
 sg13g2_tiehi _15926__1246 (.L_HI(net1246));
 sg13g2_tiehi _15925__1247 (.L_HI(net1247));
 sg13g2_tiehi _15924__1248 (.L_HI(net1248));
 sg13g2_tiehi _15923__1249 (.L_HI(net1249));
 sg13g2_tiehi _15922__1250 (.L_HI(net1250));
 sg13g2_tiehi _15921__1251 (.L_HI(net1251));
 sg13g2_tiehi _15920__1252 (.L_HI(net1252));
 sg13g2_tiehi _15919__1253 (.L_HI(net1253));
 sg13g2_tiehi _15918__1254 (.L_HI(net1254));
 sg13g2_tiehi _15917__1255 (.L_HI(net1255));
 sg13g2_tiehi _15916__1256 (.L_HI(net1256));
 sg13g2_tiehi _17049__1257 (.L_HI(net1257));
 sg13g2_tiehi _17048__1258 (.L_HI(net1258));
 sg13g2_tiehi _17047__1259 (.L_HI(net1259));
 sg13g2_tiehi _17046__1260 (.L_HI(net1260));
 sg13g2_tiehi _17045__1261 (.L_HI(net1261));
 sg13g2_tiehi _17044__1262 (.L_HI(net1262));
 sg13g2_tiehi _17043__1263 (.L_HI(net1263));
 sg13g2_tiehi _17042__1264 (.L_HI(net1264));
 sg13g2_tiehi _17330__1265 (.L_HI(net1265));
 sg13g2_tiehi _17041__1266 (.L_HI(net1266));
 sg13g2_tiehi _17252__1267 (.L_HI(net1267));
 sg13g2_tiehi _17040__1268 (.L_HI(net1268));
 sg13g2_tiehi _17039__1269 (.L_HI(net1269));
 sg13g2_tiehi _17038__1270 (.L_HI(net1270));
 sg13g2_tiehi _17037__1271 (.L_HI(net1271));
 sg13g2_tiehi _17036__1272 (.L_HI(net1272));
 sg13g2_tiehi _17035__1273 (.L_HI(net1273));
 sg13g2_tiehi _17034__1274 (.L_HI(net1274));
 sg13g2_tiehi _17033__1275 (.L_HI(net1275));
 sg13g2_tiehi _17032__1276 (.L_HI(net1276));
 sg13g2_tiehi _17031__1277 (.L_HI(net1277));
 sg13g2_tiehi _17030__1278 (.L_HI(net1278));
 sg13g2_tiehi _17029__1279 (.L_HI(net1279));
 sg13g2_tiehi _17028__1280 (.L_HI(net1280));
 sg13g2_tiehi _17027__1281 (.L_HI(net1281));
 sg13g2_tiehi _17026__1282 (.L_HI(net1282));
 sg13g2_tiehi _17025__1283 (.L_HI(net1283));
 sg13g2_tiehi _17024__1284 (.L_HI(net1284));
 sg13g2_tiehi _17023__1285 (.L_HI(net1285));
 sg13g2_tiehi _17022__1286 (.L_HI(net1286));
 sg13g2_tiehi _17021__1287 (.L_HI(net1287));
 sg13g2_tiehi _17020__1288 (.L_HI(net1288));
 sg13g2_tiehi _17019__1289 (.L_HI(net1289));
 sg13g2_tiehi _17018__1290 (.L_HI(net1290));
 sg13g2_tiehi _17017__1291 (.L_HI(net1291));
 sg13g2_tiehi _17016__1292 (.L_HI(net1292));
 sg13g2_tiehi _17015__1293 (.L_HI(net1293));
 sg13g2_tiehi _17014__1294 (.L_HI(net1294));
 sg13g2_tiehi _17013__1295 (.L_HI(net1295));
 sg13g2_tiehi _17012__1296 (.L_HI(net1296));
 sg13g2_tiehi _17011__1297 (.L_HI(net1297));
 sg13g2_tiehi _17010__1298 (.L_HI(net1298));
 sg13g2_tiehi _17009__1299 (.L_HI(net1299));
 sg13g2_tiehi _17008__1300 (.L_HI(net1300));
 sg13g2_tiehi _17007__1301 (.L_HI(net1301));
 sg13g2_tiehi _17006__1302 (.L_HI(net1302));
 sg13g2_tiehi _17005__1303 (.L_HI(net1303));
 sg13g2_tiehi _17004__1304 (.L_HI(net1304));
 sg13g2_tiehi _17003__1305 (.L_HI(net1305));
 sg13g2_tiehi _17002__1306 (.L_HI(net1306));
 sg13g2_tiehi _17001__1307 (.L_HI(net1307));
 sg13g2_tiehi _17000__1308 (.L_HI(net1308));
 sg13g2_tiehi _16999__1309 (.L_HI(net1309));
 sg13g2_tiehi _17296__1310 (.L_HI(net1310));
 sg13g2_tiehi _16998__1311 (.L_HI(net1311));
 sg13g2_tiehi _17251__1312 (.L_HI(net1312));
 sg13g2_tiehi _16997__1313 (.L_HI(net1313));
 sg13g2_tiehi _17322__1314 (.L_HI(net1314));
 sg13g2_tiehi _16996__1315 (.L_HI(net1315));
 sg13g2_tiehi _17250__1316 (.L_HI(net1316));
 sg13g2_tiehi _16995__1317 (.L_HI(net1317));
 sg13g2_tiehi _17295__1318 (.L_HI(net1318));
 sg13g2_tiehi _16994__1319 (.L_HI(net1319));
 sg13g2_tiehi _17249__1320 (.L_HI(net1320));
 sg13g2_tiehi _16993__1321 (.L_HI(net1321));
 sg13g2_tiehi _17329__1322 (.L_HI(net1322));
 sg13g2_tiehi _16992__1323 (.L_HI(net1323));
 sg13g2_tiehi _17248__1324 (.L_HI(net1324));
 sg13g2_tiehi _16991__1325 (.L_HI(net1325));
 sg13g2_tiehi _17294__1326 (.L_HI(net1326));
 sg13g2_tiehi _16990__1327 (.L_HI(net1327));
 sg13g2_tiehi _17247__1328 (.L_HI(net1328));
 sg13g2_tiehi _17074__1329 (.L_HI(net1329));
 sg13g2_tiehi _16989__1330 (.L_HI(net1330));
 sg13g2_tiehi _17321__1331 (.L_HI(net1331));
 sg13g2_tiehi _16988__1332 (.L_HI(net1332));
 sg13g2_tiehi _17246__1333 (.L_HI(net1333));
 sg13g2_tiehi _16987__1334 (.L_HI(net1334));
 sg13g2_tiehi _17293__1335 (.L_HI(net1335));
 sg13g2_tiehi _16986__1336 (.L_HI(net1336));
 sg13g2_tiehi _17245__1337 (.L_HI(net1337));
 sg13g2_tiehi _16985__1338 (.L_HI(net1338));
 sg13g2_tiehi _17320__1339 (.L_HI(net1339));
 sg13g2_tiehi _16984__1340 (.L_HI(net1340));
 sg13g2_tiehi _17244__1341 (.L_HI(net1341));
 sg13g2_tiehi _16983__1342 (.L_HI(net1342));
 sg13g2_tiehi _17292__1343 (.L_HI(net1343));
 sg13g2_tiehi _16982__1344 (.L_HI(net1344));
 sg13g2_tiehi _17243__1345 (.L_HI(net1345));
 sg13g2_tiehi _16981__1346 (.L_HI(net1346));
 sg13g2_tiehi _17291__1347 (.L_HI(net1347));
 sg13g2_tiehi _16980__1348 (.L_HI(net1348));
 sg13g2_tiehi _17242__1349 (.L_HI(net1349));
 sg13g2_tiehi _16979__1350 (.L_HI(net1350));
 sg13g2_tiehi _17290__1351 (.L_HI(net1351));
 sg13g2_tiehi _16978__1352 (.L_HI(net1352));
 sg13g2_tiehi _17241__1353 (.L_HI(net1353));
 sg13g2_tiehi _16977__1354 (.L_HI(net1354));
 sg13g2_tiehi _17289__1355 (.L_HI(net1355));
 sg13g2_tiehi _16976__1356 (.L_HI(net1356));
 sg13g2_tiehi _17240__1357 (.L_HI(net1357));
 sg13g2_tiehi _16975__1358 (.L_HI(net1358));
 sg13g2_tiehi _17319__1359 (.L_HI(net1359));
 sg13g2_tiehi _16974__1360 (.L_HI(net1360));
 sg13g2_tiehi _17239__1361 (.L_HI(net1361));
 sg13g2_tiehi _16973__1362 (.L_HI(net1362));
 sg13g2_tiehi _17288__1363 (.L_HI(net1363));
 sg13g2_tiehi _16972__1364 (.L_HI(net1364));
 sg13g2_tiehi _17238__1365 (.L_HI(net1365));
 sg13g2_tiehi _16971__1366 (.L_HI(net1366));
 sg13g2_tiehi _17318__1367 (.L_HI(net1367));
 sg13g2_tiehi _16970__1368 (.L_HI(net1368));
 sg13g2_tiehi _17237__1369 (.L_HI(net1369));
 sg13g2_tiehi _16969__1370 (.L_HI(net1370));
 sg13g2_tiehi _17287__1371 (.L_HI(net1371));
 sg13g2_tiehi _16968__1372 (.L_HI(net1372));
 sg13g2_tiehi _17236__1373 (.L_HI(net1373));
 sg13g2_tiehi _16967__1374 (.L_HI(net1374));
 sg13g2_tiehi _17317__1375 (.L_HI(net1375));
 sg13g2_tiehi _16966__1376 (.L_HI(net1376));
 sg13g2_tiehi _17235__1377 (.L_HI(net1377));
 sg13g2_tiehi _16965__1378 (.L_HI(net1378));
 sg13g2_tiehi _17286__1379 (.L_HI(net1379));
 sg13g2_tiehi _16964__1380 (.L_HI(net1380));
 sg13g2_tiehi _17234__1381 (.L_HI(net1381));
 sg13g2_tiehi _16963__1382 (.L_HI(net1382));
 sg13g2_tiehi _17316__1383 (.L_HI(net1383));
 sg13g2_tiehi _16962__1384 (.L_HI(net1384));
 sg13g2_tiehi _17233__1385 (.L_HI(net1385));
 sg13g2_tiehi _16961__1386 (.L_HI(net1386));
 sg13g2_tiehi _17285__1387 (.L_HI(net1387));
 sg13g2_tiehi _16960__1388 (.L_HI(net1388));
 sg13g2_tiehi _17232__1389 (.L_HI(net1389));
 sg13g2_tiehi _16959__1390 (.L_HI(net1390));
 sg13g2_tiehi _17315__1391 (.L_HI(net1391));
 sg13g2_tiehi _16958__1392 (.L_HI(net1392));
 sg13g2_tiehi _17231__1393 (.L_HI(net1393));
 sg13g2_tiehi _16957__1394 (.L_HI(net1394));
 sg13g2_tiehi _17284__1395 (.L_HI(net1395));
 sg13g2_tiehi _16956__1396 (.L_HI(net1396));
 sg13g2_tiehi _17230__1397 (.L_HI(net1397));
 sg13g2_tiehi _16955__1398 (.L_HI(net1398));
 sg13g2_tiehi _17314__1399 (.L_HI(net1399));
 sg13g2_tiehi _16954__1400 (.L_HI(net1400));
 sg13g2_tiehi _17229__1401 (.L_HI(net1401));
 sg13g2_tiehi _16953__1402 (.L_HI(net1402));
 sg13g2_tiehi _17283__1403 (.L_HI(net1403));
 sg13g2_tiehi _16952__1404 (.L_HI(net1404));
 sg13g2_tiehi _17228__1405 (.L_HI(net1405));
 sg13g2_tiehi _16951__1406 (.L_HI(net1406));
 sg13g2_tiehi _17313__1407 (.L_HI(net1407));
 sg13g2_tiehi _16950__1408 (.L_HI(net1408));
 sg13g2_tiehi _17227__1409 (.L_HI(net1409));
 sg13g2_tiehi _16949__1410 (.L_HI(net1410));
 sg13g2_tiehi _16948__1411 (.L_HI(net1411));
 sg13g2_tiehi _16947__1412 (.L_HI(net1412));
 sg13g2_tiehi _16946__1413 (.L_HI(net1413));
 sg13g2_tiehi _16945__1414 (.L_HI(net1414));
 sg13g2_tiehi _16944__1415 (.L_HI(net1415));
 sg13g2_tiehi _16943__1416 (.L_HI(net1416));
 sg13g2_tiehi _16942__1417 (.L_HI(net1417));
 sg13g2_tiehi _16941__1418 (.L_HI(net1418));
 sg13g2_tiehi _16940__1419 (.L_HI(net1419));
 sg13g2_tiehi _16939__1420 (.L_HI(net1420));
 sg13g2_tiehi _16938__1421 (.L_HI(net1421));
 sg13g2_tiehi _15915__1422 (.L_HI(net1422));
 sg13g2_tiehi _15929__1423 (.L_HI(net1423));
 sg13g2_tiehi _15930__1424 (.L_HI(net1424));
 sg13g2_tiehi _15931__1425 (.L_HI(net1425));
 sg13g2_tiehi _15932__1426 (.L_HI(net1426));
 sg13g2_tiehi _15933__1427 (.L_HI(net1427));
 sg13g2_tiehi _15934__1428 (.L_HI(net1428));
 sg13g2_tiehi _15935__1429 (.L_HI(net1429));
 sg13g2_tiehi _15936__1430 (.L_HI(net1430));
 sg13g2_tiehi _15937__1431 (.L_HI(net1431));
 sg13g2_tiehi _15938__1432 (.L_HI(net1432));
 sg13g2_tiehi _15939__1433 (.L_HI(net1433));
 sg13g2_inv_1 _08892__1 (.Y(net1434),
    .A(clknet_1_1__leaf_clk));
 sg13g2_buf_1 _18756_ (.A(net1),
    .X(uio_oe[0]));
 sg13g2_buf_1 _18757_ (.A(uio_oe[5]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _18758_ (.A(uio_oe[5]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _18759_ (.A(net1),
    .X(uio_oe[3]));
 sg13g2_buf_1 _18760_ (.A(uio_oe[5]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _18761_ (.A(net1),
    .X(uio_oe[6]));
 sg13g2_buf_1 _18762_ (.A(net1),
    .X(uio_oe[7]));
 sg13g2_buf_1 _18763_ (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .X(uio_out[0]));
 sg13g2_buf_1 _18764_ (.A(\i_tinyqv.mem.q_ctrl.spi_clk_out ),
    .X(uio_out[3]));
 sg13g2_buf_1 _18765_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .X(uio_out[6]));
 sg13g2_buf_1 _18766_ (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .X(uio_out[7]));
 sg13g2_buf_8 fanout1682 (.A(net1683),
    .X(net1682));
 sg13g2_buf_1 fanout1683 (.A(net1685),
    .X(net1683));
 sg13g2_buf_2 fanout1684 (.A(net1685),
    .X(net1684));
 sg13g2_buf_1 fanout1685 (.A(_04796_),
    .X(net1685));
 sg13g2_buf_8 fanout1686 (.A(net1689),
    .X(net1686));
 sg13g2_buf_8 fanout1687 (.A(net1689),
    .X(net1687));
 sg13g2_buf_1 fanout1688 (.A(net1689),
    .X(net1688));
 sg13g2_buf_8 fanout1689 (.A(_04754_),
    .X(net1689));
 sg13g2_buf_8 fanout1690 (.A(net1694),
    .X(net1690));
 sg13g2_buf_1 fanout1691 (.A(net1694),
    .X(net1691));
 sg13g2_buf_8 fanout1692 (.A(net1694),
    .X(net1692));
 sg13g2_buf_1 fanout1693 (.A(net1694),
    .X(net1693));
 sg13g2_buf_8 fanout1694 (.A(_04655_),
    .X(net1694));
 sg13g2_buf_8 fanout1695 (.A(net1696),
    .X(net1695));
 sg13g2_buf_8 fanout1696 (.A(net1698),
    .X(net1696));
 sg13g2_buf_2 fanout1697 (.A(net1698),
    .X(net1697));
 sg13g2_buf_1 fanout1698 (.A(_04654_),
    .X(net1698));
 sg13g2_buf_8 fanout1699 (.A(net1701),
    .X(net1699));
 sg13g2_buf_1 fanout1700 (.A(net1701),
    .X(net1700));
 sg13g2_buf_1 fanout1701 (.A(_04807_),
    .X(net1701));
 sg13g2_buf_2 fanout1702 (.A(_04716_),
    .X(net1702));
 sg13g2_buf_8 fanout1703 (.A(net1704),
    .X(net1703));
 sg13g2_buf_8 fanout1704 (.A(_04670_),
    .X(net1704));
 sg13g2_buf_8 fanout1705 (.A(_04669_),
    .X(net1705));
 sg13g2_buf_8 fanout1706 (.A(_04663_),
    .X(net1706));
 sg13g2_buf_8 fanout1707 (.A(net1709),
    .X(net1707));
 sg13g2_buf_1 fanout1708 (.A(net1709),
    .X(net1708));
 sg13g2_buf_1 fanout1709 (.A(_04629_),
    .X(net1709));
 sg13g2_buf_8 fanout1710 (.A(net1711),
    .X(net1710));
 sg13g2_buf_1 fanout1711 (.A(_04629_),
    .X(net1711));
 sg13g2_buf_8 fanout1712 (.A(net1714),
    .X(net1712));
 sg13g2_buf_1 fanout1713 (.A(net1714),
    .X(net1713));
 sg13g2_buf_2 fanout1714 (.A(_04629_),
    .X(net1714));
 sg13g2_buf_8 fanout1715 (.A(net1717),
    .X(net1715));
 sg13g2_buf_1 fanout1716 (.A(net1717),
    .X(net1716));
 sg13g2_buf_8 fanout1717 (.A(net1719),
    .X(net1717));
 sg13g2_buf_8 fanout1718 (.A(net1719),
    .X(net1718));
 sg13g2_buf_8 fanout1719 (.A(_04623_),
    .X(net1719));
 sg13g2_buf_8 fanout1720 (.A(_04622_),
    .X(net1720));
 sg13g2_buf_8 fanout1721 (.A(net1724),
    .X(net1721));
 sg13g2_buf_8 fanout1722 (.A(net1724),
    .X(net1722));
 sg13g2_buf_1 fanout1723 (.A(net1724),
    .X(net1723));
 sg13g2_buf_2 fanout1724 (.A(_04617_),
    .X(net1724));
 sg13g2_buf_8 fanout1725 (.A(_04618_),
    .X(net1725));
 sg13g2_buf_1 fanout1726 (.A(_04618_),
    .X(net1726));
 sg13g2_buf_8 fanout1727 (.A(net1729),
    .X(net1727));
 sg13g2_buf_8 fanout1728 (.A(net1729),
    .X(net1728));
 sg13g2_buf_8 fanout1729 (.A(_04462_),
    .X(net1729));
 sg13g2_buf_8 fanout1730 (.A(net1731),
    .X(net1730));
 sg13g2_buf_8 fanout1731 (.A(_05884_),
    .X(net1731));
 sg13g2_buf_8 fanout1732 (.A(net1733),
    .X(net1732));
 sg13g2_buf_8 fanout1733 (.A(_05284_),
    .X(net1733));
 sg13g2_buf_8 fanout1734 (.A(net1736),
    .X(net1734));
 sg13g2_buf_8 fanout1735 (.A(net1736),
    .X(net1735));
 sg13g2_buf_8 fanout1736 (.A(net1737),
    .X(net1736));
 sg13g2_buf_8 fanout1737 (.A(_06486_),
    .X(net1737));
 sg13g2_buf_8 fanout1738 (.A(net1740),
    .X(net1738));
 sg13g2_buf_8 fanout1739 (.A(net1740),
    .X(net1739));
 sg13g2_buf_8 fanout1740 (.A(net1741),
    .X(net1740));
 sg13g2_buf_8 fanout1741 (.A(_05889_),
    .X(net1741));
 sg13g2_buf_8 fanout1742 (.A(net1744),
    .X(net1742));
 sg13g2_buf_1 fanout1743 (.A(net1744),
    .X(net1743));
 sg13g2_buf_8 fanout1744 (.A(net1745),
    .X(net1744));
 sg13g2_buf_8 fanout1745 (.A(net1748),
    .X(net1745));
 sg13g2_buf_8 fanout1746 (.A(net1748),
    .X(net1746));
 sg13g2_buf_1 fanout1747 (.A(net1748),
    .X(net1747));
 sg13g2_buf_8 fanout1748 (.A(_05290_),
    .X(net1748));
 sg13g2_buf_8 fanout1749 (.A(net1750),
    .X(net1749));
 sg13g2_buf_8 fanout1750 (.A(net1751),
    .X(net1750));
 sg13g2_buf_1 fanout1751 (.A(_02807_),
    .X(net1751));
 sg13g2_buf_8 fanout1752 (.A(_02807_),
    .X(net1752));
 sg13g2_buf_8 fanout1753 (.A(_02806_),
    .X(net1753));
 sg13g2_buf_8 fanout1754 (.A(net1756),
    .X(net1754));
 sg13g2_buf_8 fanout1755 (.A(net1756),
    .X(net1755));
 sg13g2_buf_8 fanout1756 (.A(net1757),
    .X(net1756));
 sg13g2_buf_8 fanout1757 (.A(_02642_),
    .X(net1757));
 sg13g2_buf_8 fanout1758 (.A(net1759),
    .X(net1758));
 sg13g2_buf_8 fanout1759 (.A(_05281_),
    .X(net1759));
 sg13g2_buf_8 fanout1760 (.A(_05281_),
    .X(net1760));
 sg13g2_buf_8 fanout1761 (.A(net1763),
    .X(net1761));
 sg13g2_buf_8 fanout1762 (.A(net1763),
    .X(net1762));
 sg13g2_buf_8 fanout1763 (.A(_04676_),
    .X(net1763));
 sg13g2_buf_8 fanout1764 (.A(_04671_),
    .X(net1764));
 sg13g2_buf_1 fanout1765 (.A(_04671_),
    .X(net1765));
 sg13g2_buf_8 fanout1766 (.A(net1767),
    .X(net1766));
 sg13g2_buf_8 fanout1767 (.A(net1768),
    .X(net1767));
 sg13g2_buf_8 fanout1768 (.A(_06788_),
    .X(net1768));
 sg13g2_buf_8 fanout1769 (.A(net1770),
    .X(net1769));
 sg13g2_buf_8 fanout1770 (.A(net1772),
    .X(net1770));
 sg13g2_buf_8 fanout1771 (.A(net1772),
    .X(net1771));
 sg13g2_buf_8 fanout1772 (.A(_06787_),
    .X(net1772));
 sg13g2_buf_8 fanout1773 (.A(_04311_),
    .X(net1773));
 sg13g2_buf_8 fanout1774 (.A(_04310_),
    .X(net1774));
 sg13g2_buf_1 fanout1775 (.A(_04310_),
    .X(net1775));
 sg13g2_buf_8 fanout1776 (.A(_04310_),
    .X(net1776));
 sg13g2_buf_8 fanout1777 (.A(_03643_),
    .X(net1777));
 sg13g2_buf_8 fanout1778 (.A(net1779),
    .X(net1778));
 sg13g2_buf_8 fanout1779 (.A(_03641_),
    .X(net1779));
 sg13g2_buf_8 fanout1780 (.A(net1782),
    .X(net1780));
 sg13g2_buf_1 fanout1781 (.A(net1782),
    .X(net1781));
 sg13g2_buf_8 fanout1782 (.A(net1783),
    .X(net1782));
 sg13g2_buf_8 fanout1783 (.A(_06046_),
    .X(net1783));
 sg13g2_buf_8 fanout1784 (.A(net1785),
    .X(net1784));
 sg13g2_buf_8 fanout1785 (.A(net1792),
    .X(net1785));
 sg13g2_buf_8 fanout1786 (.A(net1788),
    .X(net1786));
 sg13g2_buf_1 fanout1787 (.A(net1788),
    .X(net1787));
 sg13g2_buf_1 fanout1788 (.A(net1789),
    .X(net1788));
 sg13g2_buf_1 fanout1789 (.A(net1790),
    .X(net1789));
 sg13g2_buf_2 fanout1790 (.A(net1792),
    .X(net1790));
 sg13g2_buf_8 fanout1791 (.A(net1792),
    .X(net1791));
 sg13g2_buf_2 fanout1792 (.A(net1793),
    .X(net1792));
 sg13g2_buf_8 fanout1793 (.A(_06045_),
    .X(net1793));
 sg13g2_buf_8 fanout1794 (.A(net1795),
    .X(net1794));
 sg13g2_buf_1 fanout1795 (.A(net1796),
    .X(net1795));
 sg13g2_buf_2 fanout1796 (.A(net1798),
    .X(net1796));
 sg13g2_buf_8 fanout1797 (.A(net1798),
    .X(net1797));
 sg13g2_buf_8 fanout1798 (.A(_03651_),
    .X(net1798));
 sg13g2_buf_8 fanout1799 (.A(_03637_),
    .X(net1799));
 sg13g2_buf_8 fanout1800 (.A(_03637_),
    .X(net1800));
 sg13g2_buf_8 fanout1801 (.A(_03634_),
    .X(net1801));
 sg13g2_buf_8 fanout1802 (.A(_03633_),
    .X(net1802));
 sg13g2_buf_1 fanout1803 (.A(_03633_),
    .X(net1803));
 sg13g2_buf_8 fanout1804 (.A(_03633_),
    .X(net1804));
 sg13g2_buf_8 fanout1805 (.A(_02751_),
    .X(net1805));
 sg13g2_buf_1 fanout1806 (.A(_02751_),
    .X(net1806));
 sg13g2_buf_8 fanout1807 (.A(net1809),
    .X(net1807));
 sg13g2_buf_2 fanout1808 (.A(net1809),
    .X(net1808));
 sg13g2_buf_8 fanout1809 (.A(_02557_),
    .X(net1809));
 sg13g2_buf_8 fanout1810 (.A(net1811),
    .X(net1810));
 sg13g2_buf_8 fanout1811 (.A(net1813),
    .X(net1811));
 sg13g2_buf_8 fanout1812 (.A(net1813),
    .X(net1812));
 sg13g2_buf_8 fanout1813 (.A(_02556_),
    .X(net1813));
 sg13g2_buf_8 fanout1814 (.A(net1815),
    .X(net1814));
 sg13g2_buf_8 fanout1815 (.A(_06044_),
    .X(net1815));
 sg13g2_buf_8 fanout1816 (.A(_06043_),
    .X(net1816));
 sg13g2_buf_1 fanout1817 (.A(net1818),
    .X(net1817));
 sg13g2_buf_8 fanout1818 (.A(_06043_),
    .X(net1818));
 sg13g2_buf_8 fanout1819 (.A(net1820),
    .X(net1819));
 sg13g2_buf_8 fanout1820 (.A(_03652_),
    .X(net1820));
 sg13g2_buf_8 fanout1821 (.A(_03652_),
    .X(net1821));
 sg13g2_buf_8 fanout1822 (.A(_03652_),
    .X(net1822));
 sg13g2_buf_8 fanout1823 (.A(net1824),
    .X(net1823));
 sg13g2_buf_8 fanout1824 (.A(_04314_),
    .X(net1824));
 sg13g2_buf_8 fanout1825 (.A(net1827),
    .X(net1825));
 sg13g2_buf_1 fanout1826 (.A(net1827),
    .X(net1826));
 sg13g2_buf_8 fanout1827 (.A(_04313_),
    .X(net1827));
 sg13g2_buf_2 fanout1828 (.A(net1829),
    .X(net1828));
 sg13g2_buf_8 fanout1829 (.A(net1830),
    .X(net1829));
 sg13g2_buf_8 fanout1830 (.A(net1833),
    .X(net1830));
 sg13g2_buf_8 fanout1831 (.A(net1832),
    .X(net1831));
 sg13g2_buf_8 fanout1832 (.A(net1833),
    .X(net1832));
 sg13g2_buf_2 fanout1833 (.A(net1834),
    .X(net1833));
 sg13g2_buf_2 fanout1834 (.A(_03531_),
    .X(net1834));
 sg13g2_buf_8 fanout1835 (.A(net1836),
    .X(net1835));
 sg13g2_buf_8 fanout1836 (.A(net1837),
    .X(net1836));
 sg13g2_buf_8 fanout1837 (.A(net1841),
    .X(net1837));
 sg13g2_buf_8 fanout1838 (.A(net1841),
    .X(net1838));
 sg13g2_buf_2 fanout1839 (.A(net1841),
    .X(net1839));
 sg13g2_buf_8 fanout1840 (.A(net1841),
    .X(net1840));
 sg13g2_buf_8 fanout1841 (.A(_03530_),
    .X(net1841));
 sg13g2_buf_8 fanout1842 (.A(net1843),
    .X(net1842));
 sg13g2_buf_8 fanout1843 (.A(net1844),
    .X(net1843));
 sg13g2_buf_1 fanout1844 (.A(net1846),
    .X(net1844));
 sg13g2_buf_8 fanout1845 (.A(net1846),
    .X(net1845));
 sg13g2_buf_8 fanout1846 (.A(_03529_),
    .X(net1846));
 sg13g2_buf_8 fanout1847 (.A(net1848),
    .X(net1847));
 sg13g2_buf_8 fanout1848 (.A(net1849),
    .X(net1848));
 sg13g2_buf_8 fanout1849 (.A(_03528_),
    .X(net1849));
 sg13g2_buf_8 fanout1850 (.A(net1852),
    .X(net1850));
 sg13g2_buf_1 fanout1851 (.A(net1852),
    .X(net1851));
 sg13g2_buf_8 fanout1852 (.A(_02479_),
    .X(net1852));
 sg13g2_buf_8 fanout1853 (.A(net1854),
    .X(net1853));
 sg13g2_buf_8 fanout1854 (.A(\debug_rd[3] ),
    .X(net1854));
 sg13g2_buf_8 fanout1855 (.A(_02489_),
    .X(net1855));
 sg13g2_buf_8 fanout1856 (.A(_02489_),
    .X(net1856));
 sg13g2_buf_8 fanout1857 (.A(net1858),
    .X(net1857));
 sg13g2_buf_1 fanout1858 (.A(net1859),
    .X(net1858));
 sg13g2_buf_8 fanout1859 (.A(net1860),
    .X(net1859));
 sg13g2_buf_8 fanout1860 (.A(_02488_),
    .X(net1860));
 sg13g2_buf_8 fanout1861 (.A(_02488_),
    .X(net1861));
 sg13g2_buf_2 fanout1862 (.A(_02488_),
    .X(net1862));
 sg13g2_buf_8 fanout1863 (.A(net1864),
    .X(net1863));
 sg13g2_buf_8 fanout1864 (.A(net1865),
    .X(net1864));
 sg13g2_buf_8 fanout1865 (.A(net1866),
    .X(net1865));
 sg13g2_buf_8 fanout1866 (.A(_03437_),
    .X(net1866));
 sg13g2_buf_8 fanout1867 (.A(\debug_rd[2] ),
    .X(net1867));
 sg13g2_buf_8 fanout1868 (.A(\debug_rd[2] ),
    .X(net1868));
 sg13g2_buf_8 fanout1869 (.A(net1870),
    .X(net1869));
 sg13g2_buf_8 fanout1870 (.A(net1871),
    .X(net1870));
 sg13g2_buf_8 fanout1871 (.A(_03436_),
    .X(net1871));
 sg13g2_buf_8 fanout1872 (.A(\debug_rd[1] ),
    .X(net1872));
 sg13g2_buf_8 fanout1873 (.A(\debug_rd[1] ),
    .X(net1873));
 sg13g2_buf_8 fanout1874 (.A(net1875),
    .X(net1874));
 sg13g2_buf_8 fanout1875 (.A(\debug_rd[0] ),
    .X(net1875));
 sg13g2_buf_8 fanout1876 (.A(net1877),
    .X(net1876));
 sg13g2_buf_8 fanout1877 (.A(_03623_),
    .X(net1877));
 sg13g2_buf_8 fanout1878 (.A(net1881),
    .X(net1878));
 sg13g2_buf_8 fanout1879 (.A(net1881),
    .X(net1879));
 sg13g2_buf_1 fanout1880 (.A(net1881),
    .X(net1880));
 sg13g2_buf_2 fanout1881 (.A(net1884),
    .X(net1881));
 sg13g2_buf_8 fanout1882 (.A(net1883),
    .X(net1882));
 sg13g2_buf_8 fanout1883 (.A(net1884),
    .X(net1883));
 sg13g2_buf_8 fanout1884 (.A(_03509_),
    .X(net1884));
 sg13g2_buf_8 fanout1885 (.A(net1887),
    .X(net1885));
 sg13g2_buf_1 fanout1886 (.A(net1887),
    .X(net1886));
 sg13g2_buf_2 fanout1887 (.A(net1888),
    .X(net1887));
 sg13g2_buf_8 fanout1888 (.A(net1890),
    .X(net1888));
 sg13g2_buf_8 fanout1889 (.A(net1890),
    .X(net1889));
 sg13g2_buf_8 fanout1890 (.A(_03495_),
    .X(net1890));
 sg13g2_buf_2 fanout1891 (.A(net1892),
    .X(net1891));
 sg13g2_buf_8 fanout1892 (.A(_02095_),
    .X(net1892));
 sg13g2_buf_8 fanout1893 (.A(_05488_),
    .X(net1893));
 sg13g2_buf_1 fanout1894 (.A(_05488_),
    .X(net1894));
 sg13g2_buf_8 fanout1895 (.A(net1896),
    .X(net1895));
 sg13g2_buf_8 fanout1896 (.A(_05356_),
    .X(net1896));
 sg13g2_buf_8 fanout1897 (.A(_03408_),
    .X(net1897));
 sg13g2_buf_8 fanout1898 (.A(_03408_),
    .X(net1898));
 sg13g2_buf_8 fanout1899 (.A(_06228_),
    .X(net1899));
 sg13g2_buf_8 fanout1900 (.A(_05380_),
    .X(net1900));
 sg13g2_buf_1 fanout1901 (.A(_05380_),
    .X(net1901));
 sg13g2_buf_8 fanout1902 (.A(net1903),
    .X(net1902));
 sg13g2_buf_8 fanout1903 (.A(_03407_),
    .X(net1903));
 sg13g2_buf_8 fanout1904 (.A(_03289_),
    .X(net1904));
 sg13g2_buf_1 fanout1905 (.A(_03289_),
    .X(net1905));
 sg13g2_buf_8 fanout1906 (.A(net1907),
    .X(net1906));
 sg13g2_buf_8 fanout1907 (.A(net1908),
    .X(net1907));
 sg13g2_buf_1 fanout1908 (.A(_03279_),
    .X(net1908));
 sg13g2_buf_8 fanout1909 (.A(net1910),
    .X(net1909));
 sg13g2_buf_1 fanout1910 (.A(net1911),
    .X(net1910));
 sg13g2_buf_8 fanout1911 (.A(_03266_),
    .X(net1911));
 sg13g2_buf_8 fanout1912 (.A(_03266_),
    .X(net1912));
 sg13g2_buf_8 fanout1913 (.A(net1914),
    .X(net1913));
 sg13g2_buf_2 fanout1914 (.A(_03423_),
    .X(net1914));
 sg13g2_buf_8 fanout1915 (.A(net1917),
    .X(net1915));
 sg13g2_buf_8 fanout1916 (.A(net1917),
    .X(net1916));
 sg13g2_buf_8 fanout1917 (.A(net1918),
    .X(net1917));
 sg13g2_buf_8 fanout1918 (.A(_03418_),
    .X(net1918));
 sg13g2_buf_8 fanout1919 (.A(net1921),
    .X(net1919));
 sg13g2_buf_8 fanout1920 (.A(net1921),
    .X(net1920));
 sg13g2_buf_2 fanout1921 (.A(_03284_),
    .X(net1921));
 sg13g2_buf_8 fanout1922 (.A(_03278_),
    .X(net1922));
 sg13g2_buf_8 fanout1923 (.A(_03278_),
    .X(net1923));
 sg13g2_buf_8 fanout1924 (.A(net1925),
    .X(net1924));
 sg13g2_buf_8 fanout1925 (.A(_03324_),
    .X(net1925));
 sg13g2_buf_8 fanout1926 (.A(net1927),
    .X(net1926));
 sg13g2_buf_8 fanout1927 (.A(_03183_),
    .X(net1927));
 sg13g2_buf_8 fanout1928 (.A(net1931),
    .X(net1928));
 sg13g2_buf_1 fanout1929 (.A(net1931),
    .X(net1929));
 sg13g2_buf_8 fanout1930 (.A(net1931),
    .X(net1930));
 sg13g2_buf_2 fanout1931 (.A(net1932),
    .X(net1931));
 sg13g2_buf_1 fanout1932 (.A(net1933),
    .X(net1932));
 sg13g2_buf_8 fanout1933 (.A(_03323_),
    .X(net1933));
 sg13g2_buf_8 fanout1934 (.A(net1935),
    .X(net1934));
 sg13g2_buf_2 fanout1935 (.A(net1936),
    .X(net1935));
 sg13g2_buf_8 fanout1936 (.A(net1937),
    .X(net1936));
 sg13g2_buf_8 fanout1937 (.A(net1938),
    .X(net1937));
 sg13g2_buf_1 fanout1938 (.A(net1939),
    .X(net1938));
 sg13g2_buf_8 fanout1939 (.A(_03182_),
    .X(net1939));
 sg13g2_buf_8 fanout1940 (.A(_06075_),
    .X(net1940));
 sg13g2_buf_8 fanout1941 (.A(net1942),
    .X(net1941));
 sg13g2_buf_8 fanout1942 (.A(net1943),
    .X(net1942));
 sg13g2_buf_8 fanout1943 (.A(_03158_),
    .X(net1943));
 sg13g2_buf_8 fanout1944 (.A(net1946),
    .X(net1944));
 sg13g2_buf_1 fanout1945 (.A(net1946),
    .X(net1945));
 sg13g2_buf_8 fanout1946 (.A(_03158_),
    .X(net1946));
 sg13g2_buf_8 fanout1947 (.A(_03157_),
    .X(net1947));
 sg13g2_buf_2 fanout1948 (.A(_03157_),
    .X(net1948));
 sg13g2_buf_8 fanout1949 (.A(net1950),
    .X(net1949));
 sg13g2_buf_8 fanout1950 (.A(_03157_),
    .X(net1950));
 sg13g2_buf_8 fanout1951 (.A(net1952),
    .X(net1951));
 sg13g2_buf_8 fanout1952 (.A(_02060_),
    .X(net1952));
 sg13g2_buf_8 fanout1953 (.A(net1954),
    .X(net1953));
 sg13g2_buf_8 fanout1954 (.A(_02046_),
    .X(net1954));
 sg13g2_buf_8 fanout1955 (.A(_06050_),
    .X(net1955));
 sg13g2_buf_8 fanout1956 (.A(net1957),
    .X(net1956));
 sg13g2_buf_8 fanout1957 (.A(_05658_),
    .X(net1957));
 sg13g2_buf_8 fanout1958 (.A(_01941_),
    .X(net1958));
 sg13g2_buf_8 fanout1959 (.A(net1961),
    .X(net1959));
 sg13g2_buf_1 fanout1960 (.A(net1961),
    .X(net1960));
 sg13g2_buf_2 fanout1961 (.A(net1964),
    .X(net1961));
 sg13g2_buf_8 fanout1962 (.A(net1963),
    .X(net1962));
 sg13g2_buf_8 fanout1963 (.A(net1964),
    .X(net1963));
 sg13g2_buf_8 fanout1964 (.A(_01440_),
    .X(net1964));
 sg13g2_buf_8 fanout1965 (.A(net1966),
    .X(net1965));
 sg13g2_buf_8 fanout1966 (.A(_06574_),
    .X(net1966));
 sg13g2_buf_8 fanout1967 (.A(net1968),
    .X(net1967));
 sg13g2_buf_8 fanout1968 (.A(_06559_),
    .X(net1968));
 sg13g2_buf_8 fanout1969 (.A(_06544_),
    .X(net1969));
 sg13g2_buf_8 fanout1970 (.A(_06521_),
    .X(net1970));
 sg13g2_buf_2 fanout1971 (.A(_06521_),
    .X(net1971));
 sg13g2_buf_8 fanout1972 (.A(_06049_),
    .X(net1972));
 sg13g2_buf_8 fanout1973 (.A(_06048_),
    .X(net1973));
 sg13g2_buf_8 fanout1974 (.A(_05952_),
    .X(net1974));
 sg13g2_buf_1 fanout1975 (.A(_05952_),
    .X(net1975));
 sg13g2_buf_8 fanout1976 (.A(net1977),
    .X(net1976));
 sg13g2_buf_2 fanout1977 (.A(_05945_),
    .X(net1977));
 sg13g2_buf_8 fanout1978 (.A(net1979),
    .X(net1978));
 sg13g2_buf_8 fanout1979 (.A(_05771_),
    .X(net1979));
 sg13g2_buf_8 fanout1980 (.A(net1985),
    .X(net1980));
 sg13g2_buf_8 fanout1981 (.A(net1982),
    .X(net1981));
 sg13g2_buf_8 fanout1982 (.A(net1983),
    .X(net1982));
 sg13g2_buf_8 fanout1983 (.A(net1984),
    .X(net1983));
 sg13g2_buf_8 fanout1984 (.A(net1985),
    .X(net1984));
 sg13g2_buf_8 fanout1985 (.A(_05532_),
    .X(net1985));
 sg13g2_buf_8 fanout1986 (.A(_05531_),
    .X(net1986));
 sg13g2_buf_8 fanout1987 (.A(net1989),
    .X(net1987));
 sg13g2_buf_8 fanout1988 (.A(net1989),
    .X(net1988));
 sg13g2_buf_8 fanout1989 (.A(_02918_),
    .X(net1989));
 sg13g2_buf_8 fanout1990 (.A(_02898_),
    .X(net1990));
 sg13g2_buf_1 fanout1991 (.A(_02898_),
    .X(net1991));
 sg13g2_buf_8 fanout1992 (.A(_02840_),
    .X(net1992));
 sg13g2_buf_8 fanout1993 (.A(_02728_),
    .X(net1993));
 sg13g2_buf_8 fanout1994 (.A(_02727_),
    .X(net1994));
 sg13g2_buf_1 fanout1995 (.A(_02727_),
    .X(net1995));
 sg13g2_buf_8 fanout1996 (.A(net1998),
    .X(net1996));
 sg13g2_buf_1 fanout1997 (.A(net1998),
    .X(net1997));
 sg13g2_buf_8 fanout1998 (.A(_01919_),
    .X(net1998));
 sg13g2_buf_8 fanout1999 (.A(net2000),
    .X(net1999));
 sg13g2_buf_8 fanout2000 (.A(_01459_),
    .X(net2000));
 sg13g2_buf_8 fanout2001 (.A(net2002),
    .X(net2001));
 sg13g2_buf_8 fanout2002 (.A(_01447_),
    .X(net2002));
 sg13g2_buf_8 fanout2003 (.A(net2004),
    .X(net2003));
 sg13g2_buf_8 fanout2004 (.A(_01438_),
    .X(net2004));
 sg13g2_buf_8 fanout2005 (.A(_06705_),
    .X(net2005));
 sg13g2_buf_8 fanout2006 (.A(_06519_),
    .X(net2006));
 sg13g2_buf_8 fanout2007 (.A(_05983_),
    .X(net2007));
 sg13g2_buf_8 fanout2008 (.A(_05975_),
    .X(net2008));
 sg13g2_buf_8 fanout2009 (.A(_05967_),
    .X(net2009));
 sg13g2_buf_8 fanout2010 (.A(_05959_),
    .X(net2010));
 sg13g2_buf_1 fanout2011 (.A(_05959_),
    .X(net2011));
 sg13g2_buf_8 fanout2012 (.A(_05929_),
    .X(net2012));
 sg13g2_buf_1 fanout2013 (.A(_05929_),
    .X(net2013));
 sg13g2_buf_8 fanout2014 (.A(_05524_),
    .X(net2014));
 sg13g2_buf_8 fanout2015 (.A(_05513_),
    .X(net2015));
 sg13g2_buf_8 fanout2016 (.A(_05513_),
    .X(net2016));
 sg13g2_buf_8 fanout2017 (.A(net2018),
    .X(net2017));
 sg13g2_buf_8 fanout2018 (.A(net2019),
    .X(net2018));
 sg13g2_buf_1 fanout2019 (.A(_05355_),
    .X(net2019));
 sg13g2_buf_8 fanout2020 (.A(net2021),
    .X(net2020));
 sg13g2_buf_8 fanout2021 (.A(net2023),
    .X(net2021));
 sg13g2_buf_8 fanout2022 (.A(net2023),
    .X(net2022));
 sg13g2_buf_8 fanout2023 (.A(net2028),
    .X(net2023));
 sg13g2_buf_8 fanout2024 (.A(net2025),
    .X(net2024));
 sg13g2_buf_8 fanout2025 (.A(net2028),
    .X(net2025));
 sg13g2_buf_8 fanout2026 (.A(net2027),
    .X(net2026));
 sg13g2_buf_8 fanout2027 (.A(net2028),
    .X(net2027));
 sg13g2_buf_8 fanout2028 (.A(_05248_),
    .X(net2028));
 sg13g2_buf_8 fanout2029 (.A(net2030),
    .X(net2029));
 sg13g2_buf_8 fanout2030 (.A(net2032),
    .X(net2030));
 sg13g2_buf_8 fanout2031 (.A(net2032),
    .X(net2031));
 sg13g2_buf_8 fanout2032 (.A(_05218_),
    .X(net2032));
 sg13g2_buf_8 fanout2033 (.A(net2034),
    .X(net2033));
 sg13g2_buf_8 fanout2034 (.A(net2037),
    .X(net2034));
 sg13g2_buf_8 fanout2035 (.A(net2036),
    .X(net2035));
 sg13g2_buf_8 fanout2036 (.A(net2037),
    .X(net2036));
 sg13g2_buf_8 fanout2037 (.A(_05218_),
    .X(net2037));
 sg13g2_buf_8 fanout2038 (.A(net2039),
    .X(net2038));
 sg13g2_buf_8 fanout2039 (.A(_05179_),
    .X(net2039));
 sg13g2_buf_8 fanout2040 (.A(net2049),
    .X(net2040));
 sg13g2_buf_2 fanout2041 (.A(net2049),
    .X(net2041));
 sg13g2_buf_8 fanout2042 (.A(net2045),
    .X(net2042));
 sg13g2_buf_1 fanout2043 (.A(net2045),
    .X(net2043));
 sg13g2_buf_8 fanout2044 (.A(net2045),
    .X(net2044));
 sg13g2_buf_8 fanout2045 (.A(net2049),
    .X(net2045));
 sg13g2_buf_8 fanout2046 (.A(net2049),
    .X(net2046));
 sg13g2_buf_1 fanout2047 (.A(net2048),
    .X(net2047));
 sg13g2_buf_8 fanout2048 (.A(net2049),
    .X(net2048));
 sg13g2_buf_8 fanout2049 (.A(_05178_),
    .X(net2049));
 sg13g2_buf_8 fanout2050 (.A(_03153_),
    .X(net2050));
 sg13g2_buf_8 fanout2051 (.A(_03153_),
    .X(net2051));
 sg13g2_buf_8 fanout2052 (.A(net2054),
    .X(net2052));
 sg13g2_buf_8 fanout2053 (.A(net2054),
    .X(net2053));
 sg13g2_buf_8 fanout2054 (.A(_03130_),
    .X(net2054));
 sg13g2_buf_8 fanout2055 (.A(_03126_),
    .X(net2055));
 sg13g2_buf_8 fanout2056 (.A(net2059),
    .X(net2056));
 sg13g2_buf_2 fanout2057 (.A(net2058),
    .X(net2057));
 sg13g2_buf_1 fanout2058 (.A(net2059),
    .X(net2058));
 sg13g2_buf_1 fanout2059 (.A(_02917_),
    .X(net2059));
 sg13g2_buf_8 fanout2060 (.A(net2061),
    .X(net2060));
 sg13g2_buf_8 fanout2061 (.A(net2063),
    .X(net2061));
 sg13g2_buf_8 fanout2062 (.A(net2063),
    .X(net2062));
 sg13g2_buf_8 fanout2063 (.A(_02808_),
    .X(net2063));
 sg13g2_buf_8 fanout2064 (.A(net2065),
    .X(net2064));
 sg13g2_buf_8 fanout2065 (.A(_02500_),
    .X(net2065));
 sg13g2_buf_8 fanout2066 (.A(_02500_),
    .X(net2066));
 sg13g2_buf_8 fanout2067 (.A(net2068),
    .X(net2067));
 sg13g2_buf_2 fanout2068 (.A(_02499_),
    .X(net2068));
 sg13g2_buf_2 fanout2069 (.A(net2070),
    .X(net2069));
 sg13g2_buf_2 fanout2070 (.A(net2071),
    .X(net2070));
 sg13g2_buf_1 fanout2071 (.A(_02499_),
    .X(net2071));
 sg13g2_buf_8 fanout2072 (.A(net2073),
    .X(net2072));
 sg13g2_buf_8 fanout2073 (.A(net2075),
    .X(net2073));
 sg13g2_buf_8 fanout2074 (.A(net2075),
    .X(net2074));
 sg13g2_buf_8 fanout2075 (.A(_06793_),
    .X(net2075));
 sg13g2_buf_8 fanout2076 (.A(net2077),
    .X(net2076));
 sg13g2_buf_8 fanout2077 (.A(net2080),
    .X(net2077));
 sg13g2_buf_8 fanout2078 (.A(net2079),
    .X(net2078));
 sg13g2_buf_8 fanout2079 (.A(net2080),
    .X(net2079));
 sg13g2_buf_8 fanout2080 (.A(_06793_),
    .X(net2080));
 sg13g2_buf_8 fanout2081 (.A(_05322_),
    .X(net2081));
 sg13g2_buf_8 fanout2082 (.A(net2084),
    .X(net2082));
 sg13g2_buf_2 fanout2083 (.A(net2084),
    .X(net2083));
 sg13g2_buf_8 fanout2084 (.A(_05312_),
    .X(net2084));
 sg13g2_buf_8 fanout2085 (.A(_05310_),
    .X(net2085));
 sg13g2_buf_1 fanout2086 (.A(_05310_),
    .X(net2086));
 sg13g2_buf_8 fanout2087 (.A(net2089),
    .X(net2087));
 sg13g2_buf_2 fanout2088 (.A(net2089),
    .X(net2088));
 sg13g2_buf_8 fanout2089 (.A(_05177_),
    .X(net2089));
 sg13g2_buf_8 fanout2090 (.A(_05176_),
    .X(net2090));
 sg13g2_buf_1 fanout2091 (.A(_05176_),
    .X(net2091));
 sg13g2_buf_8 fanout2092 (.A(net2095),
    .X(net2092));
 sg13g2_buf_8 fanout2093 (.A(net2094),
    .X(net2093));
 sg13g2_buf_8 fanout2094 (.A(net2095),
    .X(net2094));
 sg13g2_buf_8 fanout2095 (.A(_05176_),
    .X(net2095));
 sg13g2_buf_8 fanout2096 (.A(net2100),
    .X(net2096));
 sg13g2_buf_8 fanout2097 (.A(net2098),
    .X(net2097));
 sg13g2_buf_8 fanout2098 (.A(net2099),
    .X(net2098));
 sg13g2_buf_8 fanout2099 (.A(net2100),
    .X(net2099));
 sg13g2_buf_8 fanout2100 (.A(_03152_),
    .X(net2100));
 sg13g2_buf_8 fanout2101 (.A(net2102),
    .X(net2101));
 sg13g2_buf_8 fanout2102 (.A(_03149_),
    .X(net2102));
 sg13g2_buf_8 fanout2103 (.A(net2105),
    .X(net2103));
 sg13g2_buf_8 fanout2104 (.A(net2105),
    .X(net2104));
 sg13g2_buf_8 fanout2105 (.A(_03149_),
    .X(net2105));
 sg13g2_buf_8 fanout2106 (.A(net2108),
    .X(net2106));
 sg13g2_buf_1 fanout2107 (.A(net2108),
    .X(net2107));
 sg13g2_buf_8 fanout2108 (.A(net2109),
    .X(net2108));
 sg13g2_buf_8 fanout2109 (.A(_03129_),
    .X(net2109));
 sg13g2_buf_8 fanout2110 (.A(net2111),
    .X(net2110));
 sg13g2_buf_8 fanout2111 (.A(_03125_),
    .X(net2111));
 sg13g2_buf_8 fanout2112 (.A(net2114),
    .X(net2112));
 sg13g2_buf_8 fanout2113 (.A(_03125_),
    .X(net2113));
 sg13g2_buf_8 fanout2114 (.A(_03125_),
    .X(net2114));
 sg13g2_buf_8 fanout2115 (.A(_02896_),
    .X(net2115));
 sg13g2_buf_8 fanout2116 (.A(net2117),
    .X(net2116));
 sg13g2_buf_2 fanout2117 (.A(net2118),
    .X(net2117));
 sg13g2_buf_1 fanout2118 (.A(net2119),
    .X(net2118));
 sg13g2_buf_1 fanout2119 (.A(net2121),
    .X(net2119));
 sg13g2_buf_8 fanout2120 (.A(net2121),
    .X(net2120));
 sg13g2_buf_2 fanout2121 (.A(_02632_),
    .X(net2121));
 sg13g2_buf_8 fanout2122 (.A(_02632_),
    .X(net2122));
 sg13g2_buf_8 fanout2123 (.A(net2124),
    .X(net2123));
 sg13g2_buf_8 fanout2124 (.A(net2125),
    .X(net2124));
 sg13g2_buf_8 fanout2125 (.A(_02631_),
    .X(net2125));
 sg13g2_buf_8 fanout2126 (.A(net2127),
    .X(net2126));
 sg13g2_buf_8 fanout2127 (.A(net2128),
    .X(net2127));
 sg13g2_buf_8 fanout2128 (.A(_02553_),
    .X(net2128));
 sg13g2_buf_8 fanout2129 (.A(_02550_),
    .X(net2129));
 sg13g2_buf_8 fanout2130 (.A(_02547_),
    .X(net2130));
 sg13g2_buf_8 fanout2131 (.A(net2133),
    .X(net2131));
 sg13g2_buf_1 fanout2132 (.A(net2133),
    .X(net2132));
 sg13g2_buf_8 fanout2133 (.A(_02541_),
    .X(net2133));
 sg13g2_buf_8 fanout2134 (.A(net2135),
    .X(net2134));
 sg13g2_buf_8 fanout2135 (.A(_02540_),
    .X(net2135));
 sg13g2_buf_8 fanout2136 (.A(net2137),
    .X(net2136));
 sg13g2_buf_8 fanout2137 (.A(_02535_),
    .X(net2137));
 sg13g2_buf_8 fanout2138 (.A(_02534_),
    .X(net2138));
 sg13g2_buf_8 fanout2139 (.A(net2140),
    .X(net2139));
 sg13g2_buf_2 fanout2140 (.A(_02524_),
    .X(net2140));
 sg13g2_buf_8 fanout2141 (.A(_02523_),
    .X(net2141));
 sg13g2_buf_2 fanout2142 (.A(_02523_),
    .X(net2142));
 sg13g2_buf_8 fanout2143 (.A(net2144),
    .X(net2143));
 sg13g2_buf_8 fanout2144 (.A(_02497_),
    .X(net2144));
 sg13g2_buf_8 fanout2145 (.A(net2146),
    .X(net2145));
 sg13g2_buf_8 fanout2146 (.A(_02484_),
    .X(net2146));
 sg13g2_buf_8 fanout2147 (.A(_01754_),
    .X(net2147));
 sg13g2_buf_8 fanout2148 (.A(_07012_),
    .X(net2148));
 sg13g2_buf_1 fanout2149 (.A(_07012_),
    .X(net2149));
 sg13g2_buf_8 fanout2150 (.A(_06980_),
    .X(net2150));
 sg13g2_buf_1 fanout2151 (.A(_06980_),
    .X(net2151));
 sg13g2_buf_8 fanout2152 (.A(_06702_),
    .X(net2152));
 sg13g2_buf_8 fanout2153 (.A(net2157),
    .X(net2153));
 sg13g2_buf_8 fanout2154 (.A(net2157),
    .X(net2154));
 sg13g2_buf_8 fanout2155 (.A(net2156),
    .X(net2155));
 sg13g2_buf_8 fanout2156 (.A(net2157),
    .X(net2156));
 sg13g2_buf_8 fanout2157 (.A(_05912_),
    .X(net2157));
 sg13g2_buf_8 fanout2158 (.A(net2159),
    .X(net2158));
 sg13g2_buf_8 fanout2159 (.A(_05509_),
    .X(net2159));
 sg13g2_buf_8 fanout2160 (.A(net2163),
    .X(net2160));
 sg13g2_buf_8 fanout2161 (.A(net2162),
    .X(net2161));
 sg13g2_buf_8 fanout2162 (.A(net2163),
    .X(net2162));
 sg13g2_buf_8 fanout2163 (.A(net2165),
    .X(net2163));
 sg13g2_buf_8 fanout2164 (.A(net2165),
    .X(net2164));
 sg13g2_buf_8 fanout2165 (.A(_05307_),
    .X(net2165));
 sg13g2_buf_8 fanout2166 (.A(net2167),
    .X(net2166));
 sg13g2_buf_1 fanout2167 (.A(_05247_),
    .X(net2167));
 sg13g2_buf_8 fanout2168 (.A(net2171),
    .X(net2168));
 sg13g2_buf_8 fanout2169 (.A(net2170),
    .X(net2169));
 sg13g2_buf_8 fanout2170 (.A(net2171),
    .X(net2170));
 sg13g2_buf_8 fanout2171 (.A(net2172),
    .X(net2171));
 sg13g2_buf_8 fanout2172 (.A(_05247_),
    .X(net2172));
 sg13g2_buf_8 fanout2173 (.A(net2174),
    .X(net2173));
 sg13g2_buf_1 fanout2174 (.A(_05217_),
    .X(net2174));
 sg13g2_buf_8 fanout2175 (.A(net2178),
    .X(net2175));
 sg13g2_buf_8 fanout2176 (.A(net2177),
    .X(net2176));
 sg13g2_buf_8 fanout2177 (.A(net2178),
    .X(net2177));
 sg13g2_buf_8 fanout2178 (.A(net2179),
    .X(net2178));
 sg13g2_buf_8 fanout2179 (.A(_05217_),
    .X(net2179));
 sg13g2_buf_8 fanout2180 (.A(net2184),
    .X(net2180));
 sg13g2_buf_8 fanout2181 (.A(net2184),
    .X(net2181));
 sg13g2_buf_8 fanout2182 (.A(net2183),
    .X(net2182));
 sg13g2_buf_8 fanout2183 (.A(net2184),
    .X(net2183));
 sg13g2_buf_8 fanout2184 (.A(net2185),
    .X(net2184));
 sg13g2_buf_8 fanout2185 (.A(_02492_),
    .X(net2185));
 sg13g2_buf_8 fanout2186 (.A(_02485_),
    .X(net2186));
 sg13g2_buf_8 fanout2187 (.A(net2188),
    .X(net2187));
 sg13g2_buf_8 fanout2188 (.A(_06700_),
    .X(net2188));
 sg13g2_buf_8 fanout2189 (.A(net2190),
    .X(net2189));
 sg13g2_buf_8 fanout2190 (.A(net2194),
    .X(net2190));
 sg13g2_buf_8 fanout2191 (.A(net2194),
    .X(net2191));
 sg13g2_buf_1 fanout2192 (.A(net2194),
    .X(net2192));
 sg13g2_buf_8 fanout2193 (.A(net2194),
    .X(net2193));
 sg13g2_buf_8 fanout2194 (.A(_05534_),
    .X(net2194));
 sg13g2_buf_8 fanout2195 (.A(net2196),
    .X(net2195));
 sg13g2_buf_8 fanout2196 (.A(_05170_),
    .X(net2196));
 sg13g2_buf_8 fanout2197 (.A(net2198),
    .X(net2197));
 sg13g2_buf_8 fanout2198 (.A(_03109_),
    .X(net2198));
 sg13g2_buf_8 fanout2199 (.A(net2200),
    .X(net2199));
 sg13g2_buf_1 fanout2200 (.A(_03109_),
    .X(net2200));
 sg13g2_buf_8 fanout2201 (.A(_03109_),
    .X(net2201));
 sg13g2_buf_2 fanout2202 (.A(net2203),
    .X(net2202));
 sg13g2_buf_8 fanout2203 (.A(_02914_),
    .X(net2203));
 sg13g2_buf_8 fanout2204 (.A(_02913_),
    .X(net2204));
 sg13g2_buf_8 fanout2205 (.A(_02913_),
    .X(net2205));
 sg13g2_buf_8 fanout2206 (.A(net2209),
    .X(net2206));
 sg13g2_buf_8 fanout2207 (.A(net2209),
    .X(net2207));
 sg13g2_buf_1 fanout2208 (.A(net2209),
    .X(net2208));
 sg13g2_buf_8 fanout2209 (.A(net2210),
    .X(net2209));
 sg13g2_buf_8 fanout2210 (.A(_02913_),
    .X(net2210));
 sg13g2_buf_8 fanout2211 (.A(_02901_),
    .X(net2211));
 sg13g2_buf_8 fanout2212 (.A(_02900_),
    .X(net2212));
 sg13g2_buf_1 fanout2213 (.A(_02900_),
    .X(net2213));
 sg13g2_buf_8 fanout2214 (.A(net2216),
    .X(net2214));
 sg13g2_buf_8 fanout2215 (.A(net2216),
    .X(net2215));
 sg13g2_buf_8 fanout2216 (.A(_02495_),
    .X(net2216));
 sg13g2_buf_8 fanout2217 (.A(net2218),
    .X(net2217));
 sg13g2_buf_8 fanout2218 (.A(_02494_),
    .X(net2218));
 sg13g2_buf_8 fanout2219 (.A(net2220),
    .X(net2219));
 sg13g2_buf_8 fanout2220 (.A(net2221),
    .X(net2220));
 sg13g2_buf_8 fanout2221 (.A(net2222),
    .X(net2221));
 sg13g2_buf_8 fanout2222 (.A(net2223),
    .X(net2222));
 sg13g2_buf_8 fanout2223 (.A(_02486_),
    .X(net2223));
 sg13g2_buf_8 fanout2224 (.A(net2226),
    .X(net2224));
 sg13g2_buf_1 fanout2225 (.A(net2226),
    .X(net2225));
 sg13g2_buf_8 fanout2226 (.A(_01740_),
    .X(net2226));
 sg13g2_buf_8 fanout2227 (.A(_01739_),
    .X(net2227));
 sg13g2_buf_8 fanout2228 (.A(net2230),
    .X(net2228));
 sg13g2_buf_8 fanout2229 (.A(net2230),
    .X(net2229));
 sg13g2_buf_8 fanout2230 (.A(_01386_),
    .X(net2230));
 sg13g2_buf_8 fanout2231 (.A(net2232),
    .X(net2231));
 sg13g2_buf_8 fanout2232 (.A(_01385_),
    .X(net2232));
 sg13g2_buf_8 fanout2233 (.A(net2234),
    .X(net2233));
 sg13g2_buf_8 fanout2234 (.A(net2235),
    .X(net2234));
 sg13g2_buf_8 fanout2235 (.A(_01372_),
    .X(net2235));
 sg13g2_buf_8 fanout2236 (.A(net2237),
    .X(net2236));
 sg13g2_buf_8 fanout2237 (.A(_01371_),
    .X(net2237));
 sg13g2_buf_8 fanout2238 (.A(net2239),
    .X(net2238));
 sg13g2_buf_8 fanout2239 (.A(net2240),
    .X(net2239));
 sg13g2_buf_8 fanout2240 (.A(_01215_),
    .X(net2240));
 sg13g2_buf_8 fanout2241 (.A(net2242),
    .X(net2241));
 sg13g2_buf_8 fanout2242 (.A(_01208_),
    .X(net2242));
 sg13g2_buf_8 fanout2243 (.A(_01208_),
    .X(net2243));
 sg13g2_buf_8 fanout2244 (.A(_01206_),
    .X(net2244));
 sg13g2_buf_8 fanout2245 (.A(_01164_),
    .X(net2245));
 sg13g2_buf_8 fanout2246 (.A(net2247),
    .X(net2246));
 sg13g2_buf_8 fanout2247 (.A(net2254),
    .X(net2247));
 sg13g2_buf_8 fanout2248 (.A(net2254),
    .X(net2248));
 sg13g2_buf_1 fanout2249 (.A(net2254),
    .X(net2249));
 sg13g2_buf_8 fanout2250 (.A(net2253),
    .X(net2250));
 sg13g2_buf_1 fanout2251 (.A(net2253),
    .X(net2251));
 sg13g2_buf_8 fanout2252 (.A(net2253),
    .X(net2252));
 sg13g2_buf_8 fanout2253 (.A(net2254),
    .X(net2253));
 sg13g2_buf_8 fanout2254 (.A(_01098_),
    .X(net2254));
 sg13g2_buf_8 fanout2255 (.A(net2256),
    .X(net2255));
 sg13g2_buf_2 fanout2256 (.A(net2264),
    .X(net2256));
 sg13g2_buf_8 fanout2257 (.A(net2261),
    .X(net2257));
 sg13g2_buf_1 fanout2258 (.A(net2261),
    .X(net2258));
 sg13g2_buf_8 fanout2259 (.A(net2261),
    .X(net2259));
 sg13g2_buf_1 fanout2260 (.A(net2261),
    .X(net2260));
 sg13g2_buf_2 fanout2261 (.A(net2264),
    .X(net2261));
 sg13g2_buf_8 fanout2262 (.A(net2264),
    .X(net2262));
 sg13g2_buf_1 fanout2263 (.A(net2264),
    .X(net2263));
 sg13g2_buf_2 fanout2264 (.A(net2289),
    .X(net2264));
 sg13g2_buf_8 fanout2265 (.A(net2266),
    .X(net2265));
 sg13g2_buf_8 fanout2266 (.A(net2269),
    .X(net2266));
 sg13g2_buf_8 fanout2267 (.A(net2269),
    .X(net2267));
 sg13g2_buf_1 fanout2268 (.A(net2269),
    .X(net2268));
 sg13g2_buf_8 fanout2269 (.A(net2289),
    .X(net2269));
 sg13g2_buf_8 fanout2270 (.A(net2272),
    .X(net2270));
 sg13g2_buf_8 fanout2271 (.A(net2272),
    .X(net2271));
 sg13g2_buf_8 fanout2272 (.A(net2273),
    .X(net2272));
 sg13g2_buf_8 fanout2273 (.A(net2274),
    .X(net2273));
 sg13g2_buf_8 fanout2274 (.A(net2289),
    .X(net2274));
 sg13g2_buf_8 fanout2275 (.A(net2277),
    .X(net2275));
 sg13g2_buf_8 fanout2276 (.A(net2277),
    .X(net2276));
 sg13g2_buf_8 fanout2277 (.A(net2278),
    .X(net2277));
 sg13g2_buf_8 fanout2278 (.A(net2279),
    .X(net2278));
 sg13g2_buf_8 fanout2279 (.A(net2288),
    .X(net2279));
 sg13g2_buf_8 fanout2280 (.A(net2283),
    .X(net2280));
 sg13g2_buf_8 fanout2281 (.A(net2283),
    .X(net2281));
 sg13g2_buf_1 fanout2282 (.A(net2283),
    .X(net2282));
 sg13g2_buf_8 fanout2283 (.A(net2288),
    .X(net2283));
 sg13g2_buf_8 fanout2284 (.A(net2285),
    .X(net2284));
 sg13g2_buf_1 fanout2285 (.A(net2286),
    .X(net2285));
 sg13g2_buf_8 fanout2286 (.A(net2287),
    .X(net2286));
 sg13g2_buf_1 fanout2287 (.A(net2288),
    .X(net2287));
 sg13g2_buf_8 fanout2288 (.A(net2289),
    .X(net2288));
 sg13g2_buf_8 fanout2289 (.A(\i_debug_uart_tx.resetn ),
    .X(net2289));
 sg13g2_buf_8 fanout2290 (.A(net2291),
    .X(net2290));
 sg13g2_buf_2 fanout2291 (.A(net2292),
    .X(net2291));
 sg13g2_buf_1 fanout2292 (.A(_06699_),
    .X(net2292));
 sg13g2_buf_8 fanout2293 (.A(_06698_),
    .X(net2293));
 sg13g2_buf_8 fanout2294 (.A(_06698_),
    .X(net2294));
 sg13g2_buf_8 fanout2295 (.A(net2297),
    .X(net2295));
 sg13g2_buf_1 fanout2296 (.A(net2297),
    .X(net2296));
 sg13g2_buf_8 fanout2297 (.A(net2298),
    .X(net2297));
 sg13g2_buf_8 fanout2298 (.A(_02003_),
    .X(net2298));
 sg13g2_buf_8 fanout2299 (.A(_01911_),
    .X(net2299));
 sg13g2_buf_8 fanout2300 (.A(_01905_),
    .X(net2300));
 sg13g2_buf_1 fanout2301 (.A(_01905_),
    .X(net2301));
 sg13g2_buf_8 fanout2302 (.A(_01904_),
    .X(net2302));
 sg13g2_buf_8 fanout2303 (.A(_01404_),
    .X(net2303));
 sg13g2_buf_8 fanout2304 (.A(net2305),
    .X(net2304));
 sg13g2_buf_8 fanout2305 (.A(_01216_),
    .X(net2305));
 sg13g2_buf_8 fanout2306 (.A(_01216_),
    .X(net2306));
 sg13g2_buf_8 fanout2307 (.A(_01202_),
    .X(net2307));
 sg13g2_buf_8 fanout2308 (.A(net2309),
    .X(net2308));
 sg13g2_buf_8 fanout2309 (.A(net2312),
    .X(net2309));
 sg13g2_buf_8 fanout2310 (.A(net2312),
    .X(net2310));
 sg13g2_buf_1 fanout2311 (.A(net2312),
    .X(net2311));
 sg13g2_buf_8 fanout2312 (.A(_01201_),
    .X(net2312));
 sg13g2_buf_8 fanout2313 (.A(net2315),
    .X(net2313));
 sg13g2_buf_8 fanout2314 (.A(net2315),
    .X(net2314));
 sg13g2_buf_8 fanout2315 (.A(net2316),
    .X(net2315));
 sg13g2_buf_8 fanout2316 (.A(_01198_),
    .X(net2316));
 sg13g2_buf_8 fanout2317 (.A(_01197_),
    .X(net2317));
 sg13g2_buf_8 fanout2318 (.A(net2319),
    .X(net2318));
 sg13g2_buf_8 fanout2319 (.A(net2321),
    .X(net2319));
 sg13g2_buf_8 fanout2320 (.A(net2321),
    .X(net2320));
 sg13g2_buf_8 fanout2321 (.A(net2322),
    .X(net2321));
 sg13g2_buf_8 fanout2322 (.A(_01196_),
    .X(net2322));
 sg13g2_buf_8 fanout2323 (.A(_01195_),
    .X(net2323));
 sg13g2_buf_8 fanout2324 (.A(_01163_),
    .X(net2324));
 sg13g2_buf_8 fanout2325 (.A(net2326),
    .X(net2325));
 sg13g2_buf_8 fanout2326 (.A(net2328),
    .X(net2326));
 sg13g2_buf_8 fanout2327 (.A(net2328),
    .X(net2327));
 sg13g2_buf_8 fanout2328 (.A(_01162_),
    .X(net2328));
 sg13g2_buf_8 fanout2329 (.A(_01140_),
    .X(net2329));
 sg13g2_buf_8 fanout2330 (.A(_01128_),
    .X(net2330));
 sg13g2_buf_8 fanout2331 (.A(net2332),
    .X(net2331));
 sg13g2_buf_1 fanout2332 (.A(net2333),
    .X(net2332));
 sg13g2_buf_2 fanout2333 (.A(net2334),
    .X(net2333));
 sg13g2_buf_8 fanout2334 (.A(_01121_),
    .X(net2334));
 sg13g2_buf_8 fanout2335 (.A(_01078_),
    .X(net2335));
 sg13g2_buf_8 fanout2336 (.A(net2337),
    .X(net2336));
 sg13g2_buf_8 fanout2337 (.A(_01067_),
    .X(net2337));
 sg13g2_buf_1 fanout2338 (.A(_01067_),
    .X(net2338));
 sg13g2_buf_8 fanout2339 (.A(net2340),
    .X(net2339));
 sg13g2_buf_8 fanout2340 (.A(net2349),
    .X(net2340));
 sg13g2_buf_8 fanout2341 (.A(net2349),
    .X(net2341));
 sg13g2_buf_1 fanout2342 (.A(net2349),
    .X(net2342));
 sg13g2_buf_8 fanout2343 (.A(net2345),
    .X(net2343));
 sg13g2_buf_1 fanout2344 (.A(net2345),
    .X(net2344));
 sg13g2_buf_8 fanout2345 (.A(net2346),
    .X(net2345));
 sg13g2_buf_8 fanout2346 (.A(net2347),
    .X(net2346));
 sg13g2_buf_8 fanout2347 (.A(net2348),
    .X(net2347));
 sg13g2_buf_8 fanout2348 (.A(net2349),
    .X(net2348));
 sg13g2_buf_8 fanout2349 (.A(_01065_),
    .X(net2349));
 sg13g2_buf_8 fanout2350 (.A(_00983_),
    .X(net2350));
 sg13g2_buf_8 fanout2351 (.A(_00974_),
    .X(net2351));
 sg13g2_buf_8 fanout2352 (.A(_00969_),
    .X(net2352));
 sg13g2_buf_8 fanout2353 (.A(net2354),
    .X(net2353));
 sg13g2_buf_8 fanout2354 (.A(_00924_),
    .X(net2354));
 sg13g2_buf_8 fanout2355 (.A(net2356),
    .X(net2355));
 sg13g2_buf_8 fanout2356 (.A(debug_instr_valid),
    .X(net2356));
 sg13g2_buf_8 fanout2357 (.A(net2358),
    .X(net2357));
 sg13g2_buf_8 fanout2358 (.A(net4155),
    .X(net2358));
 sg13g2_buf_8 fanout2359 (.A(net4090),
    .X(net2359));
 sg13g2_buf_8 fanout2360 (.A(net4096),
    .X(net2360));
 sg13g2_buf_8 fanout2361 (.A(net4109),
    .X(net2361));
 sg13g2_buf_8 fanout2362 (.A(net2365),
    .X(net2362));
 sg13g2_buf_8 fanout2363 (.A(net2365),
    .X(net2363));
 sg13g2_buf_2 fanout2364 (.A(net2365),
    .X(net2364));
 sg13g2_buf_8 fanout2365 (.A(net2366),
    .X(net2365));
 sg13g2_buf_8 fanout2366 (.A(net2367),
    .X(net2366));
 sg13g2_buf_8 fanout2367 (.A(net2370),
    .X(net2367));
 sg13g2_buf_8 fanout2368 (.A(net2369),
    .X(net2368));
 sg13g2_buf_8 fanout2369 (.A(net2370),
    .X(net2369));
 sg13g2_buf_8 fanout2370 (.A(net4163),
    .X(net2370));
 sg13g2_buf_8 fanout2371 (.A(net2372),
    .X(net2371));
 sg13g2_buf_8 fanout2372 (.A(net4121),
    .X(net2372));
 sg13g2_buf_8 fanout2373 (.A(net3926),
    .X(net2373));
 sg13g2_buf_1 fanout2374 (.A(\i_tinyqv.cpu.alu_op[0] ),
    .X(net2374));
 sg13g2_buf_8 fanout2375 (.A(net2378),
    .X(net2375));
 sg13g2_buf_8 fanout2376 (.A(net2378),
    .X(net2376));
 sg13g2_buf_8 fanout2377 (.A(net2378),
    .X(net2377));
 sg13g2_buf_8 fanout2378 (.A(net3681),
    .X(net2378));
 sg13g2_buf_8 fanout2379 (.A(net2380),
    .X(net2379));
 sg13g2_buf_8 fanout2380 (.A(net2381),
    .X(net2380));
 sg13g2_buf_8 fanout2381 (.A(\i_tinyqv.cpu.counter[3] ),
    .X(net2381));
 sg13g2_buf_8 fanout2382 (.A(net2383),
    .X(net2382));
 sg13g2_buf_8 fanout2383 (.A(net2384),
    .X(net2383));
 sg13g2_buf_8 fanout2384 (.A(net3595),
    .X(net2384));
 sg13g2_buf_8 fanout2385 (.A(net4135),
    .X(net2385));
 sg13g2_buf_8 fanout2386 (.A(\addr[3] ),
    .X(net2386));
 sg13g2_buf_8 fanout2387 (.A(\addr[2] ),
    .X(net2387));
 sg13g2_buf_8 fanout2388 (.A(net4066),
    .X(net2388));
 sg13g2_buf_8 fanout2389 (.A(net2390),
    .X(net2389));
 sg13g2_buf_8 fanout2390 (.A(net4098),
    .X(net2390));
 sg13g2_buf_8 fanout2391 (.A(net2392),
    .X(net2391));
 sg13g2_buf_8 fanout2392 (.A(net4140),
    .X(net2392));
 sg13g2_buf_8 fanout2393 (.A(net2394),
    .X(net2393));
 sg13g2_buf_8 fanout2394 (.A(net4102),
    .X(net2394));
 sg13g2_buf_8 fanout2395 (.A(net2396),
    .X(net2395));
 sg13g2_buf_8 fanout2396 (.A(net4148),
    .X(net2396));
 sg13g2_buf_8 fanout2397 (.A(net2398),
    .X(net2397));
 sg13g2_buf_8 fanout2398 (.A(net4128),
    .X(net2398));
 sg13g2_buf_8 fanout2399 (.A(net4157),
    .X(net2399));
 sg13g2_buf_8 fanout2400 (.A(net2402),
    .X(net2400));
 sg13g2_buf_1 fanout2401 (.A(net2402),
    .X(net2401));
 sg13g2_buf_1 fanout2402 (.A(net2403),
    .X(net2402));
 sg13g2_buf_1 fanout2403 (.A(net2408),
    .X(net2403));
 sg13g2_buf_8 fanout2404 (.A(net2408),
    .X(net2404));
 sg13g2_buf_1 fanout2405 (.A(net2408),
    .X(net2405));
 sg13g2_buf_8 fanout2406 (.A(net2407),
    .X(net2406));
 sg13g2_buf_8 fanout2407 (.A(net2408),
    .X(net2407));
 sg13g2_buf_8 fanout2408 (.A(\i_tinyqv.cpu.was_early_branch ),
    .X(net2408));
 sg13g2_buf_8 fanout2409 (.A(net4145),
    .X(net2409));
 sg13g2_buf_8 fanout2410 (.A(net4138),
    .X(net2410));
 sg13g2_buf_8 fanout2411 (.A(net4110),
    .X(net2411));
 sg13g2_buf_8 fanout2412 (.A(net4064),
    .X(net2412));
 sg13g2_buf_8 fanout2413 (.A(net4136),
    .X(net2413));
 sg13g2_buf_8 fanout2414 (.A(net4147),
    .X(net2414));
 sg13g2_buf_8 fanout2415 (.A(net4143),
    .X(net2415));
 sg13g2_buf_8 fanout2416 (.A(net4101),
    .X(net2416));
 sg13g2_buf_8 fanout2417 (.A(net4111),
    .X(net2417));
 sg13g2_buf_8 fanout2418 (.A(net4149),
    .X(net2418));
 sg13g2_buf_8 fanout2419 (.A(net4112),
    .X(net2419));
 sg13g2_buf_8 fanout2420 (.A(net2421),
    .X(net2420));
 sg13g2_buf_8 fanout2421 (.A(net4076),
    .X(net2421));
 sg13g2_buf_8 fanout2422 (.A(net4073),
    .X(net2422));
 sg13g2_buf_1 fanout2423 (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .X(net2423));
 sg13g2_buf_8 fanout2424 (.A(net4093),
    .X(net2424));
 sg13g2_buf_2 fanout2425 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(net2425));
 sg13g2_buf_8 fanout2426 (.A(net3279),
    .X(net2426));
 sg13g2_buf_8 fanout2427 (.A(net4125),
    .X(net2427));
 sg13g2_buf_8 fanout2428 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .X(net2428));
 sg13g2_buf_8 fanout2429 (.A(net2434),
    .X(net2429));
 sg13g2_buf_8 fanout2430 (.A(net2433),
    .X(net2430));
 sg13g2_buf_8 fanout2431 (.A(net2433),
    .X(net2431));
 sg13g2_buf_2 fanout2432 (.A(net2433),
    .X(net2432));
 sg13g2_buf_8 fanout2433 (.A(net2434),
    .X(net2433));
 sg13g2_buf_8 fanout2434 (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .X(net2434));
 sg13g2_buf_8 fanout2435 (.A(\i_tinyqv.mem.q_ctrl.data_ready ),
    .X(net2435));
 sg13g2_buf_8 fanout2436 (.A(net2437),
    .X(net2436));
 sg13g2_buf_8 fanout2437 (.A(net4071),
    .X(net2437));
 sg13g2_buf_8 fanout2438 (.A(net4114),
    .X(net2438));
 sg13g2_buf_8 fanout2439 (.A(net4132),
    .X(net2439));
 sg13g2_buf_8 fanout2440 (.A(net2444),
    .X(net2440));
 sg13g2_buf_8 fanout2441 (.A(net2443),
    .X(net2441));
 sg13g2_buf_8 fanout2442 (.A(net2443),
    .X(net2442));
 sg13g2_buf_8 fanout2443 (.A(net2444),
    .X(net2443));
 sg13g2_buf_2 fanout2444 (.A(net4160),
    .X(net2444));
 sg13g2_buf_8 fanout2445 (.A(net2447),
    .X(net2445));
 sg13g2_buf_1 fanout2446 (.A(net2447),
    .X(net2446));
 sg13g2_buf_2 fanout2447 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[23] ),
    .X(net2447));
 sg13g2_buf_2 fanout2448 (.A(net2449),
    .X(net2448));
 sg13g2_buf_2 fanout2449 (.A(net2451),
    .X(net2449));
 sg13g2_buf_8 fanout2450 (.A(net2451),
    .X(net2450));
 sg13g2_buf_8 fanout2451 (.A(net4162),
    .X(net2451));
 sg13g2_buf_8 fanout2452 (.A(net3638),
    .X(net2452));
 sg13g2_buf_8 fanout2453 (.A(net3615),
    .X(net2453));
 sg13g2_buf_8 fanout2454 (.A(net3686),
    .X(net2454));
 sg13g2_buf_8 fanout2455 (.A(net3538),
    .X(net2455));
 sg13g2_buf_8 fanout2456 (.A(net3645),
    .X(net2456));
 sg13g2_buf_8 fanout2457 (.A(net3918),
    .X(net2457));
 sg13g2_buf_8 fanout2458 (.A(net4126),
    .X(net2458));
 sg13g2_buf_8 fanout2459 (.A(net4133),
    .X(net2459));
 sg13g2_buf_8 fanout2460 (.A(net3719),
    .X(net2460));
 sg13g2_buf_8 fanout2461 (.A(net2462),
    .X(net2461));
 sg13g2_buf_8 fanout2462 (.A(net4151),
    .X(net2462));
 sg13g2_buf_8 fanout2463 (.A(net4104),
    .X(net2463));
 sg13g2_buf_8 fanout2464 (.A(net3540),
    .X(net2464));
 sg13g2_buf_8 fanout2465 (.A(\i_tinyqv.cpu.i_core.i_shift.a[1] ),
    .X(net2465));
 sg13g2_buf_8 fanout2466 (.A(\i_tinyqv.cpu.i_core.i_shift.a[0] ),
    .X(net2466));
 sg13g2_buf_8 fanout2467 (.A(net2468),
    .X(net2467));
 sg13g2_buf_8 fanout2468 (.A(net2471),
    .X(net2468));
 sg13g2_buf_8 fanout2469 (.A(net2470),
    .X(net2469));
 sg13g2_buf_8 fanout2470 (.A(net2471),
    .X(net2470));
 sg13g2_buf_2 fanout2471 (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[1] ),
    .X(net2471));
 sg13g2_buf_8 fanout2472 (.A(net2473),
    .X(net2472));
 sg13g2_buf_8 fanout2473 (.A(net2474),
    .X(net2473));
 sg13g2_buf_2 fanout2474 (.A(net2476),
    .X(net2474));
 sg13g2_buf_8 fanout2475 (.A(net2476),
    .X(net2475));
 sg13g2_buf_8 fanout2476 (.A(net2480),
    .X(net2476));
 sg13g2_buf_8 fanout2477 (.A(net2479),
    .X(net2477));
 sg13g2_buf_1 fanout2478 (.A(net2479),
    .X(net2478));
 sg13g2_buf_8 fanout2479 (.A(net2480),
    .X(net2479));
 sg13g2_buf_8 fanout2480 (.A(net4159),
    .X(net2480));
 sg13g2_buf_8 fanout2481 (.A(net4023),
    .X(net2481));
 sg13g2_buf_8 fanout2482 (.A(net2483),
    .X(net2482));
 sg13g2_buf_8 fanout2483 (.A(net2485),
    .X(net2483));
 sg13g2_buf_8 fanout2484 (.A(net2485),
    .X(net2484));
 sg13g2_buf_8 fanout2485 (.A(net2499),
    .X(net2485));
 sg13g2_buf_8 fanout2486 (.A(net2488),
    .X(net2486));
 sg13g2_buf_1 fanout2487 (.A(net2488),
    .X(net2487));
 sg13g2_buf_8 fanout2488 (.A(net2499),
    .X(net2488));
 sg13g2_buf_8 fanout2489 (.A(net2491),
    .X(net2489));
 sg13g2_buf_8 fanout2490 (.A(net2491),
    .X(net2490));
 sg13g2_buf_8 fanout2491 (.A(net2499),
    .X(net2491));
 sg13g2_buf_8 fanout2492 (.A(net2493),
    .X(net2492));
 sg13g2_buf_8 fanout2493 (.A(net2494),
    .X(net2493));
 sg13g2_buf_8 fanout2494 (.A(net2499),
    .X(net2494));
 sg13g2_buf_8 fanout2495 (.A(net2496),
    .X(net2495));
 sg13g2_buf_8 fanout2496 (.A(net2497),
    .X(net2496));
 sg13g2_buf_8 fanout2497 (.A(net2498),
    .X(net2497));
 sg13g2_buf_8 fanout2498 (.A(net2499),
    .X(net2498));
 sg13g2_buf_8 fanout2499 (.A(net3628),
    .X(net2499));
 sg13g2_buf_8 fanout2500 (.A(net4117),
    .X(net2500));
 sg13g2_buf_8 fanout2501 (.A(net4113),
    .X(net2501));
 sg13g2_buf_8 fanout2502 (.A(net4129),
    .X(net2502));
 sg13g2_buf_8 fanout2503 (.A(net4127),
    .X(net2503));
 sg13g2_buf_8 fanout2504 (.A(net4127),
    .X(net2504));
 sg13g2_buf_8 fanout2505 (.A(net2506),
    .X(net2505));
 sg13g2_buf_8 fanout2506 (.A(net5),
    .X(net2506));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_tiehi _15940__14 (.L_HI(net14));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(delaynet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_buf_8 clkbuf_leaf_0_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_0_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_1_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_1_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_2_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_2_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_3_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_3_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_4_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_4_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_5_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_5_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_6_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_6_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_7_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_7_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_8_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_8_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_9_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_9_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_10_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_10_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_11_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_11_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_12_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_12_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_13_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_13_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_14_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_14_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_15_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_15_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_16_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_16_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_17_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_17_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_18_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_18_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_19_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_19_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_20_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_20_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_21_clk_regs (.A(clknet_5_3__leaf_clk_regs),
    .X(clknet_leaf_21_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_22_clk_regs (.A(clknet_5_2__leaf_clk_regs),
    .X(clknet_leaf_22_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_23_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_23_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_24_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_24_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_25_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_25_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_26_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_26_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_27_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_27_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_28_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_28_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_29_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_29_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_30_clk_regs (.A(clknet_5_9__leaf_clk_regs),
    .X(clknet_leaf_30_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_31_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_31_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_32_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_32_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_33_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_33_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_34_clk_regs (.A(clknet_5_8__leaf_clk_regs),
    .X(clknet_leaf_34_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_35_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_35_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_36_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_36_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_37_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_37_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_38_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_38_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_39_clk_regs (.A(clknet_5_10__leaf_clk_regs),
    .X(clknet_leaf_39_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_40_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_40_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_41_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_41_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_42_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_42_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_43_clk_regs (.A(clknet_5_11__leaf_clk_regs),
    .X(clknet_leaf_43_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_44_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_44_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_45_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_45_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_46_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_46_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_47_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_47_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_48_clk_regs (.A(clknet_5_14__leaf_clk_regs),
    .X(clknet_leaf_48_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_49_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_49_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_50_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_50_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_51_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_51_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_52_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_52_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_53_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_53_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_54_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_54_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_55_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_55_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_56_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_56_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_57_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_57_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_58_clk_regs (.A(clknet_5_15__leaf_clk_regs),
    .X(clknet_leaf_58_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_59_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_59_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_60_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_60_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_61_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_61_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_62_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_62_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_63_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_63_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_64_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_64_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_65_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_65_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_66_clk_regs (.A(clknet_5_13__leaf_clk_regs),
    .X(clknet_leaf_66_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_67_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_67_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_68_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_68_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_69_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_69_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_70_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_70_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_71_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_71_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_72_clk_regs (.A(clknet_5_12__leaf_clk_regs),
    .X(clknet_leaf_72_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_73_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_73_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_74_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_74_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_75_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_75_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_76_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_76_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_77_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_77_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_78_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_78_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_79_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_79_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_80_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_80_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_81_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_81_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_82_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_82_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_83_clk_regs (.A(clknet_5_30__leaf_clk_regs),
    .X(clknet_leaf_83_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_84_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_84_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_85_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_85_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_86_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_86_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_87_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_87_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_88_clk_regs (.A(clknet_5_31__leaf_clk_regs),
    .X(clknet_leaf_88_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_89_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_89_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_90_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_90_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_91_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_91_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_92_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_92_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_93_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_93_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_94_clk_regs (.A(clknet_5_26__leaf_clk_regs),
    .X(clknet_leaf_94_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_95_clk_regs (.A(clknet_5_27__leaf_clk_regs),
    .X(clknet_leaf_95_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_96_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_96_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_97_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_97_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_98_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_98_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_99_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_99_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_100_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_100_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_101_clk_regs (.A(clknet_5_28__leaf_clk_regs),
    .X(clknet_leaf_101_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_102_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_102_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_103_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_103_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_104_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_104_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_105_clk_regs (.A(clknet_5_29__leaf_clk_regs),
    .X(clknet_leaf_105_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_106_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_106_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_107_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_107_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_108_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_108_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_109_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_109_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_110_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_110_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_111_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_111_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_112_clk_regs (.A(clknet_5_22__leaf_clk_regs),
    .X(clknet_leaf_112_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_113_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_113_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_114_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_114_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_115_clk_regs (.A(clknet_5_23__leaf_clk_regs),
    .X(clknet_leaf_115_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_116_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_116_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_117_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_117_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_118_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_118_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_119_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_119_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_120_clk_regs (.A(clknet_5_21__leaf_clk_regs),
    .X(clknet_leaf_120_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_121_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_121_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_122_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_122_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_123_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_123_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_124_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_124_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_125_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_125_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_126_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_126_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_127_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_127_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_128_clk_regs (.A(clknet_5_20__leaf_clk_regs),
    .X(clknet_leaf_128_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_129_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_129_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_130_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_130_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_131_clk_regs (.A(clknet_5_17__leaf_clk_regs),
    .X(clknet_leaf_131_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_132_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_132_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_133_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_133_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_134_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_134_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_135_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_135_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_136_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_136_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_137_clk_regs (.A(clknet_5_16__leaf_clk_regs),
    .X(clknet_leaf_137_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_138_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_138_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_139_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_139_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_140_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_140_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_141_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_141_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_142_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_142_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_143_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_143_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_144_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_144_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_145_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_145_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_146_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_146_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_147_clk_regs (.A(clknet_5_25__leaf_clk_regs),
    .X(clknet_leaf_147_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_148_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_148_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_149_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_149_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_150_clk_regs (.A(clknet_5_18__leaf_clk_regs),
    .X(clknet_leaf_150_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_151_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_151_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_152_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_152_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_153_clk_regs (.A(clknet_5_24__leaf_clk_regs),
    .X(clknet_leaf_153_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_154_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_154_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_155_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_155_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_156_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_156_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_157_clk_regs (.A(clknet_5_6__leaf_clk_regs),
    .X(clknet_leaf_157_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_158_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_158_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_159_clk_regs (.A(clknet_5_7__leaf_clk_regs),
    .X(clknet_leaf_159_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_160_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_160_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_161_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_161_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_162_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_162_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_163_clk_regs (.A(clknet_5_19__leaf_clk_regs),
    .X(clknet_leaf_163_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_164_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_164_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_165_clk_regs (.A(clknet_5_5__leaf_clk_regs),
    .X(clknet_leaf_165_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_166_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_166_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_167_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_167_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_168_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_168_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_169_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_169_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_170_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_170_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_171_clk_regs (.A(clknet_5_4__leaf_clk_regs),
    .X(clknet_leaf_171_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_172_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_172_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_173_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_173_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_174_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_174_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_175_clk_regs (.A(clknet_5_1__leaf_clk_regs),
    .X(clknet_leaf_175_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_176_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_176_clk_regs));
 sg13g2_buf_8 clkbuf_leaf_177_clk_regs (.A(clknet_5_0__leaf_clk_regs),
    .X(clknet_leaf_177_clk_regs));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_0_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_0_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_1_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_1_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_2_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_2_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_3_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_3_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_4_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_4_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_5_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_5_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_6_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_6_0_clk_regs));
 sg13g2_buf_8 clkbuf_3_7_0_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_3_7_0_clk_regs));
 sg13g2_buf_8 clkbuf_5_0__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_1__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_2__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_3__f_clk_regs (.A(clknet_3_0_0_clk_regs),
    .X(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_4__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_4__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_5__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_6__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_6__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_7__f_clk_regs (.A(clknet_3_1_0_clk_regs),
    .X(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_8__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_8__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_9__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_10__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_10__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_11__f_clk_regs (.A(clknet_3_2_0_clk_regs),
    .X(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_12__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_12__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_13__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_14__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_14__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_15__f_clk_regs (.A(clknet_3_3_0_clk_regs),
    .X(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_16__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_16__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_17__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_17__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_18__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_18__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_19__f_clk_regs (.A(clknet_3_4_0_clk_regs),
    .X(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_20__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_20__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_21__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_22__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_22__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_23__f_clk_regs (.A(clknet_3_5_0_clk_regs),
    .X(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_24__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_24__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_25__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_26__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_26__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_27__f_clk_regs (.A(clknet_3_6_0_clk_regs),
    .X(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_28__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_28__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_29__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_30__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_30__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_5_31__f_clk_regs (.A(clknet_3_7_0_clk_regs),
    .X(clknet_5_31__leaf_clk_regs));
 sg13g2_buf_8 clkload0 (.A(clknet_5_3__leaf_clk_regs));
 sg13g2_buf_8 clkload1 (.A(clknet_5_5__leaf_clk_regs));
 sg13g2_buf_8 clkload2 (.A(clknet_5_7__leaf_clk_regs));
 sg13g2_buf_8 clkload3 (.A(clknet_5_9__leaf_clk_regs));
 sg13g2_buf_8 clkload4 (.A(clknet_5_11__leaf_clk_regs));
 sg13g2_buf_8 clkload5 (.A(clknet_5_13__leaf_clk_regs));
 sg13g2_buf_8 clkload6 (.A(clknet_5_15__leaf_clk_regs));
 sg13g2_buf_8 clkload7 (.A(clknet_5_19__leaf_clk_regs));
 sg13g2_buf_8 clkload8 (.A(clknet_5_21__leaf_clk_regs));
 sg13g2_buf_8 clkload9 (.A(clknet_5_23__leaf_clk_regs));
 sg13g2_buf_8 clkload10 (.A(clknet_5_25__leaf_clk_regs));
 sg13g2_buf_8 clkload11 (.A(clknet_5_27__leaf_clk_regs));
 sg13g2_buf_8 clkload12 (.A(clknet_5_29__leaf_clk_regs));
 sg13g2_buf_8 clkload13 (.A(clknet_5_31__leaf_clk_regs));
 sg13g2_inv_4 clkload14 (.A(clknet_leaf_177_clk_regs));
 sg13g2_buf_8 delaybuf_0_clk (.A(delaynet_0_clk),
    .X(clknet_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net1436));
 sg13g2_dlygate4sd3_1 hold2 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[6] ),
    .X(net1437));
 sg13g2_dlygate4sd3_1 hold3 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1438));
 sg13g2_dlygate4sd3_1 hold4 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1439));
 sg13g2_dlygate4sd3_1 hold5 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1440));
 sg13g2_dlygate4sd3_1 hold6 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[14] ),
    .X(net1441));
 sg13g2_dlygate4sd3_1 hold7 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[15] ),
    .X(net1442));
 sg13g2_dlygate4sd3_1 hold8 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1443));
 sg13g2_dlygate4sd3_1 hold9 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net1444));
 sg13g2_dlygate4sd3_1 hold10 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1445));
 sg13g2_dlygate4sd3_1 hold11 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[0] ),
    .X(net1446));
 sg13g2_dlygate4sd3_1 hold12 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[28] ),
    .X(net1447));
 sg13g2_dlygate4sd3_1 hold13 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[30] ),
    .X(net1448));
 sg13g2_dlygate4sd3_1 hold14 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net1449));
 sg13g2_dlygate4sd3_1 hold15 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net1450));
 sg13g2_dlygate4sd3_1 hold16 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net1451));
 sg13g2_dlygate4sd3_1 hold17 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[15] ),
    .X(net1452));
 sg13g2_dlygate4sd3_1 hold18 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net1453));
 sg13g2_dlygate4sd3_1 hold19 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1454));
 sg13g2_dlygate4sd3_1 hold20 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net1455));
 sg13g2_dlygate4sd3_1 hold21 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net1456));
 sg13g2_dlygate4sd3_1 hold22 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net1457));
 sg13g2_dlygate4sd3_1 hold23 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1458));
 sg13g2_dlygate4sd3_1 hold24 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1459));
 sg13g2_dlygate4sd3_1 hold25 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[4] ),
    .X(net1460));
 sg13g2_dlygate4sd3_1 hold26 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net1461));
 sg13g2_dlygate4sd3_1 hold27 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1462));
 sg13g2_dlygate4sd3_1 hold28 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1463));
 sg13g2_dlygate4sd3_1 hold29 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net1464));
 sg13g2_dlygate4sd3_1 hold30 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1465));
 sg13g2_dlygate4sd3_1 hold31 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1466));
 sg13g2_dlygate4sd3_1 hold32 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net1467));
 sg13g2_dlygate4sd3_1 hold33 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[22] ),
    .X(net1468));
 sg13g2_dlygate4sd3_1 hold34 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[27] ),
    .X(net1469));
 sg13g2_dlygate4sd3_1 hold35 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1470));
 sg13g2_dlygate4sd3_1 hold36 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net1471));
 sg13g2_dlygate4sd3_1 hold37 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1472));
 sg13g2_dlygate4sd3_1 hold38 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net1473));
 sg13g2_dlygate4sd3_1 hold39 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1474));
 sg13g2_dlygate4sd3_1 hold40 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net1475));
 sg13g2_dlygate4sd3_1 hold41 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1476));
 sg13g2_dlygate4sd3_1 hold42 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1477));
 sg13g2_dlygate4sd3_1 hold43 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[10] ),
    .X(net1478));
 sg13g2_dlygate4sd3_1 hold44 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net1479));
 sg13g2_dlygate4sd3_1 hold45 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net1480));
 sg13g2_dlygate4sd3_1 hold46 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1481));
 sg13g2_dlygate4sd3_1 hold47 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net1482));
 sg13g2_dlygate4sd3_1 hold48 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net1483));
 sg13g2_dlygate4sd3_1 hold49 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1484));
 sg13g2_dlygate4sd3_1 hold50 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1485));
 sg13g2_dlygate4sd3_1 hold51 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[4] ),
    .X(net1486));
 sg13g2_dlygate4sd3_1 hold52 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1487));
 sg13g2_dlygate4sd3_1 hold53 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net1488));
 sg13g2_dlygate4sd3_1 hold54 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net1489));
 sg13g2_dlygate4sd3_1 hold55 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net1490));
 sg13g2_dlygate4sd3_1 hold56 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1491));
 sg13g2_dlygate4sd3_1 hold57 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net1492));
 sg13g2_dlygate4sd3_1 hold58 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[12] ),
    .X(net1493));
 sg13g2_dlygate4sd3_1 hold59 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1494));
 sg13g2_dlygate4sd3_1 hold60 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1495));
 sg13g2_dlygate4sd3_1 hold61 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1496));
 sg13g2_dlygate4sd3_1 hold62 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1497));
 sg13g2_dlygate4sd3_1 hold63 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[8] ),
    .X(net1498));
 sg13g2_dlygate4sd3_1 hold64 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net1499));
 sg13g2_dlygate4sd3_1 hold65 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1500));
 sg13g2_dlygate4sd3_1 hold66 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1501));
 sg13g2_dlygate4sd3_1 hold67 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[22] ),
    .X(net1502));
 sg13g2_dlygate4sd3_1 hold68 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1503));
 sg13g2_dlygate4sd3_1 hold69 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1504));
 sg13g2_dlygate4sd3_1 hold70 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1505));
 sg13g2_dlygate4sd3_1 hold71 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1506));
 sg13g2_dlygate4sd3_1 hold72 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1507));
 sg13g2_dlygate4sd3_1 hold73 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net1508));
 sg13g2_dlygate4sd3_1 hold74 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1509));
 sg13g2_dlygate4sd3_1 hold75 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1510));
 sg13g2_dlygate4sd3_1 hold76 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net1511));
 sg13g2_dlygate4sd3_1 hold77 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1512));
 sg13g2_dlygate4sd3_1 hold78 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1513));
 sg13g2_dlygate4sd3_1 hold79 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[10] ),
    .X(net1514));
 sg13g2_dlygate4sd3_1 hold80 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1515));
 sg13g2_dlygate4sd3_1 hold81 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net1516));
 sg13g2_dlygate4sd3_1 hold82 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1517));
 sg13g2_dlygate4sd3_1 hold83 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[18] ),
    .X(net1518));
 sg13g2_dlygate4sd3_1 hold84 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net1519));
 sg13g2_dlygate4sd3_1 hold85 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[7] ),
    .X(net1520));
 sg13g2_dlygate4sd3_1 hold86 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1521));
 sg13g2_dlygate4sd3_1 hold87 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[8] ),
    .X(net1522));
 sg13g2_dlygate4sd3_1 hold88 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net1523));
 sg13g2_dlygate4sd3_1 hold89 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1524));
 sg13g2_dlygate4sd3_1 hold90 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net1525));
 sg13g2_dlygate4sd3_1 hold91 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[25] ),
    .X(net1526));
 sg13g2_dlygate4sd3_1 hold92 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1527));
 sg13g2_dlygate4sd3_1 hold93 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net1528));
 sg13g2_dlygate4sd3_1 hold94 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1529));
 sg13g2_dlygate4sd3_1 hold95 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[25] ),
    .X(net1530));
 sg13g2_dlygate4sd3_1 hold96 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1531));
 sg13g2_dlygate4sd3_1 hold97 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net1532));
 sg13g2_dlygate4sd3_1 hold98 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1533));
 sg13g2_dlygate4sd3_1 hold99 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1534));
 sg13g2_dlygate4sd3_1 hold100 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[22] ),
    .X(net1535));
 sg13g2_dlygate4sd3_1 hold101 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net1536));
 sg13g2_dlygate4sd3_1 hold102 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net1537));
 sg13g2_dlygate4sd3_1 hold103 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net1538));
 sg13g2_dlygate4sd3_1 hold104 (.A(\ui_in_sync0[4] ),
    .X(net1539));
 sg13g2_dlygate4sd3_1 hold105 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net1540));
 sg13g2_dlygate4sd3_1 hold106 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net1541));
 sg13g2_dlygate4sd3_1 hold107 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[23] ),
    .X(net1542));
 sg13g2_dlygate4sd3_1 hold108 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1543));
 sg13g2_dlygate4sd3_1 hold109 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[16] ),
    .X(net1544));
 sg13g2_dlygate4sd3_1 hold110 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1545));
 sg13g2_dlygate4sd3_1 hold111 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net1546));
 sg13g2_dlygate4sd3_1 hold112 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[29] ),
    .X(net1547));
 sg13g2_dlygate4sd3_1 hold113 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net1548));
 sg13g2_dlygate4sd3_1 hold114 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net1549));
 sg13g2_dlygate4sd3_1 hold115 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net1550));
 sg13g2_dlygate4sd3_1 hold116 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1551));
 sg13g2_dlygate4sd3_1 hold117 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1552));
 sg13g2_dlygate4sd3_1 hold118 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1553));
 sg13g2_dlygate4sd3_1 hold119 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[30] ),
    .X(net1554));
 sg13g2_dlygate4sd3_1 hold120 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1555));
 sg13g2_dlygate4sd3_1 hold121 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1556));
 sg13g2_dlygate4sd3_1 hold122 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[7] ),
    .X(net1557));
 sg13g2_dlygate4sd3_1 hold123 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net1558));
 sg13g2_dlygate4sd3_1 hold124 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net1559));
 sg13g2_dlygate4sd3_1 hold125 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[26] ),
    .X(net1560));
 sg13g2_dlygate4sd3_1 hold126 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1561));
 sg13g2_dlygate4sd3_1 hold127 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[11] ),
    .X(net1562));
 sg13g2_dlygate4sd3_1 hold128 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[30] ),
    .X(net1563));
 sg13g2_dlygate4sd3_1 hold129 (.A(\ui_in_sync0[7] ),
    .X(net1564));
 sg13g2_dlygate4sd3_1 hold130 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net1565));
 sg13g2_dlygate4sd3_1 hold131 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1566));
 sg13g2_dlygate4sd3_1 hold132 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1567));
 sg13g2_dlygate4sd3_1 hold133 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[23] ),
    .X(net1568));
 sg13g2_dlygate4sd3_1 hold134 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net1569));
 sg13g2_dlygate4sd3_1 hold135 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[17] ),
    .X(net1570));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ui_in_sync0[5] ),
    .X(net1571));
 sg13g2_dlygate4sd3_1 hold137 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1572));
 sg13g2_dlygate4sd3_1 hold138 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1573));
 sg13g2_dlygate4sd3_1 hold139 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net1574));
 sg13g2_dlygate4sd3_1 hold140 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[9] ),
    .X(net1575));
 sg13g2_dlygate4sd3_1 hold141 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net1576));
 sg13g2_dlygate4sd3_1 hold142 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[13] ),
    .X(net1577));
 sg13g2_dlygate4sd3_1 hold143 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[15] ),
    .X(net1578));
 sg13g2_dlygate4sd3_1 hold144 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net1579));
 sg13g2_dlygate4sd3_1 hold145 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1580));
 sg13g2_dlygate4sd3_1 hold146 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1581));
 sg13g2_dlygate4sd3_1 hold147 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net1582));
 sg13g2_dlygate4sd3_1 hold148 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net1583));
 sg13g2_dlygate4sd3_1 hold149 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1584));
 sg13g2_dlygate4sd3_1 hold150 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1585));
 sg13g2_dlygate4sd3_1 hold151 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net1586));
 sg13g2_dlygate4sd3_1 hold152 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net1587));
 sg13g2_dlygate4sd3_1 hold153 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1588));
 sg13g2_dlygate4sd3_1 hold154 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[3] ),
    .X(net1589));
 sg13g2_dlygate4sd3_1 hold155 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[29] ),
    .X(net1590));
 sg13g2_dlygate4sd3_1 hold156 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net1591));
 sg13g2_dlygate4sd3_1 hold157 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1592));
 sg13g2_dlygate4sd3_1 hold158 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1593));
 sg13g2_dlygate4sd3_1 hold159 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net1594));
 sg13g2_dlygate4sd3_1 hold160 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1595));
 sg13g2_dlygate4sd3_1 hold161 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[29] ),
    .X(net1596));
 sg13g2_dlygate4sd3_1 hold162 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1597));
 sg13g2_dlygate4sd3_1 hold163 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net1598));
 sg13g2_dlygate4sd3_1 hold164 (.A(\ui_in_sync0[1] ),
    .X(net1599));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ui_in_sync0[3] ),
    .X(net1600));
 sg13g2_dlygate4sd3_1 hold166 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net1601));
 sg13g2_dlygate4sd3_1 hold167 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1602));
 sg13g2_dlygate4sd3_1 hold168 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net1603));
 sg13g2_dlygate4sd3_1 hold169 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net1604));
 sg13g2_dlygate4sd3_1 hold170 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net1605));
 sg13g2_dlygate4sd3_1 hold171 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[23] ),
    .X(net1606));
 sg13g2_dlygate4sd3_1 hold172 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net1607));
 sg13g2_dlygate4sd3_1 hold173 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[8] ),
    .X(net1608));
 sg13g2_dlygate4sd3_1 hold174 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1609));
 sg13g2_dlygate4sd3_1 hold175 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net1610));
 sg13g2_dlygate4sd3_1 hold176 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[19] ),
    .X(net1611));
 sg13g2_dlygate4sd3_1 hold177 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net1612));
 sg13g2_dlygate4sd3_1 hold178 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net1613));
 sg13g2_dlygate4sd3_1 hold179 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1614));
 sg13g2_dlygate4sd3_1 hold180 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net1615));
 sg13g2_dlygate4sd3_1 hold181 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net1616));
 sg13g2_dlygate4sd3_1 hold182 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1617));
 sg13g2_dlygate4sd3_1 hold183 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1618));
 sg13g2_dlygate4sd3_1 hold184 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[24] ),
    .X(net1619));
 sg13g2_dlygate4sd3_1 hold185 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[31] ),
    .X(net1620));
 sg13g2_dlygate4sd3_1 hold186 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[1] ),
    .X(net1621));
 sg13g2_dlygate4sd3_1 hold187 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net1622));
 sg13g2_dlygate4sd3_1 hold188 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1623));
 sg13g2_dlygate4sd3_1 hold189 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net1624));
 sg13g2_dlygate4sd3_1 hold190 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net1625));
 sg13g2_dlygate4sd3_1 hold191 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1626));
 sg13g2_dlygate4sd3_1 hold192 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[18] ),
    .X(net1627));
 sg13g2_dlygate4sd3_1 hold193 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net1628));
 sg13g2_dlygate4sd3_1 hold194 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1629));
 sg13g2_dlygate4sd3_1 hold195 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net1630));
 sg13g2_dlygate4sd3_1 hold196 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[16] ),
    .X(net1631));
 sg13g2_dlygate4sd3_1 hold197 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net1632));
 sg13g2_dlygate4sd3_1 hold198 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1633));
 sg13g2_dlygate4sd3_1 hold199 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[29] ),
    .X(net1634));
 sg13g2_dlygate4sd3_1 hold200 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[21] ),
    .X(net1635));
 sg13g2_dlygate4sd3_1 hold201 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net1636));
 sg13g2_dlygate4sd3_1 hold202 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[28] ),
    .X(net1637));
 sg13g2_dlygate4sd3_1 hold203 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net1638));
 sg13g2_dlygate4sd3_1 hold204 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net1639));
 sg13g2_dlygate4sd3_1 hold205 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net1640));
 sg13g2_dlygate4sd3_1 hold206 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1641));
 sg13g2_dlygate4sd3_1 hold207 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[21] ),
    .X(net1642));
 sg13g2_dlygate4sd3_1 hold208 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1643));
 sg13g2_dlygate4sd3_1 hold209 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[19] ),
    .X(net1644));
 sg13g2_dlygate4sd3_1 hold210 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[27] ),
    .X(net1645));
 sg13g2_dlygate4sd3_1 hold211 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net1646));
 sg13g2_dlygate4sd3_1 hold212 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1647));
 sg13g2_dlygate4sd3_1 hold213 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net1648));
 sg13g2_dlygate4sd3_1 hold214 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net1649));
 sg13g2_dlygate4sd3_1 hold215 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net1650));
 sg13g2_dlygate4sd3_1 hold216 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1651));
 sg13g2_dlygate4sd3_1 hold217 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net1652));
 sg13g2_dlygate4sd3_1 hold218 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1653));
 sg13g2_dlygate4sd3_1 hold219 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net1654));
 sg13g2_dlygate4sd3_1 hold220 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net1655));
 sg13g2_dlygate4sd3_1 hold221 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net1656));
 sg13g2_dlygate4sd3_1 hold222 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net1657));
 sg13g2_dlygate4sd3_1 hold223 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net1658));
 sg13g2_dlygate4sd3_1 hold224 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[26] ),
    .X(net1659));
 sg13g2_dlygate4sd3_1 hold225 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[9] ),
    .X(net1660));
 sg13g2_dlygate4sd3_1 hold226 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1661));
 sg13g2_dlygate4sd3_1 hold227 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[12] ),
    .X(net1662));
 sg13g2_dlygate4sd3_1 hold228 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net1663));
 sg13g2_dlygate4sd3_1 hold229 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[31] ),
    .X(net1664));
 sg13g2_dlygate4sd3_1 hold230 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net1665));
 sg13g2_dlygate4sd3_1 hold231 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net1666));
 sg13g2_dlygate4sd3_1 hold232 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net1667));
 sg13g2_dlygate4sd3_1 hold233 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[12] ),
    .X(net1668));
 sg13g2_dlygate4sd3_1 hold234 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net1669));
 sg13g2_dlygate4sd3_1 hold235 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[27] ),
    .X(net1670));
 sg13g2_dlygate4sd3_1 hold236 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net1671));
 sg13g2_dlygate4sd3_1 hold237 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[8] ),
    .X(net1672));
 sg13g2_dlygate4sd3_1 hold238 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1673));
 sg13g2_dlygate4sd3_1 hold239 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1674));
 sg13g2_dlygate4sd3_1 hold240 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net1675));
 sg13g2_dlygate4sd3_1 hold241 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[19] ),
    .X(net1676));
 sg13g2_dlygate4sd3_1 hold242 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net1677));
 sg13g2_dlygate4sd3_1 hold243 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net1678));
 sg13g2_dlygate4sd3_1 hold244 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net1679));
 sg13g2_dlygate4sd3_1 hold245 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net1680));
 sg13g2_dlygate4sd3_1 hold246 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net1681));
 sg13g2_dlygate4sd3_1 hold247 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2507));
 sg13g2_dlygate4sd3_1 hold248 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2508));
 sg13g2_dlygate4sd3_1 hold249 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2509));
 sg13g2_dlygate4sd3_1 hold250 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[31] ),
    .X(net2510));
 sg13g2_dlygate4sd3_1 hold251 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[25] ),
    .X(net2511));
 sg13g2_dlygate4sd3_1 hold252 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2512));
 sg13g2_dlygate4sd3_1 hold253 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2513));
 sg13g2_dlygate4sd3_1 hold254 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[5] ),
    .X(net2514));
 sg13g2_dlygate4sd3_1 hold255 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2515));
 sg13g2_dlygate4sd3_1 hold256 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2516));
 sg13g2_dlygate4sd3_1 hold257 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2517));
 sg13g2_dlygate4sd3_1 hold258 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2518));
 sg13g2_dlygate4sd3_1 hold259 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2519));
 sg13g2_dlygate4sd3_1 hold260 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2520));
 sg13g2_dlygate4sd3_1 hold261 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[17] ),
    .X(net2521));
 sg13g2_dlygate4sd3_1 hold262 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2522));
 sg13g2_dlygate4sd3_1 hold263 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2523));
 sg13g2_dlygate4sd3_1 hold264 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2524));
 sg13g2_dlygate4sd3_1 hold265 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2525));
 sg13g2_dlygate4sd3_1 hold266 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2526));
 sg13g2_dlygate4sd3_1 hold267 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[15] ),
    .X(net2527));
 sg13g2_dlygate4sd3_1 hold268 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2528));
 sg13g2_dlygate4sd3_1 hold269 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2529));
 sg13g2_dlygate4sd3_1 hold270 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[30] ),
    .X(net2530));
 sg13g2_dlygate4sd3_1 hold271 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[12] ),
    .X(net2531));
 sg13g2_dlygate4sd3_1 hold272 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2532));
 sg13g2_dlygate4sd3_1 hold273 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[23] ),
    .X(net2533));
 sg13g2_dlygate4sd3_1 hold274 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2534));
 sg13g2_dlygate4sd3_1 hold275 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2535));
 sg13g2_dlygate4sd3_1 hold276 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2536));
 sg13g2_dlygate4sd3_1 hold277 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[24] ),
    .X(net2537));
 sg13g2_dlygate4sd3_1 hold278 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2538));
 sg13g2_dlygate4sd3_1 hold279 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[20] ),
    .X(net2539));
 sg13g2_dlygate4sd3_1 hold280 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2540));
 sg13g2_dlygate4sd3_1 hold281 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[14] ),
    .X(net2541));
 sg13g2_dlygate4sd3_1 hold282 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2542));
 sg13g2_dlygate4sd3_1 hold283 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2543));
 sg13g2_dlygate4sd3_1 hold284 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[14] ),
    .X(net2544));
 sg13g2_dlygate4sd3_1 hold285 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2545));
 sg13g2_dlygate4sd3_1 hold286 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2546));
 sg13g2_dlygate4sd3_1 hold287 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2547));
 sg13g2_dlygate4sd3_1 hold288 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2548));
 sg13g2_dlygate4sd3_1 hold289 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2549));
 sg13g2_dlygate4sd3_1 hold290 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2550));
 sg13g2_dlygate4sd3_1 hold291 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2551));
 sg13g2_dlygate4sd3_1 hold292 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[11] ),
    .X(net2552));
 sg13g2_dlygate4sd3_1 hold293 (.A(\ui_in_sync0[6] ),
    .X(net2553));
 sg13g2_dlygate4sd3_1 hold294 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[5] ),
    .X(net2554));
 sg13g2_dlygate4sd3_1 hold295 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2555));
 sg13g2_dlygate4sd3_1 hold296 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2556));
 sg13g2_dlygate4sd3_1 hold297 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2557));
 sg13g2_dlygate4sd3_1 hold298 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2558));
 sg13g2_dlygate4sd3_1 hold299 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2559));
 sg13g2_dlygate4sd3_1 hold300 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2560));
 sg13g2_dlygate4sd3_1 hold301 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[13] ),
    .X(net2561));
 sg13g2_dlygate4sd3_1 hold302 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2562));
 sg13g2_dlygate4sd3_1 hold303 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2563));
 sg13g2_dlygate4sd3_1 hold304 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[20] ),
    .X(net2564));
 sg13g2_dlygate4sd3_1 hold305 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[24] ),
    .X(net2565));
 sg13g2_dlygate4sd3_1 hold306 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2566));
 sg13g2_dlygate4sd3_1 hold307 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2567));
 sg13g2_dlygate4sd3_1 hold308 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2568));
 sg13g2_dlygate4sd3_1 hold309 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2569));
 sg13g2_dlygate4sd3_1 hold310 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2570));
 sg13g2_dlygate4sd3_1 hold311 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2571));
 sg13g2_dlygate4sd3_1 hold312 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2572));
 sg13g2_dlygate4sd3_1 hold313 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[17] ),
    .X(net2573));
 sg13g2_dlygate4sd3_1 hold314 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2574));
 sg13g2_dlygate4sd3_1 hold315 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2575));
 sg13g2_dlygate4sd3_1 hold316 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[14] ),
    .X(net2576));
 sg13g2_dlygate4sd3_1 hold317 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[9] ),
    .X(net2577));
 sg13g2_dlygate4sd3_1 hold318 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[17] ),
    .X(net2578));
 sg13g2_dlygate4sd3_1 hold319 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[13] ),
    .X(net2579));
 sg13g2_dlygate4sd3_1 hold320 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2580));
 sg13g2_dlygate4sd3_1 hold321 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2581));
 sg13g2_dlygate4sd3_1 hold322 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2582));
 sg13g2_dlygate4sd3_1 hold323 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[27] ),
    .X(net2583));
 sg13g2_dlygate4sd3_1 hold324 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[18] ),
    .X(net2584));
 sg13g2_dlygate4sd3_1 hold325 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2585));
 sg13g2_dlygate4sd3_1 hold326 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2586));
 sg13g2_dlygate4sd3_1 hold327 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[24] ),
    .X(net2587));
 sg13g2_dlygate4sd3_1 hold328 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2588));
 sg13g2_dlygate4sd3_1 hold329 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[20] ),
    .X(net2589));
 sg13g2_dlygate4sd3_1 hold330 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[26] ),
    .X(net2590));
 sg13g2_dlygate4sd3_1 hold331 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[11] ),
    .X(net2591));
 sg13g2_dlygate4sd3_1 hold332 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2592));
 sg13g2_dlygate4sd3_1 hold333 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2593));
 sg13g2_dlygate4sd3_1 hold334 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2594));
 sg13g2_dlygate4sd3_1 hold335 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2595));
 sg13g2_dlygate4sd3_1 hold336 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2596));
 sg13g2_dlygate4sd3_1 hold337 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2597));
 sg13g2_dlygate4sd3_1 hold338 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[19] ),
    .X(net2598));
 sg13g2_dlygate4sd3_1 hold339 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[20] ),
    .X(net2599));
 sg13g2_dlygate4sd3_1 hold340 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2600));
 sg13g2_dlygate4sd3_1 hold341 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2601));
 sg13g2_dlygate4sd3_1 hold342 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[25] ),
    .X(net2602));
 sg13g2_dlygate4sd3_1 hold343 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2603));
 sg13g2_dlygate4sd3_1 hold344 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2604));
 sg13g2_dlygate4sd3_1 hold345 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2605));
 sg13g2_dlygate4sd3_1 hold346 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2606));
 sg13g2_dlygate4sd3_1 hold347 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2607));
 sg13g2_dlygate4sd3_1 hold348 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2608));
 sg13g2_dlygate4sd3_1 hold349 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[22] ),
    .X(net2609));
 sg13g2_dlygate4sd3_1 hold350 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[13] ),
    .X(net2610));
 sg13g2_dlygate4sd3_1 hold351 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2611));
 sg13g2_dlygate4sd3_1 hold352 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2612));
 sg13g2_dlygate4sd3_1 hold353 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2613));
 sg13g2_dlygate4sd3_1 hold354 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2614));
 sg13g2_dlygate4sd3_1 hold355 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[18] ),
    .X(net2615));
 sg13g2_dlygate4sd3_1 hold356 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2616));
 sg13g2_dlygate4sd3_1 hold357 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2617));
 sg13g2_dlygate4sd3_1 hold358 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2618));
 sg13g2_dlygate4sd3_1 hold359 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2619));
 sg13g2_dlygate4sd3_1 hold360 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2620));
 sg13g2_dlygate4sd3_1 hold361 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2621));
 sg13g2_dlygate4sd3_1 hold362 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2622));
 sg13g2_dlygate4sd3_1 hold363 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2623));
 sg13g2_dlygate4sd3_1 hold364 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2624));
 sg13g2_dlygate4sd3_1 hold365 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[21] ),
    .X(net2625));
 sg13g2_dlygate4sd3_1 hold366 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2626));
 sg13g2_dlygate4sd3_1 hold367 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2627));
 sg13g2_dlygate4sd3_1 hold368 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2628));
 sg13g2_dlygate4sd3_1 hold369 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2629));
 sg13g2_dlygate4sd3_1 hold370 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2630));
 sg13g2_dlygate4sd3_1 hold371 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2631));
 sg13g2_dlygate4sd3_1 hold372 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[21] ),
    .X(net2632));
 sg13g2_dlygate4sd3_1 hold373 (.A(\ui_in_sync0[0] ),
    .X(net2633));
 sg13g2_dlygate4sd3_1 hold374 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2634));
 sg13g2_dlygate4sd3_1 hold375 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2635));
 sg13g2_dlygate4sd3_1 hold376 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[2] ),
    .X(net2636));
 sg13g2_dlygate4sd3_1 hold377 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2637));
 sg13g2_dlygate4sd3_1 hold378 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[11] ),
    .X(net2638));
 sg13g2_dlygate4sd3_1 hold379 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2639));
 sg13g2_dlygate4sd3_1 hold380 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2640));
 sg13g2_dlygate4sd3_1 hold381 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[28] ),
    .X(net2641));
 sg13g2_dlygate4sd3_1 hold382 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2642));
 sg13g2_dlygate4sd3_1 hold383 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2643));
 sg13g2_dlygate4sd3_1 hold384 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2644));
 sg13g2_dlygate4sd3_1 hold385 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2645));
 sg13g2_dlygate4sd3_1 hold386 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2646));
 sg13g2_dlygate4sd3_1 hold387 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2647));
 sg13g2_dlygate4sd3_1 hold388 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2648));
 sg13g2_dlygate4sd3_1 hold389 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2649));
 sg13g2_dlygate4sd3_1 hold390 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2650));
 sg13g2_dlygate4sd3_1 hold391 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[6] ),
    .X(net2651));
 sg13g2_dlygate4sd3_1 hold392 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2652));
 sg13g2_dlygate4sd3_1 hold393 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2653));
 sg13g2_dlygate4sd3_1 hold394 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[28] ),
    .X(net2654));
 sg13g2_dlygate4sd3_1 hold395 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2655));
 sg13g2_dlygate4sd3_1 hold396 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[30] ),
    .X(net2656));
 sg13g2_dlygate4sd3_1 hold397 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[29] ),
    .X(net2657));
 sg13g2_dlygate4sd3_1 hold398 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2658));
 sg13g2_dlygate4sd3_1 hold399 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2659));
 sg13g2_dlygate4sd3_1 hold400 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[26] ),
    .X(net2660));
 sg13g2_dlygate4sd3_1 hold401 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[16] ),
    .X(net2661));
 sg13g2_dlygate4sd3_1 hold402 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2662));
 sg13g2_dlygate4sd3_1 hold403 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2663));
 sg13g2_dlygate4sd3_1 hold404 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[28] ),
    .X(net2664));
 sg13g2_dlygate4sd3_1 hold405 (.A(\i_tinyqv.cpu.i_core.i_instrret.reg_buf[31] ),
    .X(net2665));
 sg13g2_dlygate4sd3_1 hold406 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[7] ),
    .X(net2666));
 sg13g2_dlygate4sd3_1 hold407 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2667));
 sg13g2_dlygate4sd3_1 hold408 (.A(\ui_in_sync0[2] ),
    .X(net2668));
 sg13g2_dlygate4sd3_1 hold409 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[31] ),
    .X(net2669));
 sg13g2_dlygate4sd3_1 hold410 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2670));
 sg13g2_dlygate4sd3_1 hold411 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2671));
 sg13g2_dlygate4sd3_1 hold412 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2672));
 sg13g2_dlygate4sd3_1 hold413 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2673));
 sg13g2_dlygate4sd3_1 hold414 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2674));
 sg13g2_dlygate4sd3_1 hold415 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2675));
 sg13g2_dlygate4sd3_1 hold416 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[9] ),
    .X(net2676));
 sg13g2_dlygate4sd3_1 hold417 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2677));
 sg13g2_dlygate4sd3_1 hold418 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[13] ),
    .X(net2678));
 sg13g2_dlygate4sd3_1 hold419 (.A(\i_tinyqv.cpu.i_timer.i_mtime.reg_buf[10] ),
    .X(net2679));
 sg13g2_dlygate4sd3_1 hold420 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2680));
 sg13g2_dlygate4sd3_1 hold421 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[16] ),
    .X(net2681));
 sg13g2_dlygate4sd3_1 hold422 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[5].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2682));
 sg13g2_dlygate4sd3_1 hold423 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[17] ),
    .X(net2683));
 sg13g2_dlygate4sd3_1 hold424 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[10] ),
    .X(net2684));
 sg13g2_dlygate4sd3_1 hold425 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[20] ),
    .X(net2685));
 sg13g2_dlygate4sd3_1 hold426 (.A(\i_tinyqv.cpu.i_core.i_cycles.reg_buf[16] ),
    .X(net2686));
 sg13g2_dlygate4sd3_1 hold427 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[13].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2687));
 sg13g2_dlygate4sd3_1 hold428 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2688));
 sg13g2_dlygate4sd3_1 hold429 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[2].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2689));
 sg13g2_dlygate4sd3_1 hold430 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[19] ),
    .X(net2690));
 sg13g2_dlygate4sd3_1 hold431 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2691));
 sg13g2_dlygate4sd3_1 hold432 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2692));
 sg13g2_dlygate4sd3_1 hold433 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2693));
 sg13g2_dlygate4sd3_1 hold434 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[14] ),
    .X(net2694));
 sg13g2_dlygate4sd3_1 hold435 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[4] ),
    .X(net2695));
 sg13g2_dlygate4sd3_1 hold436 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[15] ),
    .X(net2696));
 sg13g2_dlygate4sd3_1 hold437 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2697));
 sg13g2_dlygate4sd3_1 hold438 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[5] ),
    .X(net2698));
 sg13g2_dlygate4sd3_1 hold439 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[12] ),
    .X(net2699));
 sg13g2_dlygate4sd3_1 hold440 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2700));
 sg13g2_dlygate4sd3_1 hold441 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[23] ),
    .X(net2701));
 sg13g2_dlygate4sd3_1 hold442 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2702));
 sg13g2_dlygate4sd3_1 hold443 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2703));
 sg13g2_dlygate4sd3_1 hold444 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2704));
 sg13g2_dlygate4sd3_1 hold445 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2705));
 sg13g2_dlygate4sd3_1 hold446 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[22] ),
    .X(net2706));
 sg13g2_dlygate4sd3_1 hold447 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[11] ),
    .X(net2707));
 sg13g2_dlygate4sd3_1 hold448 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2708));
 sg13g2_dlygate4sd3_1 hold449 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2709));
 sg13g2_dlygate4sd3_1 hold450 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[21] ),
    .X(net2710));
 sg13g2_dlygate4sd3_1 hold451 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[18] ),
    .X(net2711));
 sg13g2_dlygate4sd3_1 hold452 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2712));
 sg13g2_dlygate4sd3_1 hold453 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2713));
 sg13g2_dlygate4sd3_1 hold454 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2714));
 sg13g2_dlygate4sd3_1 hold455 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2715));
 sg13g2_dlygate4sd3_1 hold456 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2716));
 sg13g2_dlygate4sd3_1 hold457 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[14].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2717));
 sg13g2_dlygate4sd3_1 hold458 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2718));
 sg13g2_dlygate4sd3_1 hold459 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[12].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2719));
 sg13g2_dlygate4sd3_1 hold460 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[6].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2720));
 sg13g2_dlygate4sd3_1 hold461 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2721));
 sg13g2_dlygate4sd3_1 hold462 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2722));
 sg13g2_dlygate4sd3_1 hold463 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2723));
 sg13g2_dlygate4sd3_1 hold464 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2724));
 sg13g2_dlygate4sd3_1 hold465 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[10].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2725));
 sg13g2_dlygate4sd3_1 hold466 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2726));
 sg13g2_dlygate4sd3_1 hold467 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[7].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2727));
 sg13g2_dlygate4sd3_1 hold468 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[8].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2728));
 sg13g2_dlygate4sd3_1 hold469 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[10] ),
    .X(net2729));
 sg13g2_dlygate4sd3_1 hold470 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[9].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2730));
 sg13g2_dlygate4sd3_1 hold471 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[4] ),
    .X(net2731));
 sg13g2_dlygate4sd3_1 hold472 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2732));
 sg13g2_dlygate4sd3_1 hold473 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[15].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2733));
 sg13g2_dlygate4sd3_1 hold474 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[9] ),
    .X(net2734));
 sg13g2_dlygate4sd3_1 hold475 (.A(\i_tinyqv.cpu.i_core.cycle_count_wide[6] ),
    .X(net2735));
 sg13g2_dlygate4sd3_1 hold476 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[11].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2736));
 sg13g2_dlygate4sd3_1 hold477 (.A(\time_count[0] ),
    .X(net2737));
 sg13g2_dlygate4sd3_1 hold478 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[24] ),
    .X(net2738));
 sg13g2_dlygate4sd3_1 hold479 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[5] ),
    .X(net2739));
 sg13g2_dlygate4sd3_1 hold480 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[8] ),
    .X(net2740));
 sg13g2_dlygate4sd3_1 hold481 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[26] ),
    .X(net2741));
 sg13g2_dlygate4sd3_1 hold482 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[27] ),
    .X(net2742));
 sg13g2_dlygate4sd3_1 hold483 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[25] ),
    .X(net2743));
 sg13g2_dlygate4sd3_1 hold484 (.A(\i_debug_uart_tx.cycle_counter[4] ),
    .X(net2744));
 sg13g2_dlygate4sd3_1 hold485 (.A(_00431_),
    .X(net2745));
 sg13g2_dlygate4sd3_1 hold486 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[6] ),
    .X(net2746));
 sg13g2_dlygate4sd3_1 hold487 (.A(\i_tinyqv.cpu.i_core.i_registers.genblk1[1].genblk1.genblk1.gen_reg_normal.reg_buf[7] ),
    .X(net2747));
 sg13g2_dlygate4sd3_1 hold488 (.A(\i_peripherals.func_sel[25] ),
    .X(net2748));
 sg13g2_dlygate4sd3_1 hold489 (.A(_00560_),
    .X(net2749));
 sg13g2_dlygate4sd3_1 hold490 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[0] ),
    .X(net2750));
 sg13g2_dlygate4sd3_1 hold491 (.A(\i_peripherals.i_user_peri39.instr[10] ),
    .X(net2751));
 sg13g2_dlygate4sd3_1 hold492 (.A(_00206_),
    .X(net2752));
 sg13g2_dlygate4sd3_1 hold493 (.A(\i_peripherals.func_sel[13] ),
    .X(net2753));
 sg13g2_dlygate4sd3_1 hold494 (.A(_00572_),
    .X(net2754));
 sg13g2_dlygate4sd3_1 hold495 (.A(\i_peripherals.func_sel[23] ),
    .X(net2755));
 sg13g2_dlygate4sd3_1 hold496 (.A(_00570_),
    .X(net2756));
 sg13g2_dlygate4sd3_1 hold497 (.A(\i_peripherals.func_sel[37] ),
    .X(net2757));
 sg13g2_dlygate4sd3_1 hold498 (.A(_00548_),
    .X(net2758));
 sg13g2_dlygate4sd3_1 hold499 (.A(\i_peripherals.func_sel[19] ),
    .X(net2759));
 sg13g2_dlygate4sd3_1 hold500 (.A(_00566_),
    .X(net2760));
 sg13g2_dlygate4sd3_1 hold501 (.A(\i_peripherals.func_sel[21] ),
    .X(net2761));
 sg13g2_dlygate4sd3_1 hold502 (.A(_00568_),
    .X(net2762));
 sg13g2_dlygate4sd3_1 hold503 (.A(\i_peripherals.func_sel[17] ),
    .X(net2763));
 sg13g2_dlygate4sd3_1 hold504 (.A(_00576_),
    .X(net2764));
 sg13g2_dlygate4sd3_1 hold505 (.A(\i_peripherals.func_sel[35] ),
    .X(net2765));
 sg13g2_dlygate4sd3_1 hold506 (.A(_00558_),
    .X(net2766));
 sg13g2_dlygate4sd3_1 hold507 (.A(\i_peripherals.func_sel[29] ),
    .X(net2767));
 sg13g2_dlygate4sd3_1 hold508 (.A(_00564_),
    .X(net2768));
 sg13g2_dlygate4sd3_1 hold509 (.A(\i_peripherals.func_sel[3] ),
    .X(net2769));
 sg13g2_dlygate4sd3_1 hold510 (.A(_00382_),
    .X(net2770));
 sg13g2_dlygate4sd3_1 hold511 (.A(\i_peripherals.i_user_peri39.instr[8] ),
    .X(net2771));
 sg13g2_dlygate4sd3_1 hold512 (.A(_00204_),
    .X(net2772));
 sg13g2_dlygate4sd3_1 hold513 (.A(\i_peripherals.func_sel[5] ),
    .X(net2773));
 sg13g2_dlygate4sd3_1 hold514 (.A(_00384_),
    .X(net2774));
 sg13g2_dlygate4sd3_1 hold515 (.A(\i_tinyqv.cpu.load_started ),
    .X(net2775));
 sg13g2_dlygate4sd3_1 hold516 (.A(_00847_),
    .X(net2776));
 sg13g2_dlygate4sd3_1 hold517 (.A(\i_peripherals.func_sel[31] ),
    .X(net2777));
 sg13g2_dlygate4sd3_1 hold518 (.A(_00554_),
    .X(net2778));
 sg13g2_dlygate4sd3_1 hold519 (.A(\i_peripherals.i_user_peri39.instr[11] ),
    .X(net2779));
 sg13g2_dlygate4sd3_1 hold520 (.A(_00207_),
    .X(net2780));
 sg13g2_dlygate4sd3_1 hold521 (.A(\i_tinyqv.mem.q_ctrl.addr[0] ),
    .X(net2781));
 sg13g2_dlygate4sd3_1 hold522 (.A(_00129_),
    .X(net2782));
 sg13g2_dlygate4sd3_1 hold523 (.A(\i_peripherals.func_sel[11] ),
    .X(net2783));
 sg13g2_dlygate4sd3_1 hold524 (.A(_00582_),
    .X(net2784));
 sg13g2_dlygate4sd3_1 hold525 (.A(\i_tinyqv.cpu.instr_data[3][11] ),
    .X(net2785));
 sg13g2_dlygate4sd3_1 hold526 (.A(_00480_),
    .X(net2786));
 sg13g2_dlygate4sd3_1 hold527 (.A(\i_tinyqv.mem.qspi_data_buf[11] ),
    .X(net2787));
 sg13g2_dlygate4sd3_1 hold528 (.A(_00679_),
    .X(net2788));
 sg13g2_dlygate4sd3_1 hold529 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_a_select ),
    .X(net2789));
 sg13g2_dlygate4sd3_1 hold530 (.A(\i_peripherals.func_sel[33] ),
    .X(net2790));
 sg13g2_dlygate4sd3_1 hold531 (.A(_00556_),
    .X(net2791));
 sg13g2_dlygate4sd3_1 hold532 (.A(\i_tinyqv.cpu.instr_data[3][13] ),
    .X(net2792));
 sg13g2_dlygate4sd3_1 hold533 (.A(_00482_),
    .X(net2793));
 sg13g2_dlygate4sd3_1 hold534 (.A(\i_debug_uart_tx.data_to_send[7] ),
    .X(net2794));
 sg13g2_dlygate4sd3_1 hold535 (.A(_00426_),
    .X(net2795));
 sg13g2_dlygate4sd3_1 hold536 (.A(\i_peripherals.func_sel[9] ),
    .X(net2796));
 sg13g2_dlygate4sd3_1 hold537 (.A(_00580_),
    .X(net2797));
 sg13g2_dlygate4sd3_1 hold538 (.A(\i_tinyqv.cpu.instr_data[3][10] ),
    .X(net2798));
 sg13g2_dlygate4sd3_1 hold539 (.A(_00479_),
    .X(net2799));
 sg13g2_dlygate4sd3_1 hold540 (.A(\i_tinyqv.mem.q_ctrl.spi_ram_b_select ),
    .X(net2800));
 sg13g2_dlygate4sd3_1 hold541 (.A(\i_tinyqv.cpu.addr_offset[3] ),
    .X(net2801));
 sg13g2_dlygate4sd3_1 hold542 (.A(_00912_),
    .X(net2802));
 sg13g2_dlygate4sd3_1 hold543 (.A(\i_peripherals.func_sel[22] ),
    .X(net2803));
 sg13g2_dlygate4sd3_1 hold544 (.A(_00569_),
    .X(net2804));
 sg13g2_dlygate4sd3_1 hold545 (.A(\i_peripherals.i_user_peri39.instr[12] ),
    .X(net2805));
 sg13g2_dlygate4sd3_1 hold546 (.A(_00208_),
    .X(net2806));
 sg13g2_dlygate4sd3_1 hold547 (.A(\i_peripherals.i_user_peri39._GEN[89] ),
    .X(net2807));
 sg13g2_dlygate4sd3_1 hold548 (.A(_00780_),
    .X(net2808));
 sg13g2_dlygate4sd3_1 hold549 (.A(\i_tinyqv.mem.q_ctrl.addr[13] ),
    .X(net2809));
 sg13g2_dlygate4sd3_1 hold550 (.A(_00643_),
    .X(net2810));
 sg13g2_dlygate4sd3_1 hold551 (.A(\i_peripherals.i_user_peri39._GEN[91] ),
    .X(net2811));
 sg13g2_dlygate4sd3_1 hold552 (.A(_00782_),
    .X(net2812));
 sg13g2_dlygate4sd3_1 hold553 (.A(\i_tinyqv.cpu.instr_data[3][4] ),
    .X(net2813));
 sg13g2_dlygate4sd3_1 hold554 (.A(_00473_),
    .X(net2814));
 sg13g2_dlygate4sd3_1 hold555 (.A(\i_peripherals.func_sel[26] ),
    .X(net2815));
 sg13g2_dlygate4sd3_1 hold556 (.A(_00561_),
    .X(net2816));
 sg13g2_dlygate4sd3_1 hold557 (.A(\i_peripherals.i_user_peri39._GEN[57] ),
    .X(net2817));
 sg13g2_dlygate4sd3_1 hold558 (.A(_00286_),
    .X(net2818));
 sg13g2_dlygate4sd3_1 hold559 (.A(\i_peripherals.i_user_peri39._GEN[93] ),
    .X(net2819));
 sg13g2_dlygate4sd3_1 hold560 (.A(_00784_),
    .X(net2820));
 sg13g2_dlygate4sd3_1 hold561 (.A(\i_peripherals.func_sel[15] ),
    .X(net2821));
 sg13g2_dlygate4sd3_1 hold562 (.A(\i_peripherals.i_user_peri39._GEN[48] ),
    .X(net2822));
 sg13g2_dlygate4sd3_1 hold563 (.A(_00277_),
    .X(net2823));
 sg13g2_dlygate4sd3_1 hold564 (.A(\i_peripherals.func_sel[40] ),
    .X(net2824));
 sg13g2_dlygate4sd3_1 hold565 (.A(_00551_),
    .X(net2825));
 sg13g2_dlygate4sd3_1 hold566 (.A(\i_peripherals.i_user_peri39._GEN[90] ),
    .X(net2826));
 sg13g2_dlygate4sd3_1 hold567 (.A(_00781_),
    .X(net2827));
 sg13g2_dlygate4sd3_1 hold568 (.A(\i_tinyqv.cpu.i_core.mepc[23] ),
    .X(net2828));
 sg13g2_dlygate4sd3_1 hold569 (.A(_00120_),
    .X(net2829));
 sg13g2_dlygate4sd3_1 hold570 (.A(\i_tinyqv.cpu.instr_data[3][7] ),
    .X(net2830));
 sg13g2_dlygate4sd3_1 hold571 (.A(_00476_),
    .X(net2831));
 sg13g2_dlygate4sd3_1 hold572 (.A(\i_tinyqv.mem.data_from_read[19] ),
    .X(net2832));
 sg13g2_dlygate4sd3_1 hold573 (.A(_00687_),
    .X(net2833));
 sg13g2_dlygate4sd3_1 hold574 (.A(\i_tinyqv.cpu.imm[28] ),
    .X(net2834));
 sg13g2_dlygate4sd3_1 hold575 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[32] ),
    .X(net2835));
 sg13g2_dlygate4sd3_1 hold576 (.A(_00173_),
    .X(net2836));
 sg13g2_dlygate4sd3_1 hold577 (.A(\i_tinyqv.cpu.i_core.mepc[20] ),
    .X(net2837));
 sg13g2_dlygate4sd3_1 hold578 (.A(_00117_),
    .X(net2838));
 sg13g2_dlygate4sd3_1 hold579 (.A(\i_tinyqv.mem.data_from_read[17] ),
    .X(net2839));
 sg13g2_dlygate4sd3_1 hold580 (.A(_00685_),
    .X(net2840));
 sg13g2_dlygate4sd3_1 hold581 (.A(\i_peripherals.i_user_peri39._GEN[85] ),
    .X(net2841));
 sg13g2_dlygate4sd3_1 hold582 (.A(_00776_),
    .X(net2842));
 sg13g2_dlygate4sd3_1 hold583 (.A(\i_tinyqv.cpu.instr_data[3][14] ),
    .X(net2843));
 sg13g2_dlygate4sd3_1 hold584 (.A(_00483_),
    .X(net2844));
 sg13g2_dlygate4sd3_1 hold585 (.A(\i_peripherals.func_sel[8] ),
    .X(net2845));
 sg13g2_dlygate4sd3_1 hold586 (.A(\i_peripherals.func_sel[27] ),
    .X(net2846));
 sg13g2_dlygate4sd3_1 hold587 (.A(\i_peripherals.i_user_peri39._GEN[81] ),
    .X(net2847));
 sg13g2_dlygate4sd3_1 hold588 (.A(_00772_),
    .X(net2848));
 sg13g2_dlygate4sd3_1 hold589 (.A(\i_peripherals.i_user_peri39._GEN[56] ),
    .X(net2849));
 sg13g2_dlygate4sd3_1 hold590 (.A(_00285_),
    .X(net2850));
 sg13g2_dlygate4sd3_1 hold591 (.A(\i_tinyqv.mem.data_from_read[16] ),
    .X(net2851));
 sg13g2_dlygate4sd3_1 hold592 (.A(_00684_),
    .X(net2852));
 sg13g2_dlygate4sd3_1 hold593 (.A(\i_peripherals.i_user_peri39._GEN[62] ),
    .X(net2853));
 sg13g2_dlygate4sd3_1 hold594 (.A(_00291_),
    .X(net2854));
 sg13g2_dlygate4sd3_1 hold595 (.A(\i_tinyqv.cpu.i_core.mie[10] ),
    .X(net2855));
 sg13g2_dlygate4sd3_1 hold596 (.A(_00437_),
    .X(net2856));
 sg13g2_dlygate4sd3_1 hold597 (.A(\i_tinyqv.cpu.additional_mem_ops[2] ),
    .X(net2857));
 sg13g2_dlygate4sd3_1 hold598 (.A(_07218_),
    .X(net2858));
 sg13g2_dlygate4sd3_1 hold599 (.A(\i_tinyqv.cpu.i_core.mepc[22] ),
    .X(net2859));
 sg13g2_dlygate4sd3_1 hold600 (.A(_00119_),
    .X(net2860));
 sg13g2_dlygate4sd3_1 hold601 (.A(\i_tinyqv.cpu.i_core.mepc[21] ),
    .X(net2861));
 sg13g2_dlygate4sd3_1 hold602 (.A(_00118_),
    .X(net2862));
 sg13g2_dlygate4sd3_1 hold603 (.A(\i_tinyqv.cpu.instr_data[3][9] ),
    .X(net2863));
 sg13g2_dlygate4sd3_1 hold604 (.A(_00478_),
    .X(net2864));
 sg13g2_dlygate4sd3_1 hold605 (.A(\i_peripherals.i_user_peri39._GEN[49] ),
    .X(net2865));
 sg13g2_dlygate4sd3_1 hold606 (.A(_00278_),
    .X(net2866));
 sg13g2_dlygate4sd3_1 hold607 (.A(\i_tinyqv.mem.data_from_read[18] ),
    .X(net2867));
 sg13g2_dlygate4sd3_1 hold608 (.A(_00686_),
    .X(net2868));
 sg13g2_dlygate4sd3_1 hold609 (.A(\i_peripherals.func_sel[32] ),
    .X(net2869));
 sg13g2_dlygate4sd3_1 hold610 (.A(\i_tinyqv.cpu.instr_data[1][0] ),
    .X(net2870));
 sg13g2_dlygate4sd3_1 hold611 (.A(_00539_),
    .X(net2871));
 sg13g2_dlygate4sd3_1 hold612 (.A(\i_peripherals.i_user_peri39._GEN[114] ),
    .X(net2872));
 sg13g2_dlygate4sd3_1 hold613 (.A(_00247_),
    .X(net2873));
 sg13g2_dlygate4sd3_1 hold614 (.A(\i_peripherals.i_user_peri39._GEN[92] ),
    .X(net2874));
 sg13g2_dlygate4sd3_1 hold615 (.A(_00783_),
    .X(net2875));
 sg13g2_dlygate4sd3_1 hold616 (.A(\i_peripherals.i_user_peri39._GEN[88] ),
    .X(net2876));
 sg13g2_dlygate4sd3_1 hold617 (.A(_00779_),
    .X(net2877));
 sg13g2_dlygate4sd3_1 hold618 (.A(\i_peripherals.i_user_peri39._GEN[79] ),
    .X(net2878));
 sg13g2_dlygate4sd3_1 hold619 (.A(_00770_),
    .X(net2879));
 sg13g2_dlygate4sd3_1 hold620 (.A(\i_peripherals.i_user_peri39._GEN[83] ),
    .X(net2880));
 sg13g2_dlygate4sd3_1 hold621 (.A(_00774_),
    .X(net2881));
 sg13g2_dlygate4sd3_1 hold622 (.A(\i_tinyqv.mem.qspi_data_buf[12] ),
    .X(net2882));
 sg13g2_dlygate4sd3_1 hold623 (.A(_00680_),
    .X(net2883));
 sg13g2_dlygate4sd3_1 hold624 (.A(\i_peripherals.i_uart.i_uart_tx.fsm_state[1] ),
    .X(net2884));
 sg13g2_dlygate4sd3_1 hold625 (.A(_00333_),
    .X(net2885));
 sg13g2_dlygate4sd3_1 hold626 (.A(\i_peripherals.i_user_peri39._GEN[122] ),
    .X(net2886));
 sg13g2_dlygate4sd3_1 hold627 (.A(_00255_),
    .X(net2887));
 sg13g2_dlygate4sd3_1 hold628 (.A(\i_peripherals.func_sel[34] ),
    .X(net2888));
 sg13g2_dlygate4sd3_1 hold629 (.A(_00557_),
    .X(net2889));
 sg13g2_dlygate4sd3_1 hold630 (.A(\i_peripherals.func_sel[16] ),
    .X(net2890));
 sg13g2_dlygate4sd3_1 hold631 (.A(_00575_),
    .X(net2891));
 sg13g2_dlygate4sd3_1 hold632 (.A(\i_peripherals.func_sel[4] ),
    .X(net2892));
 sg13g2_dlygate4sd3_1 hold633 (.A(_00383_),
    .X(net2893));
 sg13g2_dlygate4sd3_1 hold634 (.A(\i_tinyqv.cpu.i_core.mie[9] ),
    .X(net2894));
 sg13g2_dlygate4sd3_1 hold635 (.A(_00438_),
    .X(net2895));
 sg13g2_dlygate4sd3_1 hold636 (.A(\i_peripherals.i_uart.i_uart_rx.bit_sample ),
    .X(net2896));
 sg13g2_dlygate4sd3_1 hold637 (.A(_00344_),
    .X(net2897));
 sg13g2_dlygate4sd3_1 hold638 (.A(\i_peripherals.i_user_peri39._GEN[63] ),
    .X(net2898));
 sg13g2_dlygate4sd3_1 hold639 (.A(_00292_),
    .X(net2899));
 sg13g2_dlygate4sd3_1 hold640 (.A(\i_peripherals.i_user_peri39._GEN[59] ),
    .X(net2900));
 sg13g2_dlygate4sd3_1 hold641 (.A(_00288_),
    .X(net2901));
 sg13g2_dlygate4sd3_1 hold642 (.A(\i_peripherals.i_user_peri39._GEN[80] ),
    .X(net2902));
 sg13g2_dlygate4sd3_1 hold643 (.A(_00771_),
    .X(net2903));
 sg13g2_dlygate4sd3_1 hold644 (.A(\i_peripherals.i_user_peri39._GEN[39] ),
    .X(net2904));
 sg13g2_dlygate4sd3_1 hold645 (.A(_00268_),
    .X(net2905));
 sg13g2_dlygate4sd3_1 hold646 (.A(\i_tinyqv.cpu.imm[24] ),
    .X(net2906));
 sg13g2_dlygate4sd3_1 hold647 (.A(\i_tinyqv.cpu.instr_data[1][1] ),
    .X(net2907));
 sg13g2_dlygate4sd3_1 hold648 (.A(_00540_),
    .X(net2908));
 sg13g2_dlygate4sd3_1 hold649 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[12] ),
    .X(net2909));
 sg13g2_dlygate4sd3_1 hold650 (.A(_05403_),
    .X(net2910));
 sg13g2_dlygate4sd3_1 hold651 (.A(\i_peripherals.i_user_peri39._GEN[53] ),
    .X(net2911));
 sg13g2_dlygate4sd3_1 hold652 (.A(_00282_),
    .X(net2912));
 sg13g2_dlygate4sd3_1 hold653 (.A(\i_peripherals.i_user_peri39._GEN[86] ),
    .X(net2913));
 sg13g2_dlygate4sd3_1 hold654 (.A(_00777_),
    .X(net2914));
 sg13g2_dlygate4sd3_1 hold655 (.A(\i_peripherals.func_sel[20] ),
    .X(net2915));
 sg13g2_dlygate4sd3_1 hold656 (.A(\i_tinyqv.mem.q_ctrl.addr[17] ),
    .X(net2916));
 sg13g2_dlygate4sd3_1 hold657 (.A(_00647_),
    .X(net2917));
 sg13g2_dlygate4sd3_1 hold658 (.A(\i_peripherals.i_user_peri39._GEN[126] ),
    .X(net2918));
 sg13g2_dlygate4sd3_1 hold659 (.A(_00259_),
    .X(net2919));
 sg13g2_dlygate4sd3_1 hold660 (.A(\i_peripherals.func_sel[10] ),
    .X(net2920));
 sg13g2_dlygate4sd3_1 hold661 (.A(_00581_),
    .X(net2921));
 sg13g2_dlygate4sd3_1 hold662 (.A(\i_peripherals.i_user_peri39._GEN[103] ),
    .X(net2922));
 sg13g2_dlygate4sd3_1 hold663 (.A(_00236_),
    .X(net2923));
 sg13g2_dlygate4sd3_1 hold664 (.A(\i_peripherals.i_user_peri39._GEN[123] ),
    .X(net2924));
 sg13g2_dlygate4sd3_1 hold665 (.A(_00256_),
    .X(net2925));
 sg13g2_dlygate4sd3_1 hold666 (.A(\i_peripherals.i_user_peri39._GEN[112] ),
    .X(net2926));
 sg13g2_dlygate4sd3_1 hold667 (.A(_00245_),
    .X(net2927));
 sg13g2_dlygate4sd3_1 hold668 (.A(\i_peripherals.i_user_peri39._GEN[101] ),
    .X(net2928));
 sg13g2_dlygate4sd3_1 hold669 (.A(\i_tinyqv.cpu.instr_data[0][0] ),
    .X(net2929));
 sg13g2_dlygate4sd3_1 hold670 (.A(_00654_),
    .X(net2930));
 sg13g2_dlygate4sd3_1 hold671 (.A(\i_tinyqv.mem.qspi_data_buf[10] ),
    .X(net2931));
 sg13g2_dlygate4sd3_1 hold672 (.A(_00678_),
    .X(net2932));
 sg13g2_dlygate4sd3_1 hold673 (.A(\i_peripherals.i_user_peri39._GEN[125] ),
    .X(net2933));
 sg13g2_dlygate4sd3_1 hold674 (.A(_00258_),
    .X(net2934));
 sg13g2_dlygate4sd3_1 hold675 (.A(\i_peripherals.i_user_peri39._GEN[78] ),
    .X(net2935));
 sg13g2_dlygate4sd3_1 hold676 (.A(_00769_),
    .X(net2936));
 sg13g2_dlygate4sd3_1 hold677 (.A(\i_tinyqv.cpu.i_core.mcause[2] ),
    .X(net2937));
 sg13g2_dlygate4sd3_1 hold678 (.A(_02697_),
    .X(net2938));
 sg13g2_dlygate4sd3_1 hold679 (.A(\i_peripherals.i_user_peri39._GEN[120] ),
    .X(net2939));
 sg13g2_dlygate4sd3_1 hold680 (.A(_00253_),
    .X(net2940));
 sg13g2_dlygate4sd3_1 hold681 (.A(\i_peripherals.func_sel[0] ),
    .X(net2941));
 sg13g2_dlygate4sd3_1 hold682 (.A(_00379_),
    .X(net2942));
 sg13g2_dlygate4sd3_1 hold683 (.A(\i_tinyqv.cpu.instr_data[0][1] ),
    .X(net2943));
 sg13g2_dlygate4sd3_1 hold684 (.A(_00655_),
    .X(net2944));
 sg13g2_dlygate4sd3_1 hold685 (.A(\i_peripherals.i_user_peri39._GEN[0] ),
    .X(net2945));
 sg13g2_dlygate4sd3_1 hold686 (.A(\i_peripherals.gpio_out[7] ),
    .X(net2946));
 sg13g2_dlygate4sd3_1 hold687 (.A(_00378_),
    .X(net2947));
 sg13g2_dlygate4sd3_1 hold688 (.A(\i_peripherals.func_sel[38] ),
    .X(net2948));
 sg13g2_dlygate4sd3_1 hold689 (.A(\i_tinyqv.mem.qspi_data_buf[8] ),
    .X(net2949));
 sg13g2_dlygate4sd3_1 hold690 (.A(_00676_),
    .X(net2950));
 sg13g2_dlygate4sd3_1 hold691 (.A(\i_peripherals.i_user_peri39._GEN[117] ),
    .X(net2951));
 sg13g2_dlygate4sd3_1 hold692 (.A(_00250_),
    .X(net2952));
 sg13g2_dlygate4sd3_1 hold693 (.A(\i_peripherals.i_user_peri39._GEN[82] ),
    .X(net2953));
 sg13g2_dlygate4sd3_1 hold694 (.A(_00773_),
    .X(net2954));
 sg13g2_dlygate4sd3_1 hold695 (.A(\i_peripherals.i_user_peri39._GEN[60] ),
    .X(net2955));
 sg13g2_dlygate4sd3_1 hold696 (.A(_00289_),
    .X(net2956));
 sg13g2_dlygate4sd3_1 hold697 (.A(\i_tinyqv.mem.data_stall ),
    .X(net2957));
 sg13g2_dlygate4sd3_1 hold698 (.A(_06502_),
    .X(net2958));
 sg13g2_dlygate4sd3_1 hold699 (.A(_00662_),
    .X(net2959));
 sg13g2_dlygate4sd3_1 hold700 (.A(\i_peripherals.i_user_peri39._GEN[50] ),
    .X(net2960));
 sg13g2_dlygate4sd3_1 hold701 (.A(_00279_),
    .X(net2961));
 sg13g2_dlygate4sd3_1 hold702 (.A(\i_peripherals.i_user_peri39._GEN[2] ),
    .X(net2962));
 sg13g2_dlygate4sd3_1 hold703 (.A(_00231_),
    .X(net2963));
 sg13g2_dlygate4sd3_1 hold704 (.A(\i_peripherals.i_user_peri39._GEN[46] ),
    .X(net2964));
 sg13g2_dlygate4sd3_1 hold705 (.A(_00275_),
    .X(net2965));
 sg13g2_dlygate4sd3_1 hold706 (.A(\i_peripherals.gpio_out[1] ),
    .X(net2966));
 sg13g2_dlygate4sd3_1 hold707 (.A(_00372_),
    .X(net2967));
 sg13g2_dlygate4sd3_1 hold708 (.A(\i_tinyqv.cpu.i_core.load_done ),
    .X(net2968));
 sg13g2_dlygate4sd3_1 hold709 (.A(\i_peripherals.i_user_peri39._GEN[37] ),
    .X(net2969));
 sg13g2_dlygate4sd3_1 hold710 (.A(\i_peripherals.i_user_peri39._GEN[41] ),
    .X(net2970));
 sg13g2_dlygate4sd3_1 hold711 (.A(_00270_),
    .X(net2971));
 sg13g2_dlygate4sd3_1 hold712 (.A(\i_peripherals.i_user_peri39._GEN[58] ),
    .X(net2972));
 sg13g2_dlygate4sd3_1 hold713 (.A(_00287_),
    .X(net2973));
 sg13g2_dlygate4sd3_1 hold714 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[2] ),
    .X(net2974));
 sg13g2_dlygate4sd3_1 hold715 (.A(_05491_),
    .X(net2975));
 sg13g2_dlygate4sd3_1 hold716 (.A(_00360_),
    .X(net2976));
 sg13g2_dlygate4sd3_1 hold717 (.A(\i_peripherals.i_user_peri39._GEN[109] ),
    .X(net2977));
 sg13g2_dlygate4sd3_1 hold718 (.A(_00242_),
    .X(net2978));
 sg13g2_dlygate4sd3_1 hold719 (.A(\i_peripherals.i_user_peri39._GEN[124] ),
    .X(net2979));
 sg13g2_dlygate4sd3_1 hold720 (.A(_00257_),
    .X(net2980));
 sg13g2_dlygate4sd3_1 hold721 (.A(\i_peripherals.i_user_peri39._GEN[51] ),
    .X(net2981));
 sg13g2_dlygate4sd3_1 hold722 (.A(_00280_),
    .X(net2982));
 sg13g2_dlygate4sd3_1 hold723 (.A(\i_peripherals.i_user_peri39._GEN[54] ),
    .X(net2983));
 sg13g2_dlygate4sd3_1 hold724 (.A(_00283_),
    .X(net2984));
 sg13g2_dlygate4sd3_1 hold725 (.A(\i_peripherals.i_user_peri39._GEN[65] ),
    .X(net2985));
 sg13g2_dlygate4sd3_1 hold726 (.A(_00756_),
    .X(net2986));
 sg13g2_dlygate4sd3_1 hold727 (.A(\i_peripherals.i_user_peri39._GEN[61] ),
    .X(net2987));
 sg13g2_dlygate4sd3_1 hold728 (.A(_00290_),
    .X(net2988));
 sg13g2_dlygate4sd3_1 hold729 (.A(\i_tinyqv.cpu.instr_data[3][1] ),
    .X(net2989));
 sg13g2_dlygate4sd3_1 hold730 (.A(_00296_),
    .X(net2990));
 sg13g2_dlygate4sd3_1 hold731 (.A(\addr[12] ),
    .X(net2991));
 sg13g2_dlygate4sd3_1 hold732 (.A(_00860_),
    .X(net2992));
 sg13g2_dlygate4sd3_1 hold733 (.A(\i_peripherals.i_user_peri39._GEN[105] ),
    .X(net2993));
 sg13g2_dlygate4sd3_1 hold734 (.A(_00238_),
    .X(net2994));
 sg13g2_dlygate4sd3_1 hold735 (.A(\i_peripherals.i_user_peri39._GEN[102] ),
    .X(net2995));
 sg13g2_dlygate4sd3_1 hold736 (.A(_00235_),
    .X(net2996));
 sg13g2_dlygate4sd3_1 hold737 (.A(\i_tinyqv.cpu.i_core.time_hi[2] ),
    .X(net2997));
 sg13g2_dlygate4sd3_1 hold738 (.A(_00109_),
    .X(net2998));
 sg13g2_dlygate4sd3_1 hold739 (.A(_00074_),
    .X(net2999));
 sg13g2_dlygate4sd3_1 hold740 (.A(_00537_),
    .X(net3000));
 sg13g2_dlygate4sd3_1 hold741 (.A(\i_peripherals.i_user_peri39._GEN[115] ),
    .X(net3001));
 sg13g2_dlygate4sd3_1 hold742 (.A(_00248_),
    .X(net3002));
 sg13g2_dlygate4sd3_1 hold743 (.A(\i_peripherals.i_user_peri39.instr[0] ),
    .X(net3003));
 sg13g2_dlygate4sd3_1 hold744 (.A(_00196_),
    .X(net3004));
 sg13g2_dlygate4sd3_1 hold745 (.A(\i_peripherals.i_user_peri39._GEN[95] ),
    .X(net3005));
 sg13g2_dlygate4sd3_1 hold746 (.A(_00786_),
    .X(net3006));
 sg13g2_dlygate4sd3_1 hold747 (.A(\i_tinyqv.cpu.i_core.load_top_bit ),
    .X(net3007));
 sg13g2_dlygate4sd3_1 hold748 (.A(_00752_),
    .X(net3008));
 sg13g2_dlygate4sd3_1 hold749 (.A(\i_tinyqv.mem.data_from_read[20] ),
    .X(net3009));
 sg13g2_dlygate4sd3_1 hold750 (.A(_00688_),
    .X(net3010));
 sg13g2_dlygate4sd3_1 hold751 (.A(\i_peripherals.i_user_peri39._GEN[119] ),
    .X(net3011));
 sg13g2_dlygate4sd3_1 hold752 (.A(_00252_),
    .X(net3012));
 sg13g2_dlygate4sd3_1 hold753 (.A(\i_peripherals.i_user_peri39._GEN[55] ),
    .X(net3013));
 sg13g2_dlygate4sd3_1 hold754 (.A(_00284_),
    .X(net3014));
 sg13g2_dlygate4sd3_1 hold755 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[10] ),
    .X(net3015));
 sg13g2_dlygate4sd3_1 hold756 (.A(_05505_),
    .X(net3016));
 sg13g2_dlygate4sd3_1 hold757 (.A(_00368_),
    .X(net3017));
 sg13g2_dlygate4sd3_1 hold758 (.A(\i_tinyqv.mem.qspi_data_buf[9] ),
    .X(net3018));
 sg13g2_dlygate4sd3_1 hold759 (.A(_00677_),
    .X(net3019));
 sg13g2_dlygate4sd3_1 hold760 (.A(\i_peripherals.i_user_peri39._GEN[77] ),
    .X(net3020));
 sg13g2_dlygate4sd3_1 hold761 (.A(_00768_),
    .X(net3021));
 sg13g2_dlygate4sd3_1 hold762 (.A(\i_peripherals.i_user_peri39.busy_counter[0] ),
    .X(net3022));
 sg13g2_dlygate4sd3_1 hold763 (.A(_00293_),
    .X(net3023));
 sg13g2_dlygate4sd3_1 hold764 (.A(\i_peripherals.func_sel[28] ),
    .X(net3024));
 sg13g2_dlygate4sd3_1 hold765 (.A(_00563_),
    .X(net3025));
 sg13g2_dlygate4sd3_1 hold766 (.A(\i_peripherals.i_user_peri39._GEN[110] ),
    .X(net3026));
 sg13g2_dlygate4sd3_1 hold767 (.A(_00243_),
    .X(net3027));
 sg13g2_dlygate4sd3_1 hold768 (.A(\i_peripherals.i_user_peri39._GEN[45] ),
    .X(net3028));
 sg13g2_dlygate4sd3_1 hold769 (.A(_00274_),
    .X(net3029));
 sg13g2_dlygate4sd3_1 hold770 (.A(\i_peripherals.i_user_peri39._GEN[100] ),
    .X(net3030));
 sg13g2_dlygate4sd3_1 hold771 (.A(_00233_),
    .X(net3031));
 sg13g2_dlygate4sd3_1 hold772 (.A(\i_peripherals.i_user_peri39._GEN[69] ),
    .X(net3032));
 sg13g2_dlygate4sd3_1 hold773 (.A(\i_peripherals.i_user_peri39._GEN[33] ),
    .X(net3033));
 sg13g2_dlygate4sd3_1 hold774 (.A(_00262_),
    .X(net3034));
 sg13g2_dlygate4sd3_1 hold775 (.A(\i_peripherals.i_user_peri39._GEN[32] ),
    .X(net3035));
 sg13g2_dlygate4sd3_1 hold776 (.A(\i_peripherals.i_user_peri39._GEN[35] ),
    .X(net3036));
 sg13g2_dlygate4sd3_1 hold777 (.A(_00264_),
    .X(net3037));
 sg13g2_dlygate4sd3_1 hold778 (.A(\i_tinyqv.cpu.i_core.is_double_fault_r ),
    .X(net3038));
 sg13g2_dlygate4sd3_1 hold779 (.A(\i_tinyqv.cpu.imm[30] ),
    .X(net3039));
 sg13g2_dlygate4sd3_1 hold780 (.A(\i_peripherals.i_user_peri39._GEN[36] ),
    .X(net3040));
 sg13g2_dlygate4sd3_1 hold781 (.A(_00265_),
    .X(net3041));
 sg13g2_dlygate4sd3_1 hold782 (.A(\i_tinyqv.cpu.imm[27] ),
    .X(net3042));
 sg13g2_dlygate4sd3_1 hold783 (.A(\addr[22] ),
    .X(net3043));
 sg13g2_dlygate4sd3_1 hold784 (.A(_00870_),
    .X(net3044));
 sg13g2_dlygate4sd3_1 hold785 (.A(\i_tinyqv.cpu.instr_data_in[4] ),
    .X(net3045));
 sg13g2_dlygate4sd3_1 hold786 (.A(_00672_),
    .X(net3046));
 sg13g2_dlygate4sd3_1 hold787 (.A(\i_peripherals.i_user_peri39._GEN[34] ),
    .X(net3047));
 sg13g2_dlygate4sd3_1 hold788 (.A(_00263_),
    .X(net3048));
 sg13g2_dlygate4sd3_1 hold789 (.A(\i_peripherals.i_user_peri39._GEN[87] ),
    .X(net3049));
 sg13g2_dlygate4sd3_1 hold790 (.A(_00778_),
    .X(net3050));
 sg13g2_dlygate4sd3_1 hold791 (.A(\i_peripherals.i_user_peri39._GEN[127] ),
    .X(net3051));
 sg13g2_dlygate4sd3_1 hold792 (.A(_00260_),
    .X(net3052));
 sg13g2_dlygate4sd3_1 hold793 (.A(\i_tinyqv.cpu.imm[26] ),
    .X(net3053));
 sg13g2_dlygate4sd3_1 hold794 (.A(\i_peripherals.gpio_out[0] ),
    .X(net3054));
 sg13g2_dlygate4sd3_1 hold795 (.A(_00371_),
    .X(net3055));
 sg13g2_dlygate4sd3_1 hold796 (.A(\i_tinyqv.cpu.instr_data[1][14] ),
    .X(net3056));
 sg13g2_dlygate4sd3_1 hold797 (.A(_02649_),
    .X(net3057));
 sg13g2_dlygate4sd3_1 hold798 (.A(_00090_),
    .X(net3058));
 sg13g2_dlygate4sd3_1 hold799 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[28] ),
    .X(net3059));
 sg13g2_dlygate4sd3_1 hold800 (.A(\i_tinyqv.cpu.i_core.mcause[5] ),
    .X(net3060));
 sg13g2_dlygate4sd3_1 hold801 (.A(_02701_),
    .X(net3061));
 sg13g2_dlygate4sd3_1 hold802 (.A(\i_tinyqv.cpu.is_alu_reg ),
    .X(net3062));
 sg13g2_dlygate4sd3_1 hold803 (.A(\i_peripherals.i_uart.rxd_select ),
    .X(net3063));
 sg13g2_dlygate4sd3_1 hold804 (.A(_00310_),
    .X(net3064));
 sg13g2_dlygate4sd3_1 hold805 (.A(\i_peripherals.func_sel[14] ),
    .X(net3065));
 sg13g2_dlygate4sd3_1 hold806 (.A(\i_peripherals.i_user_peri39._GEN[47] ),
    .X(net3066));
 sg13g2_dlygate4sd3_1 hold807 (.A(_00276_),
    .X(net3067));
 sg13g2_dlygate4sd3_1 hold808 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[3] ),
    .X(net3068));
 sg13g2_dlygate4sd3_1 hold809 (.A(_05387_),
    .X(net3069));
 sg13g2_dlygate4sd3_1 hold810 (.A(_00322_),
    .X(net3070));
 sg13g2_dlygate4sd3_1 hold811 (.A(\i_tinyqv.cpu.imm[25] ),
    .X(net3071));
 sg13g2_dlygate4sd3_1 hold812 (.A(\i_peripherals.i_user_peri39._GEN[1] ),
    .X(net3072));
 sg13g2_dlygate4sd3_1 hold813 (.A(_00230_),
    .X(net3073));
 sg13g2_dlygate4sd3_1 hold814 (.A(\i_peripherals.func_sel[6] ),
    .X(net3074));
 sg13g2_dlygate4sd3_1 hold815 (.A(_00577_),
    .X(net3075));
 sg13g2_dlygate4sd3_1 hold816 (.A(\i_tinyqv.cpu.instr_data[2][14] ),
    .X(net3076));
 sg13g2_dlygate4sd3_1 hold817 (.A(_06780_),
    .X(net3077));
 sg13g2_dlygate4sd3_1 hold818 (.A(_00750_),
    .X(net3078));
 sg13g2_dlygate4sd3_1 hold819 (.A(\i_tinyqv.cpu.instr_data[2][11] ),
    .X(net3079));
 sg13g2_dlygate4sd3_1 hold820 (.A(_00747_),
    .X(net3080));
 sg13g2_dlygate4sd3_1 hold821 (.A(\i_tinyqv.cpu.instr_data[0][10] ),
    .X(net3081));
 sg13g2_dlygate4sd3_1 hold822 (.A(_00465_),
    .X(net3082));
 sg13g2_dlygate4sd3_1 hold823 (.A(\i_tinyqv.cpu.instr_data[0][7] ),
    .X(net3083));
 sg13g2_dlygate4sd3_1 hold824 (.A(_00462_),
    .X(net3084));
 sg13g2_dlygate4sd3_1 hold825 (.A(\i_peripherals.i_user_peri39._GEN[113] ),
    .X(net3085));
 sg13g2_dlygate4sd3_1 hold826 (.A(_00246_),
    .X(net3086));
 sg13g2_dlygate4sd3_1 hold827 (.A(\i_tinyqv.mem.qspi_data_buf[13] ),
    .X(net3087));
 sg13g2_dlygate4sd3_1 hold828 (.A(_00681_),
    .X(net3088));
 sg13g2_dlygate4sd3_1 hold829 (.A(\i_tinyqv.cpu.instr_data[1][13] ),
    .X(net3089));
 sg13g2_dlygate4sd3_1 hold830 (.A(_00089_),
    .X(net3090));
 sg13g2_dlygate4sd3_1 hold831 (.A(\i_peripherals.func_sel[2] ),
    .X(net3091));
 sg13g2_dlygate4sd3_1 hold832 (.A(_00381_),
    .X(net3092));
 sg13g2_dlygate4sd3_1 hold833 (.A(\i_peripherals.gpio_out[2] ),
    .X(net3093));
 sg13g2_dlygate4sd3_1 hold834 (.A(_00373_),
    .X(net3094));
 sg13g2_dlygate4sd3_1 hold835 (.A(\addr[16] ),
    .X(net3095));
 sg13g2_dlygate4sd3_1 hold836 (.A(_00864_),
    .X(net3096));
 sg13g2_dlygate4sd3_1 hold837 (.A(\i_tinyqv.cpu.i_core.mstatus_mpie ),
    .X(net3097));
 sg13g2_dlygate4sd3_1 hold838 (.A(_00123_),
    .X(net3098));
 sg13g2_dlygate4sd3_1 hold839 (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[0] ),
    .X(net3099));
 sg13g2_dlygate4sd3_1 hold840 (.A(\i_peripherals.i_user_peri39._GEN[70] ),
    .X(net3100));
 sg13g2_dlygate4sd3_1 hold841 (.A(_00761_),
    .X(net3101));
 sg13g2_dlygate4sd3_1 hold842 (.A(\i_peripherals.func_sel[42] ),
    .X(net3102));
 sg13g2_dlygate4sd3_1 hold843 (.A(_00541_),
    .X(net3103));
 sg13g2_dlygate4sd3_1 hold844 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[0] ),
    .X(net3104));
 sg13g2_dlygate4sd3_1 hold845 (.A(_00350_),
    .X(net3105));
 sg13g2_dlygate4sd3_1 hold846 (.A(\i_tinyqv.cpu.instr_data[2][13] ),
    .X(net3106));
 sg13g2_dlygate4sd3_1 hold847 (.A(_00749_),
    .X(net3107));
 sg13g2_dlygate4sd3_1 hold848 (.A(\i_peripherals.i_user_peri39._GEN[111] ),
    .X(net3108));
 sg13g2_dlygate4sd3_1 hold849 (.A(_00244_),
    .X(net3109));
 sg13g2_dlygate4sd3_1 hold850 (.A(\i_tinyqv.cpu.i_core.mie[4] ),
    .X(net3110));
 sg13g2_dlygate4sd3_1 hold851 (.A(\i_peripherals.i_user_peri39._GEN[64] ),
    .X(net3111));
 sg13g2_dlygate4sd3_1 hold852 (.A(_00755_),
    .X(net3112));
 sg13g2_dlygate4sd3_1 hold853 (.A(\i_tinyqv.cpu.instr_data[2][1] ),
    .X(net3113));
 sg13g2_dlygate4sd3_1 hold854 (.A(_00657_),
    .X(net3114));
 sg13g2_dlygate4sd3_1 hold855 (.A(\i_tinyqv.cpu.instr_data[2][7] ),
    .X(net3115));
 sg13g2_dlygate4sd3_1 hold856 (.A(_00743_),
    .X(net3116));
 sg13g2_dlygate4sd3_1 hold857 (.A(\i_tinyqv.cpu.instr_data[0][11] ),
    .X(net3117));
 sg13g2_dlygate4sd3_1 hold858 (.A(_00466_),
    .X(net3118));
 sg13g2_dlygate4sd3_1 hold859 (.A(\i_tinyqv.cpu.instr_data[0][4] ),
    .X(net3119));
 sg13g2_dlygate4sd3_1 hold860 (.A(\i_tinyqv.cpu.instr_data[1][9] ),
    .X(net3120));
 sg13g2_dlygate4sd3_1 hold861 (.A(_00085_),
    .X(net3121));
 sg13g2_dlygate4sd3_1 hold862 (.A(\i_tinyqv.cpu.i_core.mip[1] ),
    .X(net3122));
 sg13g2_dlygate4sd3_1 hold863 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[7] ),
    .X(net3123));
 sg13g2_dlygate4sd3_1 hold864 (.A(\i_peripherals.i_user_peri39._GEN[3] ),
    .X(net3124));
 sg13g2_dlygate4sd3_1 hold865 (.A(_00232_),
    .X(net3125));
 sg13g2_dlygate4sd3_1 hold866 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[1] ),
    .X(net3126));
 sg13g2_dlygate4sd3_1 hold867 (.A(\i_tinyqv.cpu.instr_data[1][7] ),
    .X(net3127));
 sg13g2_dlygate4sd3_1 hold868 (.A(_00083_),
    .X(net3128));
 sg13g2_dlygate4sd3_1 hold869 (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[0] ),
    .X(net3129));
 sg13g2_dlygate4sd3_1 hold870 (.A(_00121_),
    .X(net3130));
 sg13g2_dlygate4sd3_1 hold871 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[1] ),
    .X(net3131));
 sg13g2_dlygate4sd3_1 hold872 (.A(_00723_),
    .X(net3132));
 sg13g2_dlygate4sd3_1 hold873 (.A(\i_tinyqv.cpu.imm[29] ),
    .X(net3133));
 sg13g2_dlygate4sd3_1 hold874 (.A(\i_peripherals.i_user_peri39._GEN[94] ),
    .X(net3134));
 sg13g2_dlygate4sd3_1 hold875 (.A(_00785_),
    .X(net3135));
 sg13g2_dlygate4sd3_1 hold876 (.A(\i_peripherals.gpio_out[4] ),
    .X(net3136));
 sg13g2_dlygate4sd3_1 hold877 (.A(_00375_),
    .X(net3137));
 sg13g2_dlygate4sd3_1 hold878 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[2] ),
    .X(net3138));
 sg13g2_dlygate4sd3_1 hold879 (.A(_00724_),
    .X(net3139));
 sg13g2_dlygate4sd3_1 hold880 (.A(\i_tinyqv.cpu.i_core.last_interrupt_req[1] ),
    .X(net3140));
 sg13g2_dlygate4sd3_1 hold881 (.A(_00122_),
    .X(net3141));
 sg13g2_dlygate4sd3_1 hold882 (.A(\i_tinyqv.cpu.instr_data[1][11] ),
    .X(net3142));
 sg13g2_dlygate4sd3_1 hold883 (.A(_00087_),
    .X(net3143));
 sg13g2_dlygate4sd3_1 hold884 (.A(\i_peripherals.i_uart.uart_rx_buf_data[1] ),
    .X(net3144));
 sg13g2_dlygate4sd3_1 hold885 (.A(\i_tinyqv.cpu.instr_data[0][9] ),
    .X(net3145));
 sg13g2_dlygate4sd3_1 hold886 (.A(_00464_),
    .X(net3146));
 sg13g2_dlygate4sd3_1 hold887 (.A(\i_tinyqv.cpu.instr_data[0][13] ),
    .X(net3147));
 sg13g2_dlygate4sd3_1 hold888 (.A(_00468_),
    .X(net3148));
 sg13g2_dlygate4sd3_1 hold889 (.A(\i_tinyqv.mem.q_ctrl.addr[4] ),
    .X(net3149));
 sg13g2_dlygate4sd3_1 hold890 (.A(\i_peripherals.i_user_peri39._GEN[118] ),
    .X(net3150));
 sg13g2_dlygate4sd3_1 hold891 (.A(_00251_),
    .X(net3151));
 sg13g2_dlygate4sd3_1 hold892 (.A(\i_peripherals.i_user_peri39._GEN[38] ),
    .X(net3152));
 sg13g2_dlygate4sd3_1 hold893 (.A(_00267_),
    .X(net3153));
 sg13g2_dlygate4sd3_1 hold894 (.A(\addr[21] ),
    .X(net3154));
 sg13g2_dlygate4sd3_1 hold895 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[0] ),
    .X(net3155));
 sg13g2_dlygate4sd3_1 hold896 (.A(_00722_),
    .X(net3156));
 sg13g2_dlygate4sd3_1 hold897 (.A(\i_tinyqv.cpu.instr_data[2][4] ),
    .X(net3157));
 sg13g2_dlygate4sd3_1 hold898 (.A(\i_peripherals.i_user_peri39._GEN[68] ),
    .X(net3158));
 sg13g2_dlygate4sd3_1 hold899 (.A(_00759_),
    .X(net3159));
 sg13g2_dlygate4sd3_1 hold900 (.A(\i_tinyqv.cpu.instr_data[0][14] ),
    .X(net3160));
 sg13g2_dlygate4sd3_1 hold901 (.A(_05897_),
    .X(net3161));
 sg13g2_dlygate4sd3_1 hold902 (.A(_00469_),
    .X(net3162));
 sg13g2_dlygate4sd3_1 hold903 (.A(\addr[1] ),
    .X(net3163));
 sg13g2_dlygate4sd3_1 hold904 (.A(\i_tinyqv.mem.q_ctrl.addr[5] ),
    .X(net3164));
 sg13g2_dlygate4sd3_1 hold905 (.A(_00635_),
    .X(net3165));
 sg13g2_dlygate4sd3_1 hold906 (.A(\i_tinyqv.cpu.instr_data[3][0] ),
    .X(net3166));
 sg13g2_dlygate4sd3_1 hold907 (.A(_00295_),
    .X(net3167));
 sg13g2_dlygate4sd3_1 hold908 (.A(\addr[18] ),
    .X(net3168));
 sg13g2_dlygate4sd3_1 hold909 (.A(_00866_),
    .X(net3169));
 sg13g2_dlygate4sd3_1 hold910 (.A(\i_tinyqv.mem.q_ctrl.spi_in_buffer[3] ),
    .X(net3170));
 sg13g2_dlygate4sd3_1 hold911 (.A(_00725_),
    .X(net3171));
 sg13g2_dlygate4sd3_1 hold912 (.A(\addr[14] ),
    .X(net3172));
 sg13g2_dlygate4sd3_1 hold913 (.A(_00862_),
    .X(net3173));
 sg13g2_dlygate4sd3_1 hold914 (.A(\i_tinyqv.mem.q_ctrl.addr[7] ),
    .X(net3174));
 sg13g2_dlygate4sd3_1 hold915 (.A(_00637_),
    .X(net3175));
 sg13g2_dlygate4sd3_1 hold916 (.A(\addr[13] ),
    .X(net3176));
 sg13g2_dlygate4sd3_1 hold917 (.A(_00861_),
    .X(net3177));
 sg13g2_dlygate4sd3_1 hold918 (.A(\i_peripherals.i_uart.uart_rx_buf_data[5] ),
    .X(net3178));
 sg13g2_dlygate4sd3_1 hold919 (.A(_00355_),
    .X(net3179));
 sg13g2_dlygate4sd3_1 hold920 (.A(\i_peripherals.i_user_peri39._GEN[66] ),
    .X(net3180));
 sg13g2_dlygate4sd3_1 hold921 (.A(_00757_),
    .X(net3181));
 sg13g2_dlygate4sd3_1 hold922 (.A(\i_debug_uart_tx.fsm_state[1] ),
    .X(net3182));
 sg13g2_dlygate4sd3_1 hold923 (.A(_05807_),
    .X(net3183));
 sg13g2_dlygate4sd3_1 hold924 (.A(_00433_),
    .X(net3184));
 sg13g2_dlygate4sd3_1 hold925 (.A(\i_tinyqv.cpu.i_core.mcause[3] ),
    .X(net3185));
 sg13g2_dlygate4sd3_1 hold926 (.A(_02699_),
    .X(net3186));
 sg13g2_dlygate4sd3_1 hold927 (.A(\i_peripherals.gpio_out[6] ),
    .X(net3187));
 sg13g2_dlygate4sd3_1 hold928 (.A(_00377_),
    .X(net3188));
 sg13g2_dlygate4sd3_1 hold929 (.A(\i_tinyqv.cpu.i_core.mcause[4] ),
    .X(net3189));
 sg13g2_dlygate4sd3_1 hold930 (.A(_02700_),
    .X(net3190));
 sg13g2_dlygate4sd3_1 hold931 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[6] ),
    .X(net3191));
 sg13g2_dlygate4sd3_1 hold932 (.A(_05497_),
    .X(net3192));
 sg13g2_dlygate4sd3_1 hold933 (.A(_00364_),
    .X(net3193));
 sg13g2_dlygate4sd3_1 hold934 (.A(\i_peripherals.data_out[5] ),
    .X(net3194));
 sg13g2_dlygate4sd3_1 hold935 (.A(_05601_),
    .X(net3195));
 sg13g2_dlygate4sd3_1 hold936 (.A(\data_to_write[25] ),
    .X(net3196));
 sg13g2_dlygate4sd3_1 hold937 (.A(\addr[19] ),
    .X(net3197));
 sg13g2_dlygate4sd3_1 hold938 (.A(_00867_),
    .X(net3198));
 sg13g2_dlygate4sd3_1 hold939 (.A(\i_tinyqv.mem.q_ctrl.addr[1] ),
    .X(net3199));
 sg13g2_dlygate4sd3_1 hold940 (.A(_00297_),
    .X(net3200));
 sg13g2_dlygate4sd3_1 hold941 (.A(\i_debug_uart_tx.cycle_counter[0] ),
    .X(net3201));
 sg13g2_dlygate4sd3_1 hold942 (.A(_05794_),
    .X(net3202));
 sg13g2_dlygate4sd3_1 hold943 (.A(\i_debug_uart_tx.cycle_counter[1] ),
    .X(net3203));
 sg13g2_dlygate4sd3_1 hold944 (.A(\i_peripherals.data_out[15] ),
    .X(net3204));
 sg13g2_dlygate4sd3_1 hold945 (.A(_05674_),
    .X(net3205));
 sg13g2_dlygate4sd3_1 hold946 (.A(\i_peripherals.i_user_peri39._GEN[121] ),
    .X(net3206));
 sg13g2_dlygate4sd3_1 hold947 (.A(\i_tinyqv.cpu.instr_data[1][4] ),
    .X(net3207));
 sg13g2_dlygate4sd3_1 hold948 (.A(\i_tinyqv.mem.q_ctrl.addr[9] ),
    .X(net3208));
 sg13g2_dlygate4sd3_1 hold949 (.A(_00639_),
    .X(net3209));
 sg13g2_dlygate4sd3_1 hold950 (.A(\i_tinyqv.cpu.instr_data[2][9] ),
    .X(net3210));
 sg13g2_dlygate4sd3_1 hold951 (.A(_00745_),
    .X(net3211));
 sg13g2_dlygate4sd3_1 hold952 (.A(\i_tinyqv.mem.q_ctrl.addr[3] ),
    .X(net3212));
 sg13g2_dlygate4sd3_1 hold953 (.A(_05305_),
    .X(net3213));
 sg13g2_dlygate4sd3_1 hold954 (.A(_00299_),
    .X(net3214));
 sg13g2_dlygate4sd3_1 hold955 (.A(\i_peripherals.func_sel[18] ),
    .X(net3215));
 sg13g2_dlygate4sd3_1 hold956 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[0] ),
    .X(net3216));
 sg13g2_dlygate4sd3_1 hold957 (.A(_05381_),
    .X(net3217));
 sg13g2_dlygate4sd3_1 hold958 (.A(_00319_),
    .X(net3218));
 sg13g2_dlygate4sd3_1 hold959 (.A(\addr[17] ),
    .X(net3219));
 sg13g2_dlygate4sd3_1 hold960 (.A(_00865_),
    .X(net3220));
 sg13g2_dlygate4sd3_1 hold961 (.A(\i_peripherals.data_out[21] ),
    .X(net3221));
 sg13g2_dlygate4sd3_1 hold962 (.A(_05704_),
    .X(net3222));
 sg13g2_dlygate4sd3_1 hold963 (.A(\i_tinyqv.cpu.instr_data[2][0] ),
    .X(net3223));
 sg13g2_dlygate4sd3_1 hold964 (.A(_00656_),
    .X(net3224));
 sg13g2_dlygate4sd3_1 hold965 (.A(\data_to_write[24] ),
    .X(net3225));
 sg13g2_dlygate4sd3_1 hold966 (.A(\i_peripherals.data_out[17] ),
    .X(net3226));
 sg13g2_dlygate4sd3_1 hold967 (.A(_05684_),
    .X(net3227));
 sg13g2_dlygate4sd3_1 hold968 (.A(\i_peripherals.func_sel[30] ),
    .X(net3228));
 sg13g2_dlygate4sd3_1 hold969 (.A(\data_to_write[28] ),
    .X(net3229));
 sg13g2_dlygate4sd3_1 hold970 (.A(\i_tinyqv.cpu.instr_data[2][10] ),
    .X(net3230));
 sg13g2_dlygate4sd3_1 hold971 (.A(_00746_),
    .X(net3231));
 sg13g2_dlygate4sd3_1 hold972 (.A(\i_tinyqv.cpu.instr_data[0][8] ),
    .X(net3232));
 sg13g2_dlygate4sd3_1 hold973 (.A(_00463_),
    .X(net3233));
 sg13g2_dlygate4sd3_1 hold974 (.A(\i_peripherals.data_out[31] ),
    .X(net3234));
 sg13g2_dlygate4sd3_1 hold975 (.A(_05758_),
    .X(net3235));
 sg13g2_dlygate4sd3_1 hold976 (.A(\i_tinyqv.cpu.i_core.mie[8] ),
    .X(net3236));
 sg13g2_dlygate4sd3_1 hold977 (.A(\addr[15] ),
    .X(net3237));
 sg13g2_dlygate4sd3_1 hold978 (.A(_00863_),
    .X(net3238));
 sg13g2_dlygate4sd3_1 hold979 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[2] ),
    .X(net3239));
 sg13g2_dlygate4sd3_1 hold980 (.A(_00710_),
    .X(net3240));
 sg13g2_dlygate4sd3_1 hold981 (.A(\i_peripherals.i_user_peri39._GEN[71] ),
    .X(net3241));
 sg13g2_dlygate4sd3_1 hold982 (.A(_00762_),
    .X(net3242));
 sg13g2_dlygate4sd3_1 hold983 (.A(\i_peripherals.data_out[13] ),
    .X(net3243));
 sg13g2_dlygate4sd3_1 hold984 (.A(_05663_),
    .X(net3244));
 sg13g2_dlygate4sd3_1 hold985 (.A(\i_tinyqv.cpu.instr_data_in[0] ),
    .X(net3245));
 sg13g2_dlygate4sd3_1 hold986 (.A(_00668_),
    .X(net3246));
 sg13g2_dlygate4sd3_1 hold987 (.A(\i_peripherals.i_uart.uart_rx_buf_data[4] ),
    .X(net3247));
 sg13g2_dlygate4sd3_1 hold988 (.A(_00354_),
    .X(net3248));
 sg13g2_dlygate4sd3_1 hold989 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[5] ),
    .X(net3249));
 sg13g2_dlygate4sd3_1 hold990 (.A(_05391_),
    .X(net3250));
 sg13g2_dlygate4sd3_1 hold991 (.A(_00324_),
    .X(net3251));
 sg13g2_dlygate4sd3_1 hold992 (.A(\i_peripherals.i_uart.uart_rx_buf_data[2] ),
    .X(net3252));
 sg13g2_dlygate4sd3_1 hold993 (.A(_00352_),
    .X(net3253));
 sg13g2_dlygate4sd3_1 hold994 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[3] ),
    .X(net3254));
 sg13g2_dlygate4sd3_1 hold995 (.A(_00096_),
    .X(net3255));
 sg13g2_dlygate4sd3_1 hold996 (.A(\i_peripherals.data_out[25] ),
    .X(net3256));
 sg13g2_dlygate4sd3_1 hold997 (.A(_05725_),
    .X(net3257));
 sg13g2_dlygate4sd3_1 hold998 (.A(\i_peripherals.data_out[22] ),
    .X(net3258));
 sg13g2_dlygate4sd3_1 hold999 (.A(_05709_),
    .X(net3259));
 sg13g2_dlygate4sd3_1 hold1000 (.A(\i_peripherals.data_out[14] ),
    .X(net3260));
 sg13g2_dlygate4sd3_1 hold1001 (.A(_05669_),
    .X(net3261));
 sg13g2_dlygate4sd3_1 hold1002 (.A(\i_peripherals.i_user_peri39._GEN[67] ),
    .X(net3262));
 sg13g2_dlygate4sd3_1 hold1003 (.A(_00758_),
    .X(net3263));
 sg13g2_dlygate4sd3_1 hold1004 (.A(\i_peripherals.gpio_out[5] ),
    .X(net3264));
 sg13g2_dlygate4sd3_1 hold1005 (.A(_00376_),
    .X(net3265));
 sg13g2_dlygate4sd3_1 hold1006 (.A(\i_peripherals.gpio_out[3] ),
    .X(net3266));
 sg13g2_dlygate4sd3_1 hold1007 (.A(_00374_),
    .X(net3267));
 sg13g2_dlygate4sd3_1 hold1008 (.A(\i_peripherals.func_sel[24] ),
    .X(net3268));
 sg13g2_dlygate4sd3_1 hold1009 (.A(\i_peripherals.data_out[26] ),
    .X(net3269));
 sg13g2_dlygate4sd3_1 hold1010 (.A(_05730_),
    .X(net3270));
 sg13g2_dlygate4sd3_1 hold1011 (.A(\i_peripherals.data_out[1] ),
    .X(net3271));
 sg13g2_dlygate4sd3_1 hold1012 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[9] ),
    .X(net3272));
 sg13g2_dlygate4sd3_1 hold1013 (.A(_05399_),
    .X(net3273));
 sg13g2_dlygate4sd3_1 hold1014 (.A(_00328_),
    .X(net3274));
 sg13g2_dlygate4sd3_1 hold1015 (.A(\i_tinyqv.cpu.i_core.mepc[13] ),
    .X(net3275));
 sg13g2_dlygate4sd3_1 hold1016 (.A(_00498_),
    .X(net3276));
 sg13g2_dlygate4sd3_1 hold1017 (.A(\i_peripherals.func_sel[7] ),
    .X(net3277));
 sg13g2_dlygate4sd3_1 hold1018 (.A(_00578_),
    .X(net3278));
 sg13g2_dlygate4sd3_1 hold1019 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[1] ),
    .X(net3279));
 sg13g2_dlygate4sd3_1 hold1020 (.A(_00714_),
    .X(net3280));
 sg13g2_dlygate4sd3_1 hold1021 (.A(\data_to_write[31] ),
    .X(net3281));
 sg13g2_dlygate4sd3_1 hold1022 (.A(\i_peripherals.data_out[27] ),
    .X(net3282));
 sg13g2_dlygate4sd3_1 hold1023 (.A(_05736_),
    .X(net3283));
 sg13g2_dlygate4sd3_1 hold1024 (.A(\i_peripherals.data_out[18] ),
    .X(net3284));
 sg13g2_dlygate4sd3_1 hold1025 (.A(_05689_),
    .X(net3285));
 sg13g2_dlygate4sd3_1 hold1026 (.A(\i_peripherals.data_out[20] ),
    .X(net3286));
 sg13g2_dlygate4sd3_1 hold1027 (.A(_05699_),
    .X(net3287));
 sg13g2_dlygate4sd3_1 hold1028 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[7] ),
    .X(net3288));
 sg13g2_dlygate4sd3_1 hold1029 (.A(_05395_),
    .X(net3289));
 sg13g2_dlygate4sd3_1 hold1030 (.A(_00326_),
    .X(net3290));
 sg13g2_dlygate4sd3_1 hold1031 (.A(\i_tinyqv.mem.q_ctrl.addr[2] ),
    .X(net3291));
 sg13g2_dlygate4sd3_1 hold1032 (.A(_05297_),
    .X(net3292));
 sg13g2_dlygate4sd3_1 hold1033 (.A(_00298_),
    .X(net3293));
 sg13g2_dlygate4sd3_1 hold1034 (.A(\i_debug_uart_tx.data_to_send[1] ),
    .X(net3294));
 sg13g2_dlygate4sd3_1 hold1035 (.A(_05768_),
    .X(net3295));
 sg13g2_dlygate4sd3_1 hold1036 (.A(_00419_),
    .X(net3296));
 sg13g2_dlygate4sd3_1 hold1037 (.A(\i_peripherals.i_uart.uart_rx_buf_data[3] ),
    .X(net3297));
 sg13g2_dlygate4sd3_1 hold1038 (.A(_00353_),
    .X(net3298));
 sg13g2_dlygate4sd3_1 hold1039 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[2] ),
    .X(net3299));
 sg13g2_dlygate4sd3_1 hold1040 (.A(_00313_),
    .X(net3300));
 sg13g2_dlygate4sd3_1 hold1041 (.A(\i_peripherals.data_out[19] ),
    .X(net3301));
 sg13g2_dlygate4sd3_1 hold1042 (.A(_05694_),
    .X(net3302));
 sg13g2_dlygate4sd3_1 hold1043 (.A(\i_tinyqv.mem.q_ctrl.addr[22] ),
    .X(net3303));
 sg13g2_dlygate4sd3_1 hold1044 (.A(_00652_),
    .X(net3304));
 sg13g2_dlygate4sd3_1 hold1045 (.A(\i_peripherals.data_out[30] ),
    .X(net3305));
 sg13g2_dlygate4sd3_1 hold1046 (.A(_05753_),
    .X(net3306));
 sg13g2_dlygate4sd3_1 hold1047 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[8] ),
    .X(net3307));
 sg13g2_dlygate4sd3_1 hold1048 (.A(_05397_),
    .X(net3308));
 sg13g2_dlygate4sd3_1 hold1049 (.A(\addr[20] ),
    .X(net3309));
 sg13g2_dlygate4sd3_1 hold1050 (.A(\i_tinyqv.cpu.i_core.mie[0] ),
    .X(net3310));
 sg13g2_dlygate4sd3_1 hold1051 (.A(\i_tinyqv.cpu.i_core.i_shift.b[3] ),
    .X(net3311));
 sg13g2_dlygate4sd3_1 hold1052 (.A(_00488_),
    .X(net3312));
 sg13g2_dlygate4sd3_1 hold1053 (.A(\i_peripherals.data_out[16] ),
    .X(net3313));
 sg13g2_dlygate4sd3_1 hold1054 (.A(_05679_),
    .X(net3314));
 sg13g2_dlygate4sd3_1 hold1055 (.A(\i_peripherals.data_out[23] ),
    .X(net3315));
 sg13g2_dlygate4sd3_1 hold1056 (.A(_05714_),
    .X(net3316));
 sg13g2_dlygate4sd3_1 hold1057 (.A(\data_to_write[29] ),
    .X(net3317));
 sg13g2_dlygate4sd3_1 hold1058 (.A(\i_tinyqv.mem.q_ctrl.addr[23] ),
    .X(net3318));
 sg13g2_dlygate4sd3_1 hold1059 (.A(_06484_),
    .X(net3319));
 sg13g2_dlygate4sd3_1 hold1060 (.A(_00653_),
    .X(net3320));
 sg13g2_dlygate4sd3_1 hold1061 (.A(\i_tinyqv.mem.qspi_data_buf[28] ),
    .X(net3321));
 sg13g2_dlygate4sd3_1 hold1062 (.A(_00696_),
    .X(net3322));
 sg13g2_dlygate4sd3_1 hold1063 (.A(\i_peripherals.data_out[28] ),
    .X(net3323));
 sg13g2_dlygate4sd3_1 hold1064 (.A(_05741_),
    .X(net3324));
 sg13g2_dlygate4sd3_1 hold1065 (.A(\i_tinyqv.cpu.i_core.mepc[6] ),
    .X(net3325));
 sg13g2_dlygate4sd3_1 hold1066 (.A(_00491_),
    .X(net3326));
 sg13g2_dlygate4sd3_1 hold1067 (.A(\data_to_write[30] ),
    .X(net3327));
 sg13g2_dlygate4sd3_1 hold1068 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[30] ),
    .X(net3328));
 sg13g2_dlygate4sd3_1 hold1069 (.A(\data_to_write[26] ),
    .X(net3329));
 sg13g2_dlygate4sd3_1 hold1070 (.A(_00222_),
    .X(net3330));
 sg13g2_dlygate4sd3_1 hold1071 (.A(\i_peripherals.data_out_hold ),
    .X(net3331));
 sg13g2_dlygate4sd3_1 hold1072 (.A(_05760_),
    .X(net3332));
 sg13g2_dlygate4sd3_1 hold1073 (.A(\i_peripherals.data_out[7] ),
    .X(net3333));
 sg13g2_dlygate4sd3_1 hold1074 (.A(_05622_),
    .X(net3334));
 sg13g2_dlygate4sd3_1 hold1075 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[6] ),
    .X(net3335));
 sg13g2_dlygate4sd3_1 hold1076 (.A(_05393_),
    .X(net3336));
 sg13g2_dlygate4sd3_1 hold1077 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[1] ),
    .X(net3337));
 sg13g2_dlygate4sd3_1 hold1078 (.A(\i_tinyqv.cpu.i_core.mepc[19] ),
    .X(net3338));
 sg13g2_dlygate4sd3_1 hold1079 (.A(\i_tinyqv.cpu.i_core.mepc[16] ),
    .X(net3339));
 sg13g2_dlygate4sd3_1 hold1080 (.A(_00501_),
    .X(net3340));
 sg13g2_dlygate4sd3_1 hold1081 (.A(\i_peripherals.i_user_peri39.instr[25] ),
    .X(net3341));
 sg13g2_dlygate4sd3_1 hold1082 (.A(\i_tinyqv.mem.qspi_data_buf[24] ),
    .X(net3342));
 sg13g2_dlygate4sd3_1 hold1083 (.A(_00692_),
    .X(net3343));
 sg13g2_dlygate4sd3_1 hold1084 (.A(\i_tinyqv.cpu.i_core.mepc[14] ),
    .X(net3344));
 sg13g2_dlygate4sd3_1 hold1085 (.A(_00499_),
    .X(net3345));
 sg13g2_dlygate4sd3_1 hold1086 (.A(\i_tinyqv.cpu.instr_data[1][5] ),
    .X(net3346));
 sg13g2_dlygate4sd3_1 hold1087 (.A(_00081_),
    .X(net3347));
 sg13g2_dlygate4sd3_1 hold1088 (.A(\i_peripherals.func_sel[39] ),
    .X(net3348));
 sg13g2_dlygate4sd3_1 hold1089 (.A(_00550_),
    .X(net3349));
 sg13g2_dlygate4sd3_1 hold1090 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[4] ),
    .X(net3350));
 sg13g2_dlygate4sd3_1 hold1091 (.A(_05389_),
    .X(net3351));
 sg13g2_dlygate4sd3_1 hold1092 (.A(\i_peripherals.data_out[8] ),
    .X(net3352));
 sg13g2_dlygate4sd3_1 hold1093 (.A(_00393_),
    .X(net3353));
 sg13g2_dlygate4sd3_1 hold1094 (.A(\i_debug_uart_tx.cycle_counter[2] ),
    .X(net3354));
 sg13g2_dlygate4sd3_1 hold1095 (.A(\i_tinyqv.cpu.i_core.mepc[17] ),
    .X(net3355));
 sg13g2_dlygate4sd3_1 hold1096 (.A(\i_peripherals.i_uart.uart_rx_buf_data[7] ),
    .X(net3356));
 sg13g2_dlygate4sd3_1 hold1097 (.A(\i_tinyqv.cpu.i_core.mepc[7] ),
    .X(net3357));
 sg13g2_dlygate4sd3_1 hold1098 (.A(_00496_),
    .X(net3358));
 sg13g2_dlygate4sd3_1 hold1099 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[3] ),
    .X(net3359));
 sg13g2_dlygate4sd3_1 hold1100 (.A(_00338_),
    .X(net3360));
 sg13g2_dlygate4sd3_1 hold1101 (.A(\i_tinyqv.cpu.instr_data[3][6] ),
    .X(net3361));
 sg13g2_dlygate4sd3_1 hold1102 (.A(_00475_),
    .X(net3362));
 sg13g2_dlygate4sd3_1 hold1103 (.A(\i_tinyqv.cpu.instr_data[0][6] ),
    .X(net3363));
 sg13g2_dlygate4sd3_1 hold1104 (.A(_00461_),
    .X(net3364));
 sg13g2_dlygate4sd3_1 hold1105 (.A(\i_debug_uart_tx.fsm_state[3] ),
    .X(net3365));
 sg13g2_dlygate4sd3_1 hold1106 (.A(_05811_),
    .X(net3366));
 sg13g2_dlygate4sd3_1 hold1107 (.A(_00435_),
    .X(net3367));
 sg13g2_dlygate4sd3_1 hold1108 (.A(\i_peripherals.data_out[24] ),
    .X(net3368));
 sg13g2_dlygate4sd3_1 hold1109 (.A(_05720_),
    .X(net3369));
 sg13g2_dlygate4sd3_1 hold1110 (.A(\i_peripherals.i_user_peri39.instr[14] ),
    .X(net3370));
 sg13g2_dlygate4sd3_1 hold1111 (.A(_00210_),
    .X(net3371));
 sg13g2_dlygate4sd3_1 hold1112 (.A(\i_peripherals.i_user_peri39.instr[29] ),
    .X(net3372));
 sg13g2_dlygate4sd3_1 hold1113 (.A(\i_tinyqv.cpu.instr_data[1][10] ),
    .X(net3373));
 sg13g2_dlygate4sd3_1 hold1114 (.A(_00086_),
    .X(net3374));
 sg13g2_dlygate4sd3_1 hold1115 (.A(\i_peripherals.i_user_peri39.instr[28] ),
    .X(net3375));
 sg13g2_dlygate4sd3_1 hold1116 (.A(\addr[10] ),
    .X(net3376));
 sg13g2_dlygate4sd3_1 hold1117 (.A(_00858_),
    .X(net3377));
 sg13g2_dlygate4sd3_1 hold1118 (.A(\i_peripherals.func_sel[45] ),
    .X(net3378));
 sg13g2_dlygate4sd3_1 hold1119 (.A(_00544_),
    .X(net3379));
 sg13g2_dlygate4sd3_1 hold1120 (.A(\i_tinyqv.mem.q_ctrl.spi_clk_use_neg ),
    .X(net3380));
 sg13g2_dlygate4sd3_1 hold1121 (.A(\i_peripherals.i_user_peri39.instr[31] ),
    .X(net3381));
 sg13g2_dlygate4sd3_1 hold1122 (.A(\i_tinyqv.cpu.i_core.mepc[10] ),
    .X(net3382));
 sg13g2_dlygate4sd3_1 hold1123 (.A(\i_tinyqv.cpu.instr_data[1][15] ),
    .X(net3383));
 sg13g2_dlygate4sd3_1 hold1124 (.A(_00091_),
    .X(net3384));
 sg13g2_dlygate4sd3_1 hold1125 (.A(\i_tinyqv.mem.qspi_data_buf[31] ),
    .X(net3385));
 sg13g2_dlygate4sd3_1 hold1126 (.A(\data_to_write[27] ),
    .X(net3386));
 sg13g2_dlygate4sd3_1 hold1127 (.A(\i_tinyqv.cpu.i_core.mepc[12] ),
    .X(net3387));
 sg13g2_dlygate4sd3_1 hold1128 (.A(_00497_),
    .X(net3388));
 sg13g2_dlygate4sd3_1 hold1129 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[5] ),
    .X(net3389));
 sg13g2_dlygate4sd3_1 hold1130 (.A(_00316_),
    .X(net3390));
 sg13g2_dlygate4sd3_1 hold1131 (.A(\i_tinyqv.cpu.instr_data[3][12] ),
    .X(net3391));
 sg13g2_dlygate4sd3_1 hold1132 (.A(_00481_),
    .X(net3392));
 sg13g2_dlygate4sd3_1 hold1133 (.A(\i_peripherals.i_user_peri39.instr[4] ),
    .X(net3393));
 sg13g2_dlygate4sd3_1 hold1134 (.A(_00200_),
    .X(net3394));
 sg13g2_dlygate4sd3_1 hold1135 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[31] ),
    .X(net3395));
 sg13g2_dlygate4sd3_1 hold1136 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[2] ),
    .X(net3396));
 sg13g2_dlygate4sd3_1 hold1137 (.A(\i_tinyqv.cpu.i_core.mepc[3] ),
    .X(net3397));
 sg13g2_dlygate4sd3_1 hold1138 (.A(\i_tinyqv.cpu.i_core.i_shift.a[24] ),
    .X(net3398));
 sg13g2_dlygate4sd3_1 hold1139 (.A(_00533_),
    .X(net3399));
 sg13g2_dlygate4sd3_1 hold1140 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[6] ),
    .X(net3400));
 sg13g2_dlygate4sd3_1 hold1141 (.A(_00317_),
    .X(net3401));
 sg13g2_dlygate4sd3_1 hold1142 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[10] ),
    .X(net3402));
 sg13g2_dlygate4sd3_1 hold1143 (.A(\i_tinyqv.cpu.i_core.mepc[15] ),
    .X(net3403));
 sg13g2_dlygate4sd3_1 hold1144 (.A(\i_tinyqv.cpu.instr_data[1][2] ),
    .X(net3404));
 sg13g2_dlygate4sd3_1 hold1145 (.A(_00078_),
    .X(net3405));
 sg13g2_dlygate4sd3_1 hold1146 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[6] ),
    .X(net3406));
 sg13g2_dlygate4sd3_1 hold1147 (.A(\i_tinyqv.cpu.instr_data[3][2] ),
    .X(net3407));
 sg13g2_dlygate4sd3_1 hold1148 (.A(_00471_),
    .X(net3408));
 sg13g2_dlygate4sd3_1 hold1149 (.A(\i_tinyqv.cpu.i_core.mip[0] ),
    .X(net3409));
 sg13g2_dlygate4sd3_1 hold1150 (.A(\i_tinyqv.cpu.instr_data[1][6] ),
    .X(net3410));
 sg13g2_dlygate4sd3_1 hold1151 (.A(_00082_),
    .X(net3411));
 sg13g2_dlygate4sd3_1 hold1152 (.A(\i_tinyqv.cpu.instr_data[0][15] ),
    .X(net3412));
 sg13g2_dlygate4sd3_1 hold1153 (.A(_00470_),
    .X(net3413));
 sg13g2_dlygate4sd3_1 hold1154 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[4] ),
    .X(net3414));
 sg13g2_dlygate4sd3_1 hold1155 (.A(\i_peripherals.i_uart.uart_rx_buf_data[6] ),
    .X(net3415));
 sg13g2_dlygate4sd3_1 hold1156 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[29] ),
    .X(net3416));
 sg13g2_dlygate4sd3_1 hold1157 (.A(\i_peripherals.func_sel[1] ),
    .X(net3417));
 sg13g2_dlygate4sd3_1 hold1158 (.A(_00380_),
    .X(net3418));
 sg13g2_dlygate4sd3_1 hold1159 (.A(\i_peripherals.data_out[4] ),
    .X(net3419));
 sg13g2_dlygate4sd3_1 hold1160 (.A(_05591_),
    .X(net3420));
 sg13g2_dlygate4sd3_1 hold1161 (.A(\i_tinyqv.cpu.instr_data[2][6] ),
    .X(net3421));
 sg13g2_dlygate4sd3_1 hold1162 (.A(_00742_),
    .X(net3422));
 sg13g2_dlygate4sd3_1 hold1163 (.A(\i_tinyqv.mem.q_ctrl.data_req ),
    .X(net3423));
 sg13g2_dlygate4sd3_1 hold1164 (.A(_00073_),
    .X(net3424));
 sg13g2_dlygate4sd3_1 hold1165 (.A(\i_tinyqv.mem.qspi_data_buf[26] ),
    .X(net3425));
 sg13g2_dlygate4sd3_1 hold1166 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[4] ),
    .X(net3426));
 sg13g2_dlygate4sd3_1 hold1167 (.A(_00340_),
    .X(net3427));
 sg13g2_dlygate4sd3_1 hold1168 (.A(\i_tinyqv.cpu.instr_data[2][12] ),
    .X(net3428));
 sg13g2_dlygate4sd3_1 hold1169 (.A(_00748_),
    .X(net3429));
 sg13g2_dlygate4sd3_1 hold1170 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[25] ),
    .X(net3430));
 sg13g2_dlygate4sd3_1 hold1171 (.A(\time_count[4] ),
    .X(net3431));
 sg13g2_dlygate4sd3_1 hold1172 (.A(_07234_),
    .X(net3432));
 sg13g2_dlygate4sd3_1 hold1173 (.A(\i_tinyqv.mem.qspi_data_buf[25] ),
    .X(net3433));
 sg13g2_dlygate4sd3_1 hold1174 (.A(_00693_),
    .X(net3434));
 sg13g2_dlygate4sd3_1 hold1175 (.A(\data_to_write[15] ),
    .X(net3435));
 sg13g2_dlygate4sd3_1 hold1176 (.A(_00211_),
    .X(net3436));
 sg13g2_dlygate4sd3_1 hold1177 (.A(\i_tinyqv.cpu.i_core.mepc[18] ),
    .X(net3437));
 sg13g2_dlygate4sd3_1 hold1178 (.A(\i_tinyqv.cpu.instr_data[2][8] ),
    .X(net3438));
 sg13g2_dlygate4sd3_1 hold1179 (.A(_00744_),
    .X(net3439));
 sg13g2_dlygate4sd3_1 hold1180 (.A(\i_tinyqv.cpu.instr_data[2][3] ),
    .X(net3440));
 sg13g2_dlygate4sd3_1 hold1181 (.A(_00739_),
    .X(net3441));
 sg13g2_dlygate4sd3_1 hold1182 (.A(\i_tinyqv.cpu.is_store ),
    .X(net3442));
 sg13g2_dlygate4sd3_1 hold1183 (.A(_01405_),
    .X(net3443));
 sg13g2_dlygate4sd3_1 hold1184 (.A(\addr[23] ),
    .X(net3444));
 sg13g2_dlygate4sd3_1 hold1185 (.A(_00871_),
    .X(net3445));
 sg13g2_dlygate4sd3_1 hold1186 (.A(\i_peripherals.i_user_peri39.instr[3] ),
    .X(net3446));
 sg13g2_dlygate4sd3_1 hold1187 (.A(_00199_),
    .X(net3447));
 sg13g2_dlygate4sd3_1 hold1188 (.A(\i_peripherals.i_uart.i_uart_rx.fsm_state[3] ),
    .X(net3448));
 sg13g2_dlygate4sd3_1 hold1189 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[1] ),
    .X(net3449));
 sg13g2_dlygate4sd3_1 hold1190 (.A(_00312_),
    .X(net3450));
 sg13g2_dlygate4sd3_1 hold1191 (.A(\i_peripherals.i_user_peri39.instr[24] ),
    .X(net3451));
 sg13g2_dlygate4sd3_1 hold1192 (.A(\i_tinyqv.cpu.instr_data[2][2] ),
    .X(net3452));
 sg13g2_dlygate4sd3_1 hold1193 (.A(_00738_),
    .X(net3453));
 sg13g2_dlygate4sd3_1 hold1194 (.A(\i_tinyqv.mem.qspi_data_buf[27] ),
    .X(net3454));
 sg13g2_dlygate4sd3_1 hold1195 (.A(_00695_),
    .X(net3455));
 sg13g2_dlygate4sd3_1 hold1196 (.A(\i_tinyqv.cpu.instr_data[1][3] ),
    .X(net3456));
 sg13g2_dlygate4sd3_1 hold1197 (.A(_00079_),
    .X(net3457));
 sg13g2_dlygate4sd3_1 hold1198 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[7] ),
    .X(net3458));
 sg13g2_dlygate4sd3_1 hold1199 (.A(_00318_),
    .X(net3459));
 sg13g2_dlygate4sd3_1 hold1200 (.A(\i_tinyqv.cpu.i_core.mie[7] ),
    .X(net3460));
 sg13g2_dlygate4sd3_1 hold1201 (.A(\i_tinyqv.cpu.instr_data[0][5] ),
    .X(net3461));
 sg13g2_dlygate4sd3_1 hold1202 (.A(_00460_),
    .X(net3462));
 sg13g2_dlygate4sd3_1 hold1203 (.A(\i_peripherals.i_user_peri39.instr[9] ),
    .X(net3463));
 sg13g2_dlygate4sd3_1 hold1204 (.A(_00205_),
    .X(net3464));
 sg13g2_dlygate4sd3_1 hold1205 (.A(\i_tinyqv.cpu.instr_data[0][2] ),
    .X(net3465));
 sg13g2_dlygate4sd3_1 hold1206 (.A(_00457_),
    .X(net3466));
 sg13g2_dlygate4sd3_1 hold1207 (.A(\i_peripherals.i_user_peri39.instr[27] ),
    .X(net3467));
 sg13g2_dlygate4sd3_1 hold1208 (.A(\i_tinyqv.cpu.i_core.mcause[1] ),
    .X(net3468));
 sg13g2_dlygate4sd3_1 hold1209 (.A(_00111_),
    .X(net3469));
 sg13g2_dlygate4sd3_1 hold1210 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[22] ),
    .X(net3470));
 sg13g2_dlygate4sd3_1 hold1211 (.A(\i_tinyqv.cpu.i_core.mie[11] ),
    .X(net3471));
 sg13g2_dlygate4sd3_1 hold1212 (.A(\i_debug_uart_tx.data_to_send[3] ),
    .X(net3472));
 sg13g2_dlygate4sd3_1 hold1213 (.A(_05778_),
    .X(net3473));
 sg13g2_dlygate4sd3_1 hold1214 (.A(\i_peripherals.data_out[6] ),
    .X(net3474));
 sg13g2_dlygate4sd3_1 hold1215 (.A(_00391_),
    .X(net3475));
 sg13g2_dlygate4sd3_1 hold1216 (.A(\i_tinyqv.cpu.i_core.is_interrupt ),
    .X(net3476));
 sg13g2_dlygate4sd3_1 hold1217 (.A(\i_peripherals.data_out[2] ),
    .X(net3477));
 sg13g2_dlygate4sd3_1 hold1218 (.A(_00387_),
    .X(net3478));
 sg13g2_dlygate4sd3_1 hold1219 (.A(\i_tinyqv.mem.q_ctrl.delay_cycles_cfg[1] ),
    .X(net3479));
 sg13g2_dlygate4sd3_1 hold1220 (.A(\data_to_write[17] ),
    .X(net3480));
 sg13g2_dlygate4sd3_1 hold1221 (.A(_00213_),
    .X(net3481));
 sg13g2_dlygate4sd3_1 hold1222 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[0] ),
    .X(net3482));
 sg13g2_dlygate4sd3_1 hold1223 (.A(_00708_),
    .X(net3483));
 sg13g2_dlygate4sd3_1 hold1224 (.A(\i_tinyqv.cpu.i_core.mie[15] ),
    .X(net3484));
 sg13g2_dlygate4sd3_1 hold1225 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[0] ),
    .X(net3485));
 sg13g2_dlygate4sd3_1 hold1226 (.A(\i_peripherals.i_uart.i_uart_rx.recieved_data[5] ),
    .X(net3486));
 sg13g2_dlygate4sd3_1 hold1227 (.A(\i_peripherals.i_user_peri39.instr[5] ),
    .X(net3487));
 sg13g2_dlygate4sd3_1 hold1228 (.A(\i_peripherals.i_user_peri39._GEN[76] ),
    .X(net3488));
 sg13g2_dlygate4sd3_1 hold1229 (.A(_00767_),
    .X(net3489));
 sg13g2_dlygate4sd3_1 hold1230 (.A(\i_tinyqv.cpu.instr_data[0][3] ),
    .X(net3490));
 sg13g2_dlygate4sd3_1 hold1231 (.A(_00458_),
    .X(net3491));
 sg13g2_dlygate4sd3_1 hold1232 (.A(\i_peripherals.i_user_peri39.instr[30] ),
    .X(net3492));
 sg13g2_dlygate4sd3_1 hold1233 (.A(\i_tinyqv.mem.data_from_read[23] ),
    .X(net3493));
 sg13g2_dlygate4sd3_1 hold1234 (.A(_00691_),
    .X(net3494));
 sg13g2_dlygate4sd3_1 hold1235 (.A(\i_tinyqv.cpu.instr_data[3][15] ),
    .X(net3495));
 sg13g2_dlygate4sd3_1 hold1236 (.A(_00484_),
    .X(net3496));
 sg13g2_dlygate4sd3_1 hold1237 (.A(\i_peripherals.func_sel[36] ),
    .X(net3497));
 sg13g2_dlygate4sd3_1 hold1238 (.A(\i_peripherals.i_user_peri39.math_result_reg[24] ),
    .X(net3498));
 sg13g2_dlygate4sd3_1 hold1239 (.A(\i_peripherals.func_sel[47] ),
    .X(net3499));
 sg13g2_dlygate4sd3_1 hold1240 (.A(\i_peripherals.i_user_peri39._GEN[75] ),
    .X(net3500));
 sg13g2_dlygate4sd3_1 hold1241 (.A(_00766_),
    .X(net3501));
 sg13g2_dlygate4sd3_1 hold1242 (.A(\i_peripherals.i_user_peri39.instr[1] ),
    .X(net3502));
 sg13g2_dlygate4sd3_1 hold1243 (.A(_00197_),
    .X(net3503));
 sg13g2_dlygate4sd3_1 hold1244 (.A(\i_peripherals.i_user_peri39.math_result_reg[5] ),
    .X(net3504));
 sg13g2_dlygate4sd3_1 hold1245 (.A(_00147_),
    .X(net3505));
 sg13g2_dlygate4sd3_1 hold1246 (.A(\time_count[5] ),
    .X(net3506));
 sg13g2_dlygate4sd3_1 hold1247 (.A(_07236_),
    .X(net3507));
 sg13g2_dlygate4sd3_1 hold1248 (.A(\i_tinyqv.mem.q_ctrl.spi_data_oe[0] ),
    .X(net3508));
 sg13g2_dlygate4sd3_1 hold1249 (.A(_06685_),
    .X(net3509));
 sg13g2_dlygate4sd3_1 hold1250 (.A(_00719_),
    .X(net3510));
 sg13g2_dlygate4sd3_1 hold1251 (.A(\i_peripherals.i_user_peri39.instr[7] ),
    .X(net3511));
 sg13g2_dlygate4sd3_1 hold1252 (.A(_00203_),
    .X(net3512));
 sg13g2_dlygate4sd3_1 hold1253 (.A(\i_tinyqv.cpu.i_core.mepc[11] ),
    .X(net3513));
 sg13g2_dlygate4sd3_1 hold1254 (.A(\i_peripherals.i_user_peri39._GEN[84] ),
    .X(net3514));
 sg13g2_dlygate4sd3_1 hold1255 (.A(_00775_),
    .X(net3515));
 sg13g2_dlygate4sd3_1 hold1256 (.A(\i_tinyqv.mem.q_ctrl.last_ram_b_sel ),
    .X(net3516));
 sg13g2_dlygate4sd3_1 hold1257 (.A(_06680_),
    .X(net3517));
 sg13g2_dlygate4sd3_1 hold1258 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[4] ),
    .X(net3518));
 sg13g2_dlygate4sd3_1 hold1259 (.A(_05495_),
    .X(net3519));
 sg13g2_dlygate4sd3_1 hold1260 (.A(_00362_),
    .X(net3520));
 sg13g2_dlygate4sd3_1 hold1261 (.A(\i_tinyqv.cpu.instr_data[2][5] ),
    .X(net3521));
 sg13g2_dlygate4sd3_1 hold1262 (.A(_00741_),
    .X(net3522));
 sg13g2_dlygate4sd3_1 hold1263 (.A(\i_tinyqv.mem.q_ctrl.addr[14] ),
    .X(net3523));
 sg13g2_dlygate4sd3_1 hold1264 (.A(_00644_),
    .X(net3524));
 sg13g2_dlygate4sd3_1 hold1265 (.A(\i_tinyqv.cpu.instr_data[3][8] ),
    .X(net3525));
 sg13g2_dlygate4sd3_1 hold1266 (.A(_00477_),
    .X(net3526));
 sg13g2_dlygate4sd3_1 hold1267 (.A(\i_tinyqv.cpu.instr_data[1][8] ),
    .X(net3527));
 sg13g2_dlygate4sd3_1 hold1268 (.A(_00084_),
    .X(net3528));
 sg13g2_dlygate4sd3_1 hold1269 (.A(\i_peripherals.func_sel[41] ),
    .X(net3529));
 sg13g2_dlygate4sd3_1 hold1270 (.A(\i_peripherals.i_user_peri39._GEN[72] ),
    .X(net3530));
 sg13g2_dlygate4sd3_1 hold1271 (.A(_00763_),
    .X(net3531));
 sg13g2_dlygate4sd3_1 hold1272 (.A(\i_peripherals.i_uart.i_uart_tx.fsm_state[2] ),
    .X(net3532));
 sg13g2_dlygate4sd3_1 hold1273 (.A(_05412_),
    .X(net3533));
 sg13g2_dlygate4sd3_1 hold1274 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[8] ),
    .X(net3534));
 sg13g2_dlygate4sd3_1 hold1275 (.A(_05502_),
    .X(net3535));
 sg13g2_dlygate4sd3_1 hold1276 (.A(\i_tinyqv.mem.q_ctrl.addr[16] ),
    .X(net3536));
 sg13g2_dlygate4sd3_1 hold1277 (.A(_00646_),
    .X(net3537));
 sg13g2_dlygate4sd3_1 hold1278 (.A(\i_tinyqv.cpu.i_core.i_shift.a[12] ),
    .X(net3538));
 sg13g2_dlygate4sd3_1 hold1279 (.A(_00521_),
    .X(net3539));
 sg13g2_dlygate4sd3_1 hold1280 (.A(\i_tinyqv.cpu.i_core.i_shift.a[4] ),
    .X(net3540));
 sg13g2_dlygate4sd3_1 hold1281 (.A(_00509_),
    .X(net3541));
 sg13g2_dlygate4sd3_1 hold1282 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][0] ),
    .X(net3542));
 sg13g2_dlygate4sd3_1 hold1283 (.A(\i_tinyqv.mem.q_ctrl.addr[19] ),
    .X(net3543));
 sg13g2_dlygate4sd3_1 hold1284 (.A(_00649_),
    .X(net3544));
 sg13g2_dlygate4sd3_1 hold1285 (.A(\i_debug_uart_tx.data_to_send[2] ),
    .X(net3545));
 sg13g2_dlygate4sd3_1 hold1286 (.A(_00420_),
    .X(net3546));
 sg13g2_dlygate4sd3_1 hold1287 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[3] ),
    .X(net3547));
 sg13g2_dlygate4sd3_1 hold1288 (.A(_00314_),
    .X(net3548));
 sg13g2_dlygate4sd3_1 hold1289 (.A(\i_peripherals.i_user_peri39.instr[6] ),
    .X(net3549));
 sg13g2_dlygate4sd3_1 hold1290 (.A(_00202_),
    .X(net3550));
 sg13g2_dlygate4sd3_1 hold1291 (.A(\i_peripherals.func_sel[43] ),
    .X(net3551));
 sg13g2_dlygate4sd3_1 hold1292 (.A(_00542_),
    .X(net3552));
 sg13g2_dlygate4sd3_1 hold1293 (.A(\i_debug_uart_tx.cycle_counter[3] ),
    .X(net3553));
 sg13g2_dlygate4sd3_1 hold1294 (.A(\i_tinyqv.cpu.instr_data_in[1] ),
    .X(net3554));
 sg13g2_dlygate4sd3_1 hold1295 (.A(_00669_),
    .X(net3555));
 sg13g2_dlygate4sd3_1 hold1296 (.A(\i_peripherals.i_user_peri39._GEN[42] ),
    .X(net3556));
 sg13g2_dlygate4sd3_1 hold1297 (.A(_00271_),
    .X(net3557));
 sg13g2_dlygate4sd3_1 hold1298 (.A(\i_tinyqv.cpu.instr_len[1] ),
    .X(net3558));
 sg13g2_dlygate4sd3_1 hold1299 (.A(\i_peripherals.i_user_peri39._GEN[107] ),
    .X(net3559));
 sg13g2_dlygate4sd3_1 hold1300 (.A(_00240_),
    .X(net3560));
 sg13g2_dlygate4sd3_1 hold1301 (.A(\i_tinyqv.mem.q_ctrl.addr[6] ),
    .X(net3561));
 sg13g2_dlygate4sd3_1 hold1302 (.A(_00636_),
    .X(net3562));
 sg13g2_dlygate4sd3_1 hold1303 (.A(\i_peripherals.i_user_peri39._GEN[106] ),
    .X(net3563));
 sg13g2_dlygate4sd3_1 hold1304 (.A(_00239_),
    .X(net3564));
 sg13g2_dlygate4sd3_1 hold1305 (.A(\i_tinyqv.cpu.i_core.mepc[9] ),
    .X(net3565));
 sg13g2_dlygate4sd3_1 hold1306 (.A(_00494_),
    .X(net3566));
 sg13g2_dlygate4sd3_1 hold1307 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][1] ),
    .X(net3567));
 sg13g2_dlygate4sd3_1 hold1308 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[3] ),
    .X(net3568));
 sg13g2_dlygate4sd3_1 hold1309 (.A(_05493_),
    .X(net3569));
 sg13g2_dlygate4sd3_1 hold1310 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][2] ),
    .X(net3570));
 sg13g2_dlygate4sd3_1 hold1311 (.A(\i_tinyqv.cpu.instr_data[3][3] ),
    .X(net3571));
 sg13g2_dlygate4sd3_1 hold1312 (.A(_00472_),
    .X(net3572));
 sg13g2_dlygate4sd3_1 hold1313 (.A(\i_peripherals.data_out[3] ),
    .X(net3573));
 sg13g2_dlygate4sd3_1 hold1314 (.A(_05581_),
    .X(net3574));
 sg13g2_dlygate4sd3_1 hold1315 (.A(\i_tinyqv.cpu.i_core.i_shift.b[4] ),
    .X(net3575));
 sg13g2_dlygate4sd3_1 hold1316 (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .X(net3576));
 sg13g2_dlygate4sd3_1 hold1317 (.A(_02673_),
    .X(net3577));
 sg13g2_dlygate4sd3_1 hold1318 (.A(_00105_),
    .X(net3578));
 sg13g2_dlygate4sd3_1 hold1319 (.A(\i_tinyqv.cpu.i_core.mepc[4] ),
    .X(net3579));
 sg13g2_dlygate4sd3_1 hold1320 (.A(_00489_),
    .X(net3580));
 sg13g2_dlygate4sd3_1 hold1321 (.A(\i_tinyqv.cpu.i_core.mepc[8] ),
    .X(net3581));
 sg13g2_dlygate4sd3_1 hold1322 (.A(\i_peripherals.i_user_peri39._GEN[73] ),
    .X(net3582));
 sg13g2_dlygate4sd3_1 hold1323 (.A(_00764_),
    .X(net3583));
 sg13g2_dlygate4sd3_1 hold1324 (.A(\i_peripherals.i_user_peri39._GEN[104] ),
    .X(net3584));
 sg13g2_dlygate4sd3_1 hold1325 (.A(_00237_),
    .X(net3585));
 sg13g2_dlygate4sd3_1 hold1326 (.A(\i_peripherals.i_user_peri39.instr[2] ),
    .X(net3586));
 sg13g2_dlygate4sd3_1 hold1327 (.A(_00198_),
    .X(net3587));
 sg13g2_dlygate4sd3_1 hold1328 (.A(\i_peripherals.i_user_peri39._GEN[43] ),
    .X(net3588));
 sg13g2_dlygate4sd3_1 hold1329 (.A(_00272_),
    .X(net3589));
 sg13g2_dlygate4sd3_1 hold1330 (.A(\data_to_write[13] ),
    .X(net3590));
 sg13g2_dlygate4sd3_1 hold1331 (.A(\data_to_write[23] ),
    .X(net3591));
 sg13g2_dlygate4sd3_1 hold1332 (.A(_00219_),
    .X(net3592));
 sg13g2_dlygate4sd3_1 hold1333 (.A(\i_tinyqv.mem.data_from_read[22] ),
    .X(net3593));
 sg13g2_dlygate4sd3_1 hold1334 (.A(_00690_),
    .X(net3594));
 sg13g2_dlygate4sd3_1 hold1335 (.A(\i_tinyqv.cpu.counter[2] ),
    .X(net3595));
 sg13g2_dlygate4sd3_1 hold1336 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][0] ),
    .X(net3596));
 sg13g2_dlygate4sd3_1 hold1337 (.A(\i_tinyqv.cpu.instr_data[0][12] ),
    .X(net3597));
 sg13g2_dlygate4sd3_1 hold1338 (.A(_00467_),
    .X(net3598));
 sg13g2_dlygate4sd3_1 hold1339 (.A(\i_tinyqv.mem.q_ctrl.addr[8] ),
    .X(net3599));
 sg13g2_dlygate4sd3_1 hold1340 (.A(_00638_),
    .X(net3600));
 sg13g2_dlygate4sd3_1 hold1341 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[1] ),
    .X(net3601));
 sg13g2_dlygate4sd3_1 hold1342 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[5] ),
    .X(net3602));
 sg13g2_dlygate4sd3_1 hold1343 (.A(\i_tinyqv.mem.q_ctrl.addr[12] ),
    .X(net3603));
 sg13g2_dlygate4sd3_1 hold1344 (.A(\i_tinyqv.mem.q_ctrl.addr[10] ),
    .X(net3604));
 sg13g2_dlygate4sd3_1 hold1345 (.A(\i_peripherals.data_out[10] ),
    .X(net3605));
 sg13g2_dlygate4sd3_1 hold1346 (.A(_00395_),
    .X(net3606));
 sg13g2_dlygate4sd3_1 hold1347 (.A(\data_to_write[18] ),
    .X(net3607));
 sg13g2_dlygate4sd3_1 hold1348 (.A(_00214_),
    .X(net3608));
 sg13g2_dlygate4sd3_1 hold1349 (.A(\i_peripherals.i_user_peri39._GEN[40] ),
    .X(net3609));
 sg13g2_dlygate4sd3_1 hold1350 (.A(_00269_),
    .X(net3610));
 sg13g2_dlygate4sd3_1 hold1351 (.A(\i_tinyqv.mem.qspi_data_buf[29] ),
    .X(net3611));
 sg13g2_dlygate4sd3_1 hold1352 (.A(_00697_),
    .X(net3612));
 sg13g2_dlygate4sd3_1 hold1353 (.A(\i_tinyqv.mem.data_from_read[21] ),
    .X(net3613));
 sg13g2_dlygate4sd3_1 hold1354 (.A(_00689_),
    .X(net3614));
 sg13g2_dlygate4sd3_1 hold1355 (.A(\i_tinyqv.cpu.i_core.i_shift.a[14] ),
    .X(net3615));
 sg13g2_dlygate4sd3_1 hold1356 (.A(_00523_),
    .X(net3616));
 sg13g2_dlygate4sd3_1 hold1357 (.A(\i_peripherals.func_sel[12] ),
    .X(net3617));
 sg13g2_dlygate4sd3_1 hold1358 (.A(_00571_),
    .X(net3618));
 sg13g2_dlygate4sd3_1 hold1359 (.A(\i_peripherals.data_out[29] ),
    .X(net3619));
 sg13g2_dlygate4sd3_1 hold1360 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][0] ),
    .X(net3620));
 sg13g2_dlygate4sd3_1 hold1361 (.A(\i_tinyqv.cpu.imm[23] ),
    .X(net3621));
 sg13g2_dlygate4sd3_1 hold1362 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][0] ),
    .X(net3622));
 sg13g2_dlygate4sd3_1 hold1363 (.A(\i_tinyqv.cpu.instr_data[1][12] ),
    .X(net3623));
 sg13g2_dlygate4sd3_1 hold1364 (.A(_00088_),
    .X(net3624));
 sg13g2_dlygate4sd3_1 hold1365 (.A(\i_peripherals.data_out[0] ),
    .X(net3625));
 sg13g2_dlygate4sd3_1 hold1366 (.A(_00385_),
    .X(net3626));
 sg13g2_dlygate4sd3_1 hold1367 (.A(\i_tinyqv.cpu.i_core.mie[13] ),
    .X(net3627));
 sg13g2_dlygate4sd3_1 hold1368 (.A(\i_tinyqv.cpu.i_core.i_cycles.rstn ),
    .X(net3628));
 sg13g2_dlygate4sd3_1 hold1369 (.A(\i_tinyqv.mem.qspi_data_buf[14] ),
    .X(net3629));
 sg13g2_dlygate4sd3_1 hold1370 (.A(_00682_),
    .X(net3630));
 sg13g2_dlygate4sd3_1 hold1371 (.A(\i_tinyqv.cpu.imm[31] ),
    .X(net3631));
 sg13g2_dlygate4sd3_1 hold1372 (.A(\i_peripherals.i_user_peri39.instr[13] ),
    .X(net3632));
 sg13g2_dlygate4sd3_1 hold1373 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][3] ),
    .X(net3633));
 sg13g2_dlygate4sd3_1 hold1374 (.A(\i_peripherals.i_user_peri39._GEN[108] ),
    .X(net3634));
 sg13g2_dlygate4sd3_1 hold1375 (.A(_00241_),
    .X(net3635));
 sg13g2_dlygate4sd3_1 hold1376 (.A(\i_tinyqv.cpu.instr_data_in[3] ),
    .X(net3636));
 sg13g2_dlygate4sd3_1 hold1377 (.A(_00671_),
    .X(net3637));
 sg13g2_dlygate4sd3_1 hold1378 (.A(\i_tinyqv.cpu.i_core.i_shift.a[15] ),
    .X(net3638));
 sg13g2_dlygate4sd3_1 hold1379 (.A(_00524_),
    .X(net3639));
 sg13g2_dlygate4sd3_1 hold1380 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][1] ),
    .X(net3640));
 sg13g2_dlygate4sd3_1 hold1381 (.A(_00046_),
    .X(net3641));
 sg13g2_dlygate4sd3_1 hold1382 (.A(\data_to_write[21] ),
    .X(net3642));
 sg13g2_dlygate4sd3_1 hold1383 (.A(\data_to_write[22] ),
    .X(net3643));
 sg13g2_dlygate4sd3_1 hold1384 (.A(_00218_),
    .X(net3644));
 sg13g2_dlygate4sd3_1 hold1385 (.A(\i_tinyqv.cpu.i_core.i_shift.a[11] ),
    .X(net3645));
 sg13g2_dlygate4sd3_1 hold1386 (.A(\i_tinyqv.mem.continue_txn ),
    .X(net3646));
 sg13g2_dlygate4sd3_1 hold1387 (.A(_00665_),
    .X(net3647));
 sg13g2_dlygate4sd3_1 hold1388 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[11] ),
    .X(net3648));
 sg13g2_dlygate4sd3_1 hold1389 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[3] ),
    .X(net3649));
 sg13g2_dlygate4sd3_1 hold1390 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][0] ),
    .X(net3650));
 sg13g2_dlygate4sd3_1 hold1391 (.A(\i_tinyqv.cpu.i_core.i_shift.a[28] ),
    .X(net3651));
 sg13g2_dlygate4sd3_1 hold1392 (.A(\i_tinyqv.cpu.is_branch ),
    .X(net3652));
 sg13g2_dlygate4sd3_1 hold1393 (.A(\i_tinyqv.cpu.instr_data[3][5] ),
    .X(net3653));
 sg13g2_dlygate4sd3_1 hold1394 (.A(_00474_),
    .X(net3654));
 sg13g2_dlygate4sd3_1 hold1395 (.A(\i_tinyqv.mem.q_ctrl.addr[18] ),
    .X(net3655));
 sg13g2_dlygate4sd3_1 hold1396 (.A(\i_tinyqv.mem.q_ctrl.addr[11] ),
    .X(net3656));
 sg13g2_dlygate4sd3_1 hold1397 (.A(_00641_),
    .X(net3657));
 sg13g2_dlygate4sd3_1 hold1398 (.A(\i_tinyqv.cpu.i_core.imm_lo[0] ),
    .X(net3658));
 sg13g2_dlygate4sd3_1 hold1399 (.A(\i_tinyqv.mem.qspi_data_buf[30] ),
    .X(net3659));
 sg13g2_dlygate4sd3_1 hold1400 (.A(_00698_),
    .X(net3660));
 sg13g2_dlygate4sd3_1 hold1401 (.A(\i_peripherals.i_user_peri39.math_result_reg[22] ),
    .X(net3661));
 sg13g2_dlygate4sd3_1 hold1402 (.A(\i_peripherals.i_user_peri39.math_result_reg[12] ),
    .X(net3662));
 sg13g2_dlygate4sd3_1 hold1403 (.A(_00154_),
    .X(net3663));
 sg13g2_dlygate4sd3_1 hold1404 (.A(\i_tinyqv.mem.qspi_data_buf[15] ),
    .X(net3664));
 sg13g2_dlygate4sd3_1 hold1405 (.A(\i_tinyqv.cpu.i_core.mie[14] ),
    .X(net3665));
 sg13g2_dlygate4sd3_1 hold1406 (.A(\addr[6] ),
    .X(net3666));
 sg13g2_dlygate4sd3_1 hold1407 (.A(_00854_),
    .X(net3667));
 sg13g2_dlygate4sd3_1 hold1408 (.A(\i_peripherals.i_user_peri39._GEN[44] ),
    .X(net3668));
 sg13g2_dlygate4sd3_1 hold1409 (.A(_00273_),
    .X(net3669));
 sg13g2_dlygate4sd3_1 hold1410 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][2] ),
    .X(net3670));
 sg13g2_dlygate4sd3_1 hold1411 (.A(\i_debug_uart_tx.data_to_send[4] ),
    .X(net3671));
 sg13g2_dlygate4sd3_1 hold1412 (.A(\i_peripherals.i_user_peri39._GEN[74] ),
    .X(net3672));
 sg13g2_dlygate4sd3_1 hold1413 (.A(_00765_),
    .X(net3673));
 sg13g2_dlygate4sd3_1 hold1414 (.A(\data_to_write[16] ),
    .X(net3674));
 sg13g2_dlygate4sd3_1 hold1415 (.A(_00212_),
    .X(net3675));
 sg13g2_dlygate4sd3_1 hold1416 (.A(\i_tinyqv.cpu.i_core.time_hi[0] ),
    .X(net3676));
 sg13g2_dlygate4sd3_1 hold1417 (.A(_02680_),
    .X(net3677));
 sg13g2_dlygate4sd3_1 hold1418 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][1] ),
    .X(net3678));
 sg13g2_dlygate4sd3_1 hold1419 (.A(\i_peripherals.i_user_peri39.math_result_reg[8] ),
    .X(net3679));
 sg13g2_dlygate4sd3_1 hold1420 (.A(_00150_),
    .X(net3680));
 sg13g2_dlygate4sd3_1 hold1421 (.A(\i_tinyqv.cpu.counter[4] ),
    .X(net3681));
 sg13g2_dlygate4sd3_1 hold1422 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][1] ),
    .X(net3682));
 sg13g2_dlygate4sd3_1 hold1423 (.A(\i_peripherals.i_user_peri39._GEN[116] ),
    .X(net3683));
 sg13g2_dlygate4sd3_1 hold1424 (.A(_00249_),
    .X(net3684));
 sg13g2_dlygate4sd3_1 hold1425 (.A(\i_tinyqv.mem.q_ctrl.addr[21] ),
    .X(net3685));
 sg13g2_dlygate4sd3_1 hold1426 (.A(\i_tinyqv.cpu.i_core.i_shift.a[13] ),
    .X(net3686));
 sg13g2_dlygate4sd3_1 hold1427 (.A(_00522_),
    .X(net3687));
 sg13g2_dlygate4sd3_1 hold1428 (.A(\data_to_write[14] ),
    .X(net3688));
 sg13g2_dlygate4sd3_1 hold1429 (.A(\i_tinyqv.cpu.data_ready_latch ),
    .X(net3689));
 sg13g2_dlygate4sd3_1 hold1430 (.A(\i_peripherals.i_uart.baud_divider[8] ),
    .X(net3690));
 sg13g2_dlygate4sd3_1 hold1431 (.A(_00583_),
    .X(net3691));
 sg13g2_dlygate4sd3_1 hold1432 (.A(\i_peripherals.i_user_peri39.math_result_reg[6] ),
    .X(net3692));
 sg13g2_dlygate4sd3_1 hold1433 (.A(_00148_),
    .X(net3693));
 sg13g2_dlygate4sd3_1 hold1434 (.A(\i_debug_uart_tx.data_to_send[0] ),
    .X(net3694));
 sg13g2_dlygate4sd3_1 hold1435 (.A(_05761_),
    .X(net3695));
 sg13g2_dlygate4sd3_1 hold1436 (.A(_00418_),
    .X(net3696));
 sg13g2_dlygate4sd3_1 hold1437 (.A(\i_tinyqv.cpu.i_core.i_shift.a[29] ),
    .X(net3697));
 sg13g2_dlygate4sd3_1 hold1438 (.A(\i_peripherals.i_user_peri39.instr[21] ),
    .X(net3698));
 sg13g2_dlygate4sd3_1 hold1439 (.A(\i_tinyqv.cpu.mem_op_increment_reg ),
    .X(net3699));
 sg13g2_dlygate4sd3_1 hold1440 (.A(\i_tinyqv.cpu.is_auipc ),
    .X(net3700));
 sg13g2_dlygate4sd3_1 hold1441 (.A(\time_count[6] ),
    .X(net3701));
 sg13g2_dlygate4sd3_1 hold1442 (.A(\i_peripherals.i_user_peri39.busy_counter[1] ),
    .X(net3702));
 sg13g2_dlygate4sd3_1 hold1443 (.A(_00294_),
    .X(net3703));
 sg13g2_dlygate4sd3_1 hold1444 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[27] ),
    .X(net3704));
 sg13g2_dlygate4sd3_1 hold1445 (.A(_06016_),
    .X(net3705));
 sg13g2_dlygate4sd3_1 hold1446 (.A(_00594_),
    .X(net3706));
 sg13g2_dlygate4sd3_1 hold1447 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[1] ),
    .X(net3707));
 sg13g2_dlygate4sd3_1 hold1448 (.A(_06632_),
    .X(net3708));
 sg13g2_dlygate4sd3_1 hold1449 (.A(_00706_),
    .X(net3709));
 sg13g2_dlygate4sd3_1 hold1450 (.A(\i_tinyqv.cpu.i_core.mie[5] ),
    .X(net3710));
 sg13g2_dlygate4sd3_1 hold1451 (.A(\i_tinyqv.cpu.instr_data[2][15] ),
    .X(net3711));
 sg13g2_dlygate4sd3_1 hold1452 (.A(_00751_),
    .X(net3712));
 sg13g2_dlygate4sd3_1 hold1453 (.A(\i_tinyqv.cpu.no_write_in_progress ),
    .X(net3713));
 sg13g2_dlygate4sd3_1 hold1454 (.A(\i_peripherals.i_user_peri39.math_result_reg[30] ),
    .X(net3714));
 sg13g2_dlygate4sd3_1 hold1455 (.A(_00172_),
    .X(net3715));
 sg13g2_dlygate4sd3_1 hold1456 (.A(\i_peripherals.i_user_peri39.math_result_reg[27] ),
    .X(net3716));
 sg13g2_dlygate4sd3_1 hold1457 (.A(\i_peripherals.i_user_peri39.math_result_reg[21] ),
    .X(net3717));
 sg13g2_dlygate4sd3_1 hold1458 (.A(_00163_),
    .X(net3718));
 sg13g2_dlygate4sd3_1 hold1459 (.A(\i_tinyqv.cpu.i_core.i_shift.a[7] ),
    .X(net3719));
 sg13g2_dlygate4sd3_1 hold1460 (.A(_00512_),
    .X(net3720));
 sg13g2_dlygate4sd3_1 hold1461 (.A(\i_tinyqv.cpu.i_core.i_shift.a[16] ),
    .X(net3721));
 sg13g2_dlygate4sd3_1 hold1462 (.A(_00525_),
    .X(net3722));
 sg13g2_dlygate4sd3_1 hold1463 (.A(\i_peripherals.func_sel[46] ),
    .X(net3723));
 sg13g2_dlygate4sd3_1 hold1464 (.A(_00545_),
    .X(net3724));
 sg13g2_dlygate4sd3_1 hold1465 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[12][3] ),
    .X(net3725));
 sg13g2_dlygate4sd3_1 hold1466 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][0] ),
    .X(net3726));
 sg13g2_dlygate4sd3_1 hold1467 (.A(\i_peripherals.i_uart.baud_divider[10] ),
    .X(net3727));
 sg13g2_dlygate4sd3_1 hold1468 (.A(_00585_),
    .X(net3728));
 sg13g2_dlygate4sd3_1 hold1469 (.A(\i_tinyqv.cpu.i_core.cycle_count[2] ),
    .X(net3729));
 sg13g2_dlygate4sd3_1 hold1470 (.A(_02656_),
    .X(net3730));
 sg13g2_dlygate4sd3_1 hold1471 (.A(_00094_),
    .X(net3731));
 sg13g2_dlygate4sd3_1 hold1472 (.A(\i_tinyqv.cpu.data_ready_sync ),
    .X(net3732));
 sg13g2_dlygate4sd3_1 hold1473 (.A(\i_peripherals.i_user_peri39.math_result_reg[11] ),
    .X(net3733));
 sg13g2_dlygate4sd3_1 hold1474 (.A(_00153_),
    .X(net3734));
 sg13g2_dlygate4sd3_1 hold1475 (.A(\i_peripherals.i_user_peri39._GEN[52] ),
    .X(net3735));
 sg13g2_dlygate4sd3_1 hold1476 (.A(_00281_),
    .X(net3736));
 sg13g2_dlygate4sd3_1 hold1477 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][0] ),
    .X(net3737));
 sg13g2_dlygate4sd3_1 hold1478 (.A(\i_peripherals.data_out[9] ),
    .X(net3738));
 sg13g2_dlygate4sd3_1 hold1479 (.A(_00394_),
    .X(net3739));
 sg13g2_dlygate4sd3_1 hold1480 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[11] ),
    .X(net3740));
 sg13g2_dlygate4sd3_1 hold1481 (.A(_05507_),
    .X(net3741));
 sg13g2_dlygate4sd3_1 hold1482 (.A(\i_tinyqv.mem.q_ctrl.addr[20] ),
    .X(net3742));
 sg13g2_dlygate4sd3_1 hold1483 (.A(\i_peripherals.i_user_peri39.math_result_reg[2] ),
    .X(net3743));
 sg13g2_dlygate4sd3_1 hold1484 (.A(_00144_),
    .X(net3744));
 sg13g2_dlygate4sd3_1 hold1485 (.A(\i_peripherals.i_user_peri39.math_result_reg[23] ),
    .X(net3745));
 sg13g2_dlygate4sd3_1 hold1486 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][3] ),
    .X(net3746));
 sg13g2_dlygate4sd3_1 hold1487 (.A(\i_peripherals.i_user_peri39.instr[20] ),
    .X(net3747));
 sg13g2_dlygate4sd3_1 hold1488 (.A(_00216_),
    .X(net3748));
 sg13g2_dlygate4sd3_1 hold1489 (.A(\i_peripherals.i_user_peri39.math_result_reg[0] ),
    .X(net3749));
 sg13g2_dlygate4sd3_1 hold1490 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[9] ),
    .X(net3750));
 sg13g2_dlygate4sd3_1 hold1491 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[7] ),
    .X(net3751));
 sg13g2_dlygate4sd3_1 hold1492 (.A(_05499_),
    .X(net3752));
 sg13g2_dlygate4sd3_1 hold1493 (.A(\i_tinyqv.mem.q_ctrl.spi_clk_pos ),
    .X(net3753));
 sg13g2_dlygate4sd3_1 hold1494 (.A(_00707_),
    .X(net3754));
 sg13g2_dlygate4sd3_1 hold1495 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][1] ),
    .X(net3755));
 sg13g2_dlygate4sd3_1 hold1496 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[2] ),
    .X(net3756));
 sg13g2_dlygate4sd3_1 hold1497 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][1] ),
    .X(net3757));
 sg13g2_dlygate4sd3_1 hold1498 (.A(\i_peripherals.i_uart.i_uart_tx.fsm_state[0] ),
    .X(net3758));
 sg13g2_dlygate4sd3_1 hold1499 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[26] ),
    .X(net3759));
 sg13g2_dlygate4sd3_1 hold1500 (.A(\i_tinyqv.cpu.i_timer.i_mtime.data[1] ),
    .X(net3760));
 sg13g2_dlygate4sd3_1 hold1501 (.A(_02839_),
    .X(net3761));
 sg13g2_dlygate4sd3_1 hold1502 (.A(_00134_),
    .X(net3762));
 sg13g2_dlygate4sd3_1 hold1503 (.A(\i_peripherals.i_uart.i_uart_tx.data_to_send[0] ),
    .X(net3763));
 sg13g2_dlygate4sd3_1 hold1504 (.A(_00311_),
    .X(net3764));
 sg13g2_dlygate4sd3_1 hold1505 (.A(\i_tinyqv.cpu.i_core.mepc[5] ),
    .X(net3765));
 sg13g2_dlygate4sd3_1 hold1506 (.A(_00490_),
    .X(net3766));
 sg13g2_dlygate4sd3_1 hold1507 (.A(\i_tinyqv.cpu.is_jal ),
    .X(net3767));
 sg13g2_dlygate4sd3_1 hold1508 (.A(\i_peripherals.i_user_peri39.math_result_reg[19] ),
    .X(net3768));
 sg13g2_dlygate4sd3_1 hold1509 (.A(_00161_),
    .X(net3769));
 sg13g2_dlygate4sd3_1 hold1510 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[9] ),
    .X(net3770));
 sg13g2_dlygate4sd3_1 hold1511 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][2] ),
    .X(net3771));
 sg13g2_dlygate4sd3_1 hold1512 (.A(\data_to_write[19] ),
    .X(net3772));
 sg13g2_dlygate4sd3_1 hold1513 (.A(_00215_),
    .X(net3773));
 sg13g2_dlygate4sd3_1 hold1514 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[15] ),
    .X(net3774));
 sg13g2_dlygate4sd3_1 hold1515 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[1] ),
    .X(net3775));
 sg13g2_dlygate4sd3_1 hold1516 (.A(\i_peripherals.func_sel[44] ),
    .X(net3776));
 sg13g2_dlygate4sd3_1 hold1517 (.A(_00543_),
    .X(net3777));
 sg13g2_dlygate4sd3_1 hold1518 (.A(\i_tinyqv.mem.q_ctrl.addr[15] ),
    .X(net3778));
 sg13g2_dlygate4sd3_1 hold1519 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[6][3] ),
    .X(net3779));
 sg13g2_dlygate4sd3_1 hold1520 (.A(\i_tinyqv.cpu.i_core.mcause[0] ),
    .X(net3780));
 sg13g2_dlygate4sd3_1 hold1521 (.A(_00110_),
    .X(net3781));
 sg13g2_dlygate4sd3_1 hold1522 (.A(\time_limit[6] ),
    .X(net3782));
 sg13g2_dlygate4sd3_1 hold1523 (.A(_00006_),
    .X(net3783));
 sg13g2_dlygate4sd3_1 hold1524 (.A(\i_peripherals.i_uart.baud_divider[12] ),
    .X(net3784));
 sg13g2_dlygate4sd3_1 hold1525 (.A(_00587_),
    .X(net3785));
 sg13g2_dlygate4sd3_1 hold1526 (.A(\i_tinyqv.cpu.i_core.i_shift.a[19] ),
    .X(net3786));
 sg13g2_dlygate4sd3_1 hold1527 (.A(_00528_),
    .X(net3787));
 sg13g2_dlygate4sd3_1 hold1528 (.A(\i_tinyqv.cpu.imm[22] ),
    .X(net3788));
 sg13g2_dlygate4sd3_1 hold1529 (.A(\addr[24] ),
    .X(net3789));
 sg13g2_dlygate4sd3_1 hold1530 (.A(\i_peripherals.i_user_peri39.math_result_reg[20] ),
    .X(net3790));
 sg13g2_dlygate4sd3_1 hold1531 (.A(_00162_),
    .X(net3791));
 sg13g2_dlygate4sd3_1 hold1532 (.A(\i_tinyqv.mem.q_ctrl.read_cycles_count[0] ),
    .X(net3792));
 sg13g2_dlygate4sd3_1 hold1533 (.A(_00705_),
    .X(net3793));
 sg13g2_dlygate4sd3_1 hold1534 (.A(\i_peripherals.i_user_peri39.math_result_reg[15] ),
    .X(net3794));
 sg13g2_dlygate4sd3_1 hold1535 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[14][1] ),
    .X(net3795));
 sg13g2_dlygate4sd3_1 hold1536 (.A(\i_debug_uart_tx.data_to_send[5] ),
    .X(net3796));
 sg13g2_dlygate4sd3_1 hold1537 (.A(_00423_),
    .X(net3797));
 sg13g2_dlygate4sd3_1 hold1538 (.A(\i_tinyqv.cpu.data_read_n[0] ),
    .X(net3798));
 sg13g2_dlygate4sd3_1 hold1539 (.A(_00844_),
    .X(net3799));
 sg13g2_dlygate4sd3_1 hold1540 (.A(\i_tinyqv.cpu.data_read_n[1] ),
    .X(net3800));
 sg13g2_dlygate4sd3_1 hold1541 (.A(_00845_),
    .X(net3801));
 sg13g2_dlygate4sd3_1 hold1542 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][0] ),
    .X(net3802));
 sg13g2_dlygate4sd3_1 hold1543 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[6] ),
    .X(net3803));
 sg13g2_dlygate4sd3_1 hold1544 (.A(_00180_),
    .X(net3804));
 sg13g2_dlygate4sd3_1 hold1545 (.A(\i_tinyqv.cpu.i_core.mie[12] ),
    .X(net3805));
 sg13g2_dlygate4sd3_1 hold1546 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][3] ),
    .X(net3806));
 sg13g2_dlygate4sd3_1 hold1547 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[20] ),
    .X(net3807));
 sg13g2_dlygate4sd3_1 hold1548 (.A(\i_tinyqv.cpu.i_core.mie[3] ),
    .X(net3808));
 sg13g2_dlygate4sd3_1 hold1549 (.A(\i_tinyqv.cpu.i_core.mie[6] ),
    .X(net3809));
 sg13g2_dlygate4sd3_1 hold1550 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[10] ),
    .X(net3810));
 sg13g2_dlygate4sd3_1 hold1551 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[7] ),
    .X(net3811));
 sg13g2_dlygate4sd3_1 hold1552 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[19] ),
    .X(net3812));
 sg13g2_dlygate4sd3_1 hold1553 (.A(\i_tinyqv.cpu.i_core.i_shift.a[20] ),
    .X(net3813));
 sg13g2_dlygate4sd3_1 hold1554 (.A(\i_tinyqv.mem.q_ctrl.nibbles_remaining[1] ),
    .X(net3814));
 sg13g2_dlygate4sd3_1 hold1555 (.A(_00709_),
    .X(net3815));
 sg13g2_dlygate4sd3_1 hold1556 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][2] ),
    .X(net3816));
 sg13g2_dlygate4sd3_1 hold1557 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][2] ),
    .X(net3817));
 sg13g2_dlygate4sd3_1 hold1558 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][1] ),
    .X(net3818));
 sg13g2_dlygate4sd3_1 hold1559 (.A(\i_tinyqv.cpu.instr_len[2] ),
    .X(net3819));
 sg13g2_dlygate4sd3_1 hold1560 (.A(\i_tinyqv.cpu.instr_data_start[15] ),
    .X(net3820));
 sg13g2_dlygate4sd3_1 hold1561 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[18] ),
    .X(net3821));
 sg13g2_dlygate4sd3_1 hold1562 (.A(\i_peripherals.data_out[11] ),
    .X(net3822));
 sg13g2_dlygate4sd3_1 hold1563 (.A(_00396_),
    .X(net3823));
 sg13g2_dlygate4sd3_1 hold1564 (.A(\i_tinyqv.cpu.is_lui ),
    .X(net3824));
 sg13g2_dlygate4sd3_1 hold1565 (.A(\i_tinyqv.cpu.is_alu_imm ),
    .X(net3825));
 sg13g2_dlygate4sd3_1 hold1566 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][2] ),
    .X(net3826));
 sg13g2_dlygate4sd3_1 hold1567 (.A(\addr[7] ),
    .X(net3827));
 sg13g2_dlygate4sd3_1 hold1568 (.A(_00855_),
    .X(net3828));
 sg13g2_dlygate4sd3_1 hold1569 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][3] ),
    .X(net3829));
 sg13g2_dlygate4sd3_1 hold1570 (.A(\i_peripherals.i_user_peri39.math_result_reg[1] ),
    .X(net3830));
 sg13g2_dlygate4sd3_1 hold1571 (.A(\i_tinyqv.cpu.imm[19] ),
    .X(net3831));
 sg13g2_dlygate4sd3_1 hold1572 (.A(\i_tinyqv.cpu.i_core.i_shift.a[17] ),
    .X(net3832));
 sg13g2_dlygate4sd3_1 hold1573 (.A(_00526_),
    .X(net3833));
 sg13g2_dlygate4sd3_1 hold1574 (.A(\i_peripherals.i_user_peri39.math_result_reg[3] ),
    .X(net3834));
 sg13g2_dlygate4sd3_1 hold1575 (.A(\i_peripherals.i_uart.i_uart_rx.fsm_state[2] ),
    .X(net3835));
 sg13g2_dlygate4sd3_1 hold1576 (.A(_05482_),
    .X(net3836));
 sg13g2_dlygate4sd3_1 hold1577 (.A(_00348_),
    .X(net3837));
 sg13g2_dlygate4sd3_1 hold1578 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][0] ),
    .X(net3838));
 sg13g2_dlygate4sd3_1 hold1579 (.A(\i_tinyqv.cpu.additional_mem_ops[1] ),
    .X(net3839));
 sg13g2_dlygate4sd3_1 hold1580 (.A(_00909_),
    .X(net3840));
 sg13g2_dlygate4sd3_1 hold1581 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[2] ),
    .X(net3841));
 sg13g2_dlygate4sd3_1 hold1582 (.A(_00176_),
    .X(net3842));
 sg13g2_dlygate4sd3_1 hold1583 (.A(\i_tinyqv.cpu.is_system ),
    .X(net3843));
 sg13g2_dlygate4sd3_1 hold1584 (.A(\i_tinyqv.cpu.instr_data_in[2] ),
    .X(net3844));
 sg13g2_dlygate4sd3_1 hold1585 (.A(_00670_),
    .X(net3845));
 sg13g2_dlygate4sd3_1 hold1586 (.A(\i_peripherals.i_user_peri39.math_result_reg[10] ),
    .X(net3846));
 sg13g2_dlygate4sd3_1 hold1587 (.A(\i_tinyqv.cpu.imm[20] ),
    .X(net3847));
 sg13g2_dlygate4sd3_1 hold1588 (.A(\i_tinyqv.cpu.i_core.i_shift.a[18] ),
    .X(net3848));
 sg13g2_dlygate4sd3_1 hold1589 (.A(_00527_),
    .X(net3849));
 sg13g2_dlygate4sd3_1 hold1590 (.A(\i_peripherals.i_user_peri39.math_result_reg[14] ),
    .X(net3850));
 sg13g2_dlygate4sd3_1 hold1591 (.A(_00156_),
    .X(net3851));
 sg13g2_dlygate4sd3_1 hold1592 (.A(\addr[0] ),
    .X(net3852));
 sg13g2_dlygate4sd3_1 hold1593 (.A(_00848_),
    .X(net3853));
 sg13g2_dlygate4sd3_1 hold1594 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[1][2] ),
    .X(net3854));
 sg13g2_dlygate4sd3_1 hold1595 (.A(\i_peripherals.i_user_peri39.math_result_reg[16] ),
    .X(net3855));
 sg13g2_dlygate4sd3_1 hold1596 (.A(_00158_),
    .X(net3856));
 sg13g2_dlygate4sd3_1 hold1597 (.A(\i_tinyqv.mem.q_ctrl.spi_flash_select ),
    .X(net3857));
 sg13g2_dlygate4sd3_1 hold1598 (.A(\i_peripherals.i_user_peri39.math_result_reg[17] ),
    .X(net3858));
 sg13g2_dlygate4sd3_1 hold1599 (.A(_00159_),
    .X(net3859));
 sg13g2_dlygate4sd3_1 hold1600 (.A(\i_peripherals.i_uart.baud_divider[5] ),
    .X(net3860));
 sg13g2_dlygate4sd3_1 hold1601 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[8] ),
    .X(net3861));
 sg13g2_dlygate4sd3_1 hold1602 (.A(\i_tinyqv.cpu.i_core.i_shift.b[2] ),
    .X(net3862));
 sg13g2_dlygate4sd3_1 hold1603 (.A(debug_register_data),
    .X(net3863));
 sg13g2_dlygate4sd3_1 hold1604 (.A(_00456_),
    .X(net3864));
 sg13g2_dlygate4sd3_1 hold1605 (.A(\i_tinyqv.cpu.i_core.mie[2] ),
    .X(net3865));
 sg13g2_dlygate4sd3_1 hold1606 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[0] ),
    .X(net3866));
 sg13g2_dlygate4sd3_1 hold1607 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[5] ),
    .X(net3867));
 sg13g2_dlygate4sd3_1 hold1608 (.A(\i_peripherals.i_user_peri39.math_result_reg[28] ),
    .X(net3868));
 sg13g2_dlygate4sd3_1 hold1609 (.A(\i_peripherals.i_user_peri39.math_result_reg[29] ),
    .X(net3869));
 sg13g2_dlygate4sd3_1 hold1610 (.A(\i_peripherals.data_out[12] ),
    .X(net3870));
 sg13g2_dlygate4sd3_1 hold1611 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[4] ),
    .X(net3871));
 sg13g2_dlygate4sd3_1 hold1612 (.A(_00178_),
    .X(net3872));
 sg13g2_dlygate4sd3_1 hold1613 (.A(\i_tinyqv.cpu.instr_data_start[9] ),
    .X(net3873));
 sg13g2_dlygate4sd3_1 hold1614 (.A(\i_tinyqv.cpu.i_core.cycle[1] ),
    .X(net3874));
 sg13g2_dlygate4sd3_1 hold1615 (.A(\i_peripherals.i_user_peri39.math_result_reg[13] ),
    .X(net3875));
 sg13g2_dlygate4sd3_1 hold1616 (.A(_00155_),
    .X(net3876));
 sg13g2_dlygate4sd3_1 hold1617 (.A(\i_peripherals.i_uart.baud_divider[2] ),
    .X(net3877));
 sg13g2_dlygate4sd3_1 hold1618 (.A(_00302_),
    .X(net3878));
 sg13g2_dlygate4sd3_1 hold1619 (.A(\gpio_out_sel[6] ),
    .X(net3879));
 sg13g2_dlygate4sd3_1 hold1620 (.A(_00000_),
    .X(net3880));
 sg13g2_dlygate4sd3_1 hold1621 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[7][3] ),
    .X(net3881));
 sg13g2_dlygate4sd3_1 hold1622 (.A(\i_tinyqv.mem.data_txn_len[1] ),
    .X(net3882));
 sg13g2_dlygate4sd3_1 hold1623 (.A(_06508_),
    .X(net3883));
 sg13g2_dlygate4sd3_1 hold1624 (.A(_00664_),
    .X(net3884));
 sg13g2_dlygate4sd3_1 hold1625 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][3] ),
    .X(net3885));
 sg13g2_dlygate4sd3_1 hold1626 (.A(\i_peripherals.i_user_peri39.math_result_reg[18] ),
    .X(net3886));
 sg13g2_dlygate4sd3_1 hold1627 (.A(\i_tinyqv.cpu.i_core.imm_lo[2] ),
    .X(net3887));
 sg13g2_dlygate4sd3_1 hold1628 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[0] ),
    .X(net3888));
 sg13g2_dlygate4sd3_1 hold1629 (.A(_02665_),
    .X(net3889));
 sg13g2_dlygate4sd3_1 hold1630 (.A(_00099_),
    .X(net3890));
 sg13g2_dlygate4sd3_1 hold1631 (.A(\i_tinyqv.cpu.i_core.imm_lo[7] ),
    .X(net3891));
 sg13g2_dlygate4sd3_1 hold1632 (.A(\i_peripherals.i_uart.baud_divider[11] ),
    .X(net3892));
 sg13g2_dlygate4sd3_1 hold1633 (.A(_00586_),
    .X(net3893));
 sg13g2_dlygate4sd3_1 hold1634 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][0] ),
    .X(net3894));
 sg13g2_dlygate4sd3_1 hold1635 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[16] ),
    .X(net3895));
 sg13g2_dlygate4sd3_1 hold1636 (.A(\i_tinyqv.cpu.instr_data_start[8] ),
    .X(net3896));
 sg13g2_dlygate4sd3_1 hold1637 (.A(\i_peripherals.i_uart.baud_divider[0] ),
    .X(net3897));
 sg13g2_dlygate4sd3_1 hold1638 (.A(_00300_),
    .X(net3898));
 sg13g2_dlygate4sd3_1 hold1639 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[2] ),
    .X(net3899));
 sg13g2_dlygate4sd3_1 hold1640 (.A(_02667_),
    .X(net3900));
 sg13g2_dlygate4sd3_1 hold1641 (.A(_00101_),
    .X(net3901));
 sg13g2_dlygate4sd3_1 hold1642 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][0] ),
    .X(net3902));
 sg13g2_dlygate4sd3_1 hold1643 (.A(\i_tinyqv.cpu.i_core.mstatus_mie ),
    .X(net3903));
 sg13g2_dlygate4sd3_1 hold1644 (.A(\i_tinyqv.cpu.imm[13] ),
    .X(net3904));
 sg13g2_dlygate4sd3_1 hold1645 (.A(\i_peripherals.i_user_peri39.math_result_reg[25] ),
    .X(net3905));
 sg13g2_dlygate4sd3_1 hold1646 (.A(_00167_),
    .X(net3906));
 sg13g2_dlygate4sd3_1 hold1647 (.A(\i_tinyqv.cpu.imm[12] ),
    .X(net3907));
 sg13g2_dlygate4sd3_1 hold1648 (.A(\i_tinyqv.cpu.i_core.mie[1] ),
    .X(net3908));
 sg13g2_dlygate4sd3_1 hold1649 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[9][1] ),
    .X(net3909));
 sg13g2_dlygate4sd3_1 hold1650 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[5] ),
    .X(net3910));
 sg13g2_dlygate4sd3_1 hold1651 (.A(\i_tinyqv.cpu.imm[17] ),
    .X(net3911));
 sg13g2_dlygate4sd3_1 hold1652 (.A(\i_tinyqv.cpu.i_timer.time_pulse_r ),
    .X(net3912));
 sg13g2_dlygate4sd3_1 hold1653 (.A(_02835_),
    .X(net3913));
 sg13g2_dlygate4sd3_1 hold1654 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[2] ),
    .X(net3914));
 sg13g2_dlygate4sd3_1 hold1655 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][2] ),
    .X(net3915));
 sg13g2_dlygate4sd3_1 hold1656 (.A(\i_tinyqv.cpu.addr_offset[2] ),
    .X(net3916));
 sg13g2_dlygate4sd3_1 hold1657 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[1] ),
    .X(net3917));
 sg13g2_dlygate4sd3_1 hold1658 (.A(\i_tinyqv.cpu.i_core.i_shift.a[10] ),
    .X(net3918));
 sg13g2_dlygate4sd3_1 hold1659 (.A(\i_tinyqv.cpu.imm[18] ),
    .X(net3919));
 sg13g2_dlygate4sd3_1 hold1660 (.A(\i_tinyqv.cpu.i_core.mie[16] ),
    .X(net3920));
 sg13g2_dlygate4sd3_1 hold1661 (.A(\i_peripherals.i_uart.baud_divider[7] ),
    .X(net3921));
 sg13g2_dlygate4sd3_1 hold1662 (.A(_00307_),
    .X(net3922));
 sg13g2_dlygate4sd3_1 hold1663 (.A(\i_tinyqv.cpu.i_core.i_instrret.data[1] ),
    .X(net3923));
 sg13g2_dlygate4sd3_1 hold1664 (.A(\i_peripherals.i_uart.baud_divider[9] ),
    .X(net3924));
 sg13g2_dlygate4sd3_1 hold1665 (.A(_00584_),
    .X(net3925));
 sg13g2_dlygate4sd3_1 hold1666 (.A(\i_tinyqv.cpu.alu_op[0] ),
    .X(net3926));
 sg13g2_dlygate4sd3_1 hold1667 (.A(\i_peripherals.i_user_peri39.math_result_reg[4] ),
    .X(net3927));
 sg13g2_dlygate4sd3_1 hold1668 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][3] ),
    .X(net3928));
 sg13g2_dlygate4sd3_1 hold1669 (.A(\i_tinyqv.cpu.i_core.i_shift.a[21] ),
    .X(net3929));
 sg13g2_dlygate4sd3_1 hold1670 (.A(_00530_),
    .X(net3930));
 sg13g2_dlygate4sd3_1 hold1671 (.A(\i_tinyqv.cpu.i_core.i_shift.a[25] ),
    .X(net3931));
 sg13g2_dlygate4sd3_1 hold1672 (.A(\i_tinyqv.cpu.instr_data_in[7] ),
    .X(net3932));
 sg13g2_dlygate4sd3_1 hold1673 (.A(_00675_),
    .X(net3933));
 sg13g2_dlygate4sd3_1 hold1674 (.A(\i_peripherals.i_uart.baud_divider[3] ),
    .X(net3934));
 sg13g2_dlygate4sd3_1 hold1675 (.A(_00303_),
    .X(net3935));
 sg13g2_dlygate4sd3_1 hold1676 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][2] ),
    .X(net3936));
 sg13g2_dlygate4sd3_1 hold1677 (.A(\i_peripherals.i_user_peri39.busy_counter[2] ),
    .X(net3937));
 sg13g2_dlygate4sd3_1 hold1678 (.A(\i_peripherals.i_uart.baud_divider[1] ),
    .X(net3938));
 sg13g2_dlygate4sd3_1 hold1679 (.A(_00301_),
    .X(net3939));
 sg13g2_dlygate4sd3_1 hold1680 (.A(\addr[25] ),
    .X(net3940));
 sg13g2_dlygate4sd3_1 hold1681 (.A(\i_tinyqv.cpu.i_core.i_shift.a[23] ),
    .X(net3941));
 sg13g2_dlygate4sd3_1 hold1682 (.A(_00532_),
    .X(net3942));
 sg13g2_dlygate4sd3_1 hold1683 (.A(\i_tinyqv.cpu.i_core.cycle_count[3] ),
    .X(net3943));
 sg13g2_dlygate4sd3_1 hold1684 (.A(_02658_),
    .X(net3944));
 sg13g2_dlygate4sd3_1 hold1685 (.A(\i_tinyqv.mem.data_txn_len[0] ),
    .X(net3945));
 sg13g2_dlygate4sd3_1 hold1686 (.A(_06505_),
    .X(net3946));
 sg13g2_dlygate4sd3_1 hold1687 (.A(_00663_),
    .X(net3947));
 sg13g2_dlygate4sd3_1 hold1688 (.A(\i_tinyqv.cpu.i_timer.i_mtime.data[0] ),
    .X(net3948));
 sg13g2_dlygate4sd3_1 hold1689 (.A(_06490_),
    .X(net3949));
 sg13g2_dlygate4sd3_1 hold1690 (.A(\i_tinyqv.cpu.i_core.i_shift.a[22] ),
    .X(net3950));
 sg13g2_dlygate4sd3_1 hold1691 (.A(_00531_),
    .X(net3951));
 sg13g2_dlygate4sd3_1 hold1692 (.A(\i_peripherals.i_user_peri39.math_result_reg[26] ),
    .X(net3952));
 sg13g2_dlygate4sd3_1 hold1693 (.A(_00168_),
    .X(net3953));
 sg13g2_dlygate4sd3_1 hold1694 (.A(\i_tinyqv.cpu.instr_data_in[11] ),
    .X(net3954));
 sg13g2_dlygate4sd3_1 hold1695 (.A(_00729_),
    .X(net3955));
 sg13g2_dlygate4sd3_1 hold1696 (.A(\i_debug_uart_tx.fsm_state[2] ),
    .X(net3956));
 sg13g2_dlygate4sd3_1 hold1697 (.A(_05810_),
    .X(net3957));
 sg13g2_dlygate4sd3_1 hold1698 (.A(_00434_),
    .X(net3958));
 sg13g2_dlygate4sd3_1 hold1699 (.A(\i_peripherals.i_user_peri39.math_result_reg[7] ),
    .X(net3959));
 sg13g2_dlygate4sd3_1 hold1700 (.A(\addr[9] ),
    .X(net3960));
 sg13g2_dlygate4sd3_1 hold1701 (.A(\i_tinyqv.cpu.imm[16] ),
    .X(net3961));
 sg13g2_dlygate4sd3_1 hold1702 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][0] ),
    .X(net3962));
 sg13g2_dlygate4sd3_1 hold1703 (.A(\i_tinyqv.cpu.instr_data_start[22] ),
    .X(net3963));
 sg13g2_dlygate4sd3_1 hold1704 (.A(\i_tinyqv.cpu.i_core.mem_op[2] ),
    .X(net3964));
 sg13g2_dlygate4sd3_1 hold1705 (.A(\i_tinyqv.cpu.imm[21] ),
    .X(net3965));
 sg13g2_dlygate4sd3_1 hold1706 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[4] ),
    .X(net3966));
 sg13g2_dlygate4sd3_1 hold1707 (.A(\i_tinyqv.mem.q_ctrl.stop_txn_reg ),
    .X(net3967));
 sg13g2_dlygate4sd3_1 hold1708 (.A(_00712_),
    .X(net3968));
 sg13g2_dlygate4sd3_1 hold1709 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][2] ),
    .X(net3969));
 sg13g2_dlygate4sd3_1 hold1710 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[1] ),
    .X(net3970));
 sg13g2_dlygate4sd3_1 hold1711 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][1] ),
    .X(net3971));
 sg13g2_dlygate4sd3_1 hold1712 (.A(\i_tinyqv.cpu.instr_data_start[21] ),
    .X(net3972));
 sg13g2_dlygate4sd3_1 hold1713 (.A(\i_tinyqv.cpu.i_core.mip[16] ),
    .X(net3973));
 sg13g2_dlygate4sd3_1 hold1714 (.A(_00136_),
    .X(net3974));
 sg13g2_dlygate4sd3_1 hold1715 (.A(\addr[3] ),
    .X(net3975));
 sg13g2_dlygate4sd3_1 hold1716 (.A(\i_peripherals.i_uart.i_uart_rx.fsm_state[1] ),
    .X(net3976));
 sg13g2_dlygate4sd3_1 hold1717 (.A(_05327_),
    .X(net3977));
 sg13g2_dlygate4sd3_1 hold1718 (.A(_05485_),
    .X(net3978));
 sg13g2_dlygate4sd3_1 hold1719 (.A(\i_tinyqv.cpu.i_core.imm_lo[10] ),
    .X(net3979));
 sg13g2_dlygate4sd3_1 hold1720 (.A(\i_tinyqv.cpu.i_core.i_shift.a[27] ),
    .X(net3980));
 sg13g2_dlygate4sd3_1 hold1721 (.A(_00536_),
    .X(net3981));
 sg13g2_dlygate4sd3_1 hold1722 (.A(\i_peripherals.i_uart.i_uart_tx.fsm_state[3] ),
    .X(net3982));
 sg13g2_dlygate4sd3_1 hold1723 (.A(\time_count[2] ),
    .X(net3983));
 sg13g2_dlygate4sd3_1 hold1724 (.A(_07230_),
    .X(net3984));
 sg13g2_dlygate4sd3_1 hold1725 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[12] ),
    .X(net3985));
 sg13g2_dlygate4sd3_1 hold1726 (.A(\i_peripherals.i_uart.baud_divider[4] ),
    .X(net3986));
 sg13g2_dlygate4sd3_1 hold1727 (.A(_00304_),
    .X(net3987));
 sg13g2_dlygate4sd3_1 hold1728 (.A(\i_debug_uart_tx.fsm_state[0] ),
    .X(net3988));
 sg13g2_dlygate4sd3_1 hold1729 (.A(_00432_),
    .X(net3989));
 sg13g2_dlygate4sd3_1 hold1730 (.A(\i_tinyqv.cpu.instr_data_in[9] ),
    .X(net3990));
 sg13g2_dlygate4sd3_1 hold1731 (.A(_06718_),
    .X(net3991));
 sg13g2_dlygate4sd3_1 hold1732 (.A(_00727_),
    .X(net3992));
 sg13g2_dlygate4sd3_1 hold1733 (.A(\i_tinyqv.cpu.i_core.i_shift.a[2] ),
    .X(net3993));
 sg13g2_dlygate4sd3_1 hold1734 (.A(_00511_),
    .X(net3994));
 sg13g2_dlygate4sd3_1 hold1735 (.A(\i_tinyqv.cpu.imm[15] ),
    .X(net3995));
 sg13g2_dlygate4sd3_1 hold1736 (.A(\i_tinyqv.cpu.instr_data_in[14] ),
    .X(net3996));
 sg13g2_dlygate4sd3_1 hold1737 (.A(_00732_),
    .X(net3997));
 sg13g2_dlygate4sd3_1 hold1738 (.A(\i_tinyqv.cpu.imm[14] ),
    .X(net3998));
 sg13g2_dlygate4sd3_1 hold1739 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][3] ),
    .X(net3999));
 sg13g2_dlygate4sd3_1 hold1740 (.A(\i_peripherals.i_user_peri39.math_result_reg[9] ),
    .X(net4000));
 sg13g2_dlygate4sd3_1 hold1741 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[10][3] ),
    .X(net4001));
 sg13g2_dlygate4sd3_1 hold1742 (.A(debug_data_continue),
    .X(net4002));
 sg13g2_dlygate4sd3_1 hold1743 (.A(_02637_),
    .X(net4003));
 sg13g2_dlygate4sd3_1 hold1744 (.A(_00019_),
    .X(net4004));
 sg13g2_dlygate4sd3_1 hold1745 (.A(\addr[11] ),
    .X(net4005));
 sg13g2_dlygate4sd3_1 hold1746 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[5][0] ),
    .X(net4006));
 sg13g2_dlygate4sd3_1 hold1747 (.A(\i_tinyqv.cpu.i_core.imm_lo[3] ),
    .X(net4007));
 sg13g2_dlygate4sd3_1 hold1748 (.A(\i_tinyqv.cpu.is_jalr ),
    .X(net4008));
 sg13g2_dlygate4sd3_1 hold1749 (.A(\i_tinyqv.cpu.i_core.imm_lo[4] ),
    .X(net4009));
 sg13g2_dlygate4sd3_1 hold1750 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][3] ),
    .X(net4010));
 sg13g2_dlygate4sd3_1 hold1751 (.A(\i_tinyqv.cpu.instr_data_start[5] ),
    .X(net4011));
 sg13g2_dlygate4sd3_1 hold1752 (.A(\i_tinyqv.cpu.additional_mem_ops[0] ),
    .X(net4012));
 sg13g2_dlygate4sd3_1 hold1753 (.A(\addr[26] ),
    .X(net4013));
 sg13g2_dlygate4sd3_1 hold1754 (.A(_07076_),
    .X(net4014));
 sg13g2_dlygate4sd3_1 hold1755 (.A(\i_peripherals.i_uart.baud_divider[6] ),
    .X(net4015));
 sg13g2_dlygate4sd3_1 hold1756 (.A(_00306_),
    .X(net4016));
 sg13g2_dlygate4sd3_1 hold1757 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[15][2] ),
    .X(net4017));
 sg13g2_dlygate4sd3_1 hold1758 (.A(\i_tinyqv.cpu.i_core.i_shift.a[26] ),
    .X(net4018));
 sg13g2_dlygate4sd3_1 hold1759 (.A(_00535_),
    .X(net4019));
 sg13g2_dlygate4sd3_1 hold1760 (.A(\time_count[3] ),
    .X(net4020));
 sg13g2_dlygate4sd3_1 hold1761 (.A(_07232_),
    .X(net4021));
 sg13g2_dlygate4sd3_1 hold1762 (.A(_00919_),
    .X(net4022));
 sg13g2_dlygate4sd3_1 hold1763 (.A(\i_peripherals.i_uart.i_uart_rx.fsm_state[0] ),
    .X(net4023));
 sg13g2_dlygate4sd3_1 hold1764 (.A(\i_tinyqv.cpu.alu_op[3] ),
    .X(net4024));
 sg13g2_dlygate4sd3_1 hold1765 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][2] ),
    .X(net4025));
 sg13g2_dlygate4sd3_1 hold1766 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[11][1] ),
    .X(net4026));
 sg13g2_dlygate4sd3_1 hold1767 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][2] ),
    .X(net4027));
 sg13g2_dlygate4sd3_1 hold1768 (.A(\i_tinyqv.mem.qspi_data_byte_idx[0] ),
    .X(net4028));
 sg13g2_dlygate4sd3_1 hold1769 (.A(_00666_),
    .X(net4029));
 sg13g2_dlygate4sd3_1 hold1770 (.A(\i_tinyqv.mem.qspi_data_byte_idx[1] ),
    .X(net4030));
 sg13g2_dlygate4sd3_1 hold1771 (.A(_06517_),
    .X(net4031));
 sg13g2_dlygate4sd3_1 hold1772 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[14] ),
    .X(net4032));
 sg13g2_dlygate4sd3_1 hold1773 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[7] ),
    .X(net4033));
 sg13g2_dlygate4sd3_1 hold1774 (.A(\data_to_write[9] ),
    .X(net4034));
 sg13g2_dlygate4sd3_1 hold1775 (.A(\data_to_write[20] ),
    .X(net4035));
 sg13g2_dlygate4sd3_1 hold1776 (.A(\i_tinyqv.cpu.instr_data_start[23] ),
    .X(net4036));
 sg13g2_dlygate4sd3_1 hold1777 (.A(\i_peripherals.i_uart.i_uart_rx.cycle_counter[12] ),
    .X(net4037));
 sg13g2_dlygate4sd3_1 hold1778 (.A(\i_tinyqv.cpu.i_timer.i_mtime.data[3] ),
    .X(net4038));
 sg13g2_dlygate4sd3_1 hold1779 (.A(_00135_),
    .X(net4039));
 sg13g2_dlygate4sd3_1 hold1780 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[8][3] ),
    .X(net4040));
 sg13g2_dlygate4sd3_1 hold1781 (.A(\i_tinyqv.cpu.i_core.i_shift.a[31] ),
    .X(net4041));
 sg13g2_dlygate4sd3_1 hold1782 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[3] ),
    .X(net4042));
 sg13g2_dlygate4sd3_1 hold1783 (.A(\i_tinyqv.cpu.i_core.imm_lo[5] ),
    .X(net4043));
 sg13g2_dlygate4sd3_1 hold1784 (.A(\addr[8] ),
    .X(net4044));
 sg13g2_dlygate4sd3_1 hold1785 (.A(\i_tinyqv.cpu.i_core.cycle_count[1] ),
    .X(net4045));
 sg13g2_dlygate4sd3_1 hold1786 (.A(_02654_),
    .X(net4046));
 sg13g2_dlygate4sd3_1 hold1787 (.A(_00093_),
    .X(net4047));
 sg13g2_dlygate4sd3_1 hold1788 (.A(\i_tinyqv.cpu.i_core.imm_lo[6] ),
    .X(net4048));
 sg13g2_dlygate4sd3_1 hold1789 (.A(\i_tinyqv.cpu.i_core.mem_op[1] ),
    .X(net4049));
 sg13g2_dlygate4sd3_1 hold1790 (.A(_00843_),
    .X(net4050));
 sg13g2_dlygate4sd3_1 hold1791 (.A(\i_tinyqv.cpu.data_write_n[0] ),
    .X(net4051));
 sg13g2_dlygate4sd3_1 hold1792 (.A(_00842_),
    .X(net4052));
 sg13g2_dlygate4sd3_1 hold1793 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[21] ),
    .X(net4053));
 sg13g2_dlygate4sd3_1 hold1794 (.A(\i_tinyqv.cpu.instr_data_start[11] ),
    .X(net4054));
 sg13g2_dlygate4sd3_1 hold1795 (.A(\i_tinyqv.cpu.instr_data_in[6] ),
    .X(net4055));
 sg13g2_dlygate4sd3_1 hold1796 (.A(_00674_),
    .X(net4056));
 sg13g2_dlygate4sd3_1 hold1797 (.A(\i_tinyqv.cpu.instr_fetch_started ),
    .X(net4057));
 sg13g2_dlygate4sd3_1 hold1798 (.A(_06969_),
    .X(net4058));
 sg13g2_dlygate4sd3_1 hold1799 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[2][1] ),
    .X(net4059));
 sg13g2_dlygate4sd3_1 hold1800 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[17] ),
    .X(net4060));
 sg13g2_dlygate4sd3_1 hold1801 (.A(\addr[5] ),
    .X(net4061));
 sg13g2_dlygate4sd3_1 hold1802 (.A(_00853_),
    .X(net4062));
 sg13g2_dlygate4sd3_1 hold1803 (.A(\i_tinyqv.cpu.instr_data_start[6] ),
    .X(net4063));
 sg13g2_dlygate4sd3_1 hold1804 (.A(\i_tinyqv.cpu.instr_data_start[16] ),
    .X(net4064));
 sg13g2_dlygate4sd3_1 hold1805 (.A(\i_tinyqv.cpu.i_core.i_registers.reg_access[13][1] ),
    .X(net4065));
 sg13g2_dlygate4sd3_1 hold1806 (.A(\addr[2] ),
    .X(net4066));
 sg13g2_dlygate4sd3_1 hold1807 (.A(\i_tinyqv.cpu.i_core.i_cycles.cy ),
    .X(net4067));
 sg13g2_dlygate4sd3_1 hold1808 (.A(_02650_),
    .X(net4068));
 sg13g2_dlygate4sd3_1 hold1809 (.A(_00092_),
    .X(net4069));
 sg13g2_dlygate4sd3_1 hold1810 (.A(\i_tinyqv.cpu.instr_data_start[18] ),
    .X(net4070));
 sg13g2_dlygate4sd3_1 hold1811 (.A(\i_tinyqv.mem.q_ctrl.is_writing ),
    .X(net4071));
 sg13g2_dlygate4sd3_1 hold1812 (.A(_00704_),
    .X(net4072));
 sg13g2_dlygate4sd3_1 hold1813 (.A(\i_tinyqv.cpu.instr_data_in[8] ),
    .X(net4073));
 sg13g2_dlygate4sd3_1 hold1814 (.A(\i_tinyqv.cpu.instr_data_start[12] ),
    .X(net4074));
 sg13g2_dlygate4sd3_1 hold1815 (.A(\i_tinyqv.cpu.i_core.i_registers.rs1[3] ),
    .X(net4075));
 sg13g2_dlygate4sd3_1 hold1816 (.A(\i_tinyqv.cpu.instr_data_in[12] ),
    .X(net4076));
 sg13g2_dlygate4sd3_1 hold1817 (.A(\i_tinyqv.cpu.pc[2] ),
    .X(net4077));
 sg13g2_dlygate4sd3_1 hold1818 (.A(\i_tinyqv.cpu.pc[1] ),
    .X(net4078));
 sg13g2_dlygate4sd3_1 hold1819 (.A(\i_tinyqv.cpu.i_core.time_hi[1] ),
    .X(net4079));
 sg13g2_dlygate4sd3_1 hold1820 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[13] ),
    .X(net4080));
 sg13g2_dlygate4sd3_1 hold1821 (.A(\time_count[1] ),
    .X(net4081));
 sg13g2_dlygate4sd3_1 hold1822 (.A(\data_to_write[6] ),
    .X(net4082));
 sg13g2_dlygate4sd3_1 hold1823 (.A(_00425_),
    .X(net4083));
 sg13g2_dlygate4sd3_1 hold1824 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[11] ),
    .X(net4084));
 sg13g2_dlygate4sd3_1 hold1825 (.A(\addr[27] ),
    .X(net4085));
 sg13g2_dlygate4sd3_1 hold1826 (.A(\i_tinyqv.cpu.instr_data_in[5] ),
    .X(net4086));
 sg13g2_dlygate4sd3_1 hold1827 (.A(_00673_),
    .X(net4087));
 sg13g2_dlygate4sd3_1 hold1828 (.A(\i_peripherals.i_uart.uart_rx_buffered ),
    .X(net4088));
 sg13g2_dlygate4sd3_1 hold1829 (.A(\i_tinyqv.cpu.i_core.imm_lo[11] ),
    .X(net4089));
 sg13g2_dlygate4sd3_1 hold1830 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[2] ),
    .X(net4090));
 sg13g2_dlygate4sd3_1 hold1831 (.A(\time_limit[5] ),
    .X(net4091));
 sg13g2_dlygate4sd3_1 hold1832 (.A(_00005_),
    .X(net4092));
 sg13g2_dlygate4sd3_1 hold1833 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[2] ),
    .X(net4093));
 sg13g2_dlygate4sd3_1 hold1834 (.A(_00715_),
    .X(net4094));
 sg13g2_dlygate4sd3_1 hold1835 (.A(\data_to_write[8] ),
    .X(net4095));
 sg13g2_dlygate4sd3_1 hold1836 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[1] ),
    .X(net4096));
 sg13g2_dlygate4sd3_1 hold1837 (.A(\i_tinyqv.cpu.i_core.imm_lo[8] ),
    .X(net4097));
 sg13g2_dlygate4sd3_1 hold1838 (.A(\data_to_write[5] ),
    .X(net4098));
 sg13g2_dlygate4sd3_1 hold1839 (.A(\i_tinyqv.cpu.instr_data_in[13] ),
    .X(net4099));
 sg13g2_dlygate4sd3_1 hold1840 (.A(\i_peripherals.data_ready_r ),
    .X(net4100));
 sg13g2_dlygate4sd3_1 hold1841 (.A(\i_tinyqv.cpu.instr_data_start[7] ),
    .X(net4101));
 sg13g2_dlygate4sd3_1 hold1842 (.A(\data_to_write[3] ),
    .X(net4102));
 sg13g2_dlygate4sd3_1 hold1843 (.A(_00003_),
    .X(net4103));
 sg13g2_dlygate4sd3_1 hold1844 (.A(\i_tinyqv.cpu.i_core.i_shift.a[5] ),
    .X(net4104));
 sg13g2_dlygate4sd3_1 hold1845 (.A(_00510_),
    .X(net4105));
 sg13g2_dlygate4sd3_1 hold1846 (.A(\i_tinyqv.cpu.i_timer.mtimecmp[6] ),
    .X(net4106));
 sg13g2_dlygate4sd3_1 hold1847 (.A(\data_to_write[10] ),
    .X(net4107));
 sg13g2_dlygate4sd3_1 hold1848 (.A(\data_to_write[11] ),
    .X(net4108));
 sg13g2_dlygate4sd3_1 hold1849 (.A(\i_tinyqv.cpu.i_core.i_registers.rs2[0] ),
    .X(net4109));
 sg13g2_dlygate4sd3_1 hold1850 (.A(\i_tinyqv.cpu.instr_data_start[17] ),
    .X(net4110));
 sg13g2_dlygate4sd3_1 hold1851 (.A(\i_tinyqv.cpu.instr_data_start[4] ),
    .X(net4111));
 sg13g2_dlygate4sd3_1 hold1852 (.A(\i_tinyqv.cpu.instr_data_in[15] ),
    .X(net4112));
 sg13g2_dlygate4sd3_1 hold1853 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[2] ),
    .X(net4113));
 sg13g2_dlygate4sd3_1 hold1854 (.A(\i_tinyqv.mem.instr_active ),
    .X(net4114));
 sg13g2_dlygate4sd3_1 hold1855 (.A(_06590_),
    .X(net4115));
 sg13g2_dlygate4sd3_1 hold1856 (.A(_00701_),
    .X(net4116));
 sg13g2_dlygate4sd3_1 hold1857 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .X(net4117));
 sg13g2_dlygate4sd3_1 hold1858 (.A(\i_tinyqv.cpu.i_core.imm_lo[9] ),
    .X(net4118));
 sg13g2_dlygate4sd3_1 hold1859 (.A(\time_limit[2] ),
    .X(net4119));
 sg13g2_dlygate4sd3_1 hold1860 (.A(_00002_),
    .X(net4120));
 sg13g2_dlygate4sd3_1 hold1861 (.A(\i_tinyqv.cpu.alu_op[1] ),
    .X(net4121));
 sg13g2_dlygate4sd3_1 hold1862 (.A(\time_limit[4] ),
    .X(net4122));
 sg13g2_dlygate4sd3_1 hold1863 (.A(_00004_),
    .X(net4123));
 sg13g2_dlygate4sd3_1 hold1864 (.A(\data_to_write[12] ),
    .X(net4124));
 sg13g2_dlygate4sd3_1 hold1865 (.A(\i_tinyqv.mem.q_ctrl.fsm_state[0] ),
    .X(net4125));
 sg13g2_dlygate4sd3_1 hold1866 (.A(\i_tinyqv.cpu.i_core.i_shift.a[9] ),
    .X(net4126));
 sg13g2_dlygate4sd3_1 hold1867 (.A(\i_tinyqv.cpu.i_core.cycle[0] ),
    .X(net4127));
 sg13g2_dlygate4sd3_1 hold1868 (.A(\data_to_write[1] ),
    .X(net4128));
 sg13g2_dlygate4sd3_1 hold1869 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .X(net4129));
 sg13g2_dlygate4sd3_1 hold1870 (.A(\gpio_out_sel[7] ),
    .X(net4130));
 sg13g2_dlygate4sd3_1 hold1871 (.A(_00001_),
    .X(net4131));
 sg13g2_dlygate4sd3_1 hold1872 (.A(\i_tinyqv.cpu.i_core.imm_lo[1] ),
    .X(net4132));
 sg13g2_dlygate4sd3_1 hold1873 (.A(\i_tinyqv.cpu.i_core.i_shift.a[8] ),
    .X(net4133));
 sg13g2_dlygate4sd3_1 hold1874 (.A(\i_tinyqv.cpu.instr_data_in[10] ),
    .X(net4134));
 sg13g2_dlygate4sd3_1 hold1875 (.A(\addr[4] ),
    .X(net4135));
 sg13g2_dlygate4sd3_1 hold1876 (.A(\i_tinyqv.cpu.instr_data_start[14] ),
    .X(net4136));
 sg13g2_dlygate4sd3_1 hold1877 (.A(\i_tinyqv.mem.qspi_write_done ),
    .X(net4137));
 sg13g2_dlygate4sd3_1 hold1878 (.A(\i_tinyqv.cpu.instr_data_start[19] ),
    .X(net4138));
 sg13g2_dlygate4sd3_1 hold1879 (.A(\i_tinyqv.cpu.instr_fetch_running ),
    .X(net4139));
 sg13g2_dlygate4sd3_1 hold1880 (.A(\data_to_write[4] ),
    .X(net4140));
 sg13g2_dlygate4sd3_1 hold1881 (.A(\i_debug_uart_tx.data_to_send[6] ),
    .X(net4141));
 sg13g2_dlygate4sd3_1 hold1882 (.A(\i_tinyqv.cpu.i_timer.i_mtime.data[2] ),
    .X(net4142));
 sg13g2_dlygate4sd3_1 hold1883 (.A(\i_tinyqv.cpu.instr_data_start[10] ),
    .X(net4143));
 sg13g2_dlygate4sd3_1 hold1884 (.A(\i_tinyqv.cpu.is_load ),
    .X(net4144));
 sg13g2_dlygate4sd3_1 hold1885 (.A(\i_tinyqv.cpu.instr_data_start[20] ),
    .X(net4145));
 sg13g2_dlygate4sd3_1 hold1886 (.A(_06947_),
    .X(net4146));
 sg13g2_dlygate4sd3_1 hold1887 (.A(\i_tinyqv.cpu.instr_data_start[13] ),
    .X(net4147));
 sg13g2_dlygate4sd3_1 hold1888 (.A(\data_to_write[2] ),
    .X(net4148));
 sg13g2_dlygate4sd3_1 hold1889 (.A(\i_tinyqv.cpu.instr_data_start[3] ),
    .X(net4149));
 sg13g2_dlygate4sd3_1 hold1890 (.A(\data_to_write[7] ),
    .X(net4150));
 sg13g2_dlygate4sd3_1 hold1891 (.A(\i_tinyqv.cpu.i_core.i_shift.a[6] ),
    .X(net4151));
 sg13g2_dlygate4sd3_1 hold1892 (.A(\i_tinyqv.cpu.instr_write_offset[1] ),
    .X(net4152));
 sg13g2_dlygate4sd3_1 hold1893 (.A(_02580_),
    .X(net4153));
 sg13g2_dlygate4sd3_1 hold1894 (.A(\i_tinyqv.cpu.i_core.mem_op[0] ),
    .X(net4154));
 sg13g2_dlygate4sd3_1 hold1895 (.A(debug_instr_valid),
    .X(net4155));
 sg13g2_dlygate4sd3_1 hold1896 (.A(\i_tinyqv.cpu.instr_fetch_running ),
    .X(net4156));
 sg13g2_dlygate4sd3_1 hold1897 (.A(\data_to_write[0] ),
    .X(net4157));
 sg13g2_dlygate4sd3_1 hold1898 (.A(\i_tinyqv.cpu.instr_write_offset[3] ),
    .X(net4158));
 sg13g2_dlygate4sd3_1 hold1899 (.A(\i_tinyqv.cpu.i_core.i_shift.adjusted_shift_amt[0] ),
    .X(net4159));
 sg13g2_dlygate4sd3_1 hold1900 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[24] ),
    .X(net4160));
 sg13g2_dlygate4sd3_1 hold1901 (.A(\i_tinyqv.cpu.i_core.multiplier.accum[0] ),
    .X(net4161));
 sg13g2_dlygate4sd3_1 hold1902 (.A(\i_peripherals.i_user_peri39.stage1_math_rec[23] ),
    .X(net4162));
 sg13g2_dlygate4sd3_1 hold1903 (.A(\i_tinyqv.cpu.alu_op[2] ),
    .X(net4163));
 sg13g2_dlygate4sd3_1 hold1904 (.A(\i_peripherals.i_user_peri39.busy_counter[1] ),
    .X(net4164));
 sg13g2_dlygate4sd3_1 hold1905 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[0] ),
    .X(net4165));
 sg13g2_dlygate4sd3_1 hold1906 (.A(\i_tinyqv.cpu.i_core.i_registers.rd[3] ),
    .X(net4166));
 sg13g2_dlygate4sd3_1 hold1907 (.A(_02400_),
    .X(net4167));
 sg13g2_dlygate4sd3_1 hold1908 (.A(\i_peripherals.i_user_peri39.busy_counter[2] ),
    .X(net4168));
 sg13g2_dlygate4sd3_1 hold1909 (.A(\time_count[1] ),
    .X(net4169));
 sg13g2_dlygate4sd3_1 hold1910 (.A(\i_peripherals.i_uart.i_uart_tx.cycle_counter[2] ),
    .X(net4170));
 sg13g2_dlygate4sd3_1 hold1911 (.A(\i_peripherals.i_user_peri39.busy_counter[2] ),
    .X(net4171));
 sg13g2_antennanp ANTENNA_1 (.A(net2739));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_69 ();
 sg13g2_fill_2 FILLER_0_76 ();
 sg13g2_decap_4 FILLER_0_83 ();
 sg13g2_fill_1 FILLER_0_87 ();
 sg13g2_fill_2 FILLER_0_115 ();
 sg13g2_fill_1 FILLER_0_117 ();
 sg13g2_decap_4 FILLER_0_125 ();
 sg13g2_fill_2 FILLER_0_129 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_fill_1 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_170 ();
 sg13g2_decap_8 FILLER_0_177 ();
 sg13g2_decap_8 FILLER_0_184 ();
 sg13g2_decap_8 FILLER_0_195 ();
 sg13g2_decap_8 FILLER_0_202 ();
 sg13g2_fill_1 FILLER_0_209 ();
 sg13g2_decap_8 FILLER_0_215 ();
 sg13g2_fill_1 FILLER_0_222 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_fill_2 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_fill_2 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_318 ();
 sg13g2_decap_4 FILLER_0_325 ();
 sg13g2_fill_2 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_4 FILLER_0_356 ();
 sg13g2_fill_2 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_decap_8 FILLER_0_373 ();
 sg13g2_fill_1 FILLER_0_380 ();
 sg13g2_fill_2 FILLER_0_408 ();
 sg13g2_fill_1 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_442 ();
 sg13g2_fill_2 FILLER_0_458 ();
 sg13g2_decap_4 FILLER_0_487 ();
 sg13g2_fill_2 FILLER_0_491 ();
 sg13g2_decap_8 FILLER_0_520 ();
 sg13g2_fill_1 FILLER_0_527 ();
 sg13g2_fill_2 FILLER_0_568 ();
 sg13g2_fill_1 FILLER_0_570 ();
 sg13g2_decap_8 FILLER_0_575 ();
 sg13g2_fill_1 FILLER_0_582 ();
 sg13g2_decap_8 FILLER_0_587 ();
 sg13g2_decap_8 FILLER_0_594 ();
 sg13g2_fill_1 FILLER_0_610 ();
 sg13g2_decap_8 FILLER_0_619 ();
 sg13g2_decap_4 FILLER_0_626 ();
 sg13g2_fill_1 FILLER_0_630 ();
 sg13g2_fill_2 FILLER_0_685 ();
 sg13g2_fill_1 FILLER_0_687 ();
 sg13g2_fill_2 FILLER_0_715 ();
 sg13g2_fill_1 FILLER_0_717 ();
 sg13g2_fill_1 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_800 ();
 sg13g2_decap_8 FILLER_0_807 ();
 sg13g2_fill_1 FILLER_0_814 ();
 sg13g2_decap_8 FILLER_0_873 ();
 sg13g2_decap_8 FILLER_0_880 ();
 sg13g2_fill_2 FILLER_0_887 ();
 sg13g2_decap_8 FILLER_0_893 ();
 sg13g2_decap_8 FILLER_0_900 ();
 sg13g2_decap_4 FILLER_0_907 ();
 sg13g2_fill_2 FILLER_0_911 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_4 FILLER_0_924 ();
 sg13g2_fill_2 FILLER_0_928 ();
 sg13g2_fill_2 FILLER_0_984 ();
 sg13g2_decap_8 FILLER_0_990 ();
 sg13g2_decap_8 FILLER_0_997 ();
 sg13g2_fill_2 FILLER_0_1004 ();
 sg13g2_fill_1 FILLER_0_1006 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_fill_1 FILLER_0_1049 ();
 sg13g2_fill_2 FILLER_0_1117 ();
 sg13g2_fill_2 FILLER_0_1146 ();
 sg13g2_fill_1 FILLER_0_1148 ();
 sg13g2_fill_1 FILLER_0_1176 ();
 sg13g2_fill_2 FILLER_0_1226 ();
 sg13g2_fill_1 FILLER_0_1228 ();
 sg13g2_decap_8 FILLER_0_1233 ();
 sg13g2_fill_2 FILLER_0_1240 ();
 sg13g2_decap_4 FILLER_0_1269 ();
 sg13g2_fill_1 FILLER_0_1273 ();
 sg13g2_fill_2 FILLER_0_1283 ();
 sg13g2_decap_8 FILLER_0_1298 ();
 sg13g2_fill_1 FILLER_0_1305 ();
 sg13g2_fill_1 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_decap_8 FILLER_0_1358 ();
 sg13g2_decap_4 FILLER_0_1365 ();
 sg13g2_fill_2 FILLER_0_1369 ();
 sg13g2_fill_2 FILLER_0_1469 ();
 sg13g2_fill_2 FILLER_0_1507 ();
 sg13g2_decap_8 FILLER_0_1531 ();
 sg13g2_decap_8 FILLER_0_1538 ();
 sg13g2_decap_8 FILLER_0_1545 ();
 sg13g2_decap_8 FILLER_0_1552 ();
 sg13g2_decap_8 FILLER_0_1559 ();
 sg13g2_decap_8 FILLER_0_1566 ();
 sg13g2_decap_8 FILLER_0_1573 ();
 sg13g2_decap_8 FILLER_0_1580 ();
 sg13g2_decap_8 FILLER_0_1587 ();
 sg13g2_decap_8 FILLER_0_1594 ();
 sg13g2_decap_8 FILLER_0_1601 ();
 sg13g2_decap_8 FILLER_0_1608 ();
 sg13g2_decap_8 FILLER_0_1615 ();
 sg13g2_decap_8 FILLER_0_1622 ();
 sg13g2_decap_8 FILLER_0_1629 ();
 sg13g2_decap_8 FILLER_0_1636 ();
 sg13g2_decap_8 FILLER_0_1643 ();
 sg13g2_decap_8 FILLER_0_1650 ();
 sg13g2_decap_8 FILLER_0_1657 ();
 sg13g2_decap_8 FILLER_0_1664 ();
 sg13g2_decap_8 FILLER_0_1671 ();
 sg13g2_decap_8 FILLER_0_1678 ();
 sg13g2_decap_8 FILLER_0_1685 ();
 sg13g2_decap_8 FILLER_0_1692 ();
 sg13g2_decap_8 FILLER_0_1699 ();
 sg13g2_decap_8 FILLER_0_1706 ();
 sg13g2_decap_8 FILLER_0_1713 ();
 sg13g2_decap_8 FILLER_0_1720 ();
 sg13g2_decap_8 FILLER_0_1727 ();
 sg13g2_decap_8 FILLER_0_1734 ();
 sg13g2_decap_8 FILLER_0_1741 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_decap_4 FILLER_0_1762 ();
 sg13g2_fill_2 FILLER_0_1766 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_4 FILLER_1_28 ();
 sg13g2_fill_2 FILLER_1_45 ();
 sg13g2_decap_8 FILLER_1_51 ();
 sg13g2_fill_2 FILLER_1_58 ();
 sg13g2_fill_1 FILLER_1_60 ();
 sg13g2_decap_4 FILLER_1_88 ();
 sg13g2_fill_1 FILLER_1_92 ();
 sg13g2_decap_8 FILLER_1_97 ();
 sg13g2_decap_8 FILLER_1_109 ();
 sg13g2_decap_4 FILLER_1_132 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_fill_2 FILLER_1_147 ();
 sg13g2_fill_1 FILLER_1_149 ();
 sg13g2_fill_1 FILLER_1_227 ();
 sg13g2_decap_8 FILLER_1_232 ();
 sg13g2_decap_8 FILLER_1_239 ();
 sg13g2_fill_2 FILLER_1_259 ();
 sg13g2_fill_1 FILLER_1_261 ();
 sg13g2_fill_2 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_fill_2 FILLER_1_322 ();
 sg13g2_fill_1 FILLER_1_324 ();
 sg13g2_decap_4 FILLER_1_352 ();
 sg13g2_fill_2 FILLER_1_392 ();
 sg13g2_fill_2 FILLER_1_419 ();
 sg13g2_fill_1 FILLER_1_431 ();
 sg13g2_decap_4 FILLER_1_459 ();
 sg13g2_fill_1 FILLER_1_463 ();
 sg13g2_decap_8 FILLER_1_472 ();
 sg13g2_fill_2 FILLER_1_479 ();
 sg13g2_decap_8 FILLER_1_485 ();
 sg13g2_fill_1 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_537 ();
 sg13g2_decap_8 FILLER_1_544 ();
 sg13g2_fill_1 FILLER_1_641 ();
 sg13g2_fill_2 FILLER_1_651 ();
 sg13g2_fill_1 FILLER_1_653 ();
 sg13g2_fill_2 FILLER_1_667 ();
 sg13g2_fill_2 FILLER_1_678 ();
 sg13g2_fill_1 FILLER_1_680 ();
 sg13g2_fill_1 FILLER_1_734 ();
 sg13g2_decap_8 FILLER_1_765 ();
 sg13g2_fill_1 FILLER_1_772 ();
 sg13g2_fill_2 FILLER_1_786 ();
 sg13g2_fill_1 FILLER_1_788 ();
 sg13g2_fill_1 FILLER_1_825 ();
 sg13g2_fill_2 FILLER_1_830 ();
 sg13g2_fill_1 FILLER_1_832 ();
 sg13g2_fill_2 FILLER_1_855 ();
 sg13g2_decap_8 FILLER_1_947 ();
 sg13g2_fill_1 FILLER_1_954 ();
 sg13g2_decap_4 FILLER_1_972 ();
 sg13g2_fill_1 FILLER_1_976 ();
 sg13g2_fill_2 FILLER_1_1044 ();
 sg13g2_fill_1 FILLER_1_1046 ();
 sg13g2_fill_1 FILLER_1_1074 ();
 sg13g2_fill_2 FILLER_1_1097 ();
 sg13g2_fill_1 FILLER_1_1099 ();
 sg13g2_decap_4 FILLER_1_1136 ();
 sg13g2_fill_2 FILLER_1_1166 ();
 sg13g2_fill_1 FILLER_1_1168 ();
 sg13g2_decap_4 FILLER_1_1199 ();
 sg13g2_fill_1 FILLER_1_1257 ();
 sg13g2_fill_1 FILLER_1_1338 ();
 sg13g2_fill_1 FILLER_1_1366 ();
 sg13g2_fill_1 FILLER_1_1394 ();
 sg13g2_decap_4 FILLER_1_1417 ();
 sg13g2_fill_1 FILLER_1_1421 ();
 sg13g2_decap_8 FILLER_1_1444 ();
 sg13g2_fill_1 FILLER_1_1451 ();
 sg13g2_fill_2 FILLER_1_1488 ();
 sg13g2_fill_1 FILLER_1_1517 ();
 sg13g2_fill_2 FILLER_1_1545 ();
 sg13g2_fill_1 FILLER_1_1547 ();
 sg13g2_decap_8 FILLER_1_1552 ();
 sg13g2_decap_8 FILLER_1_1559 ();
 sg13g2_decap_4 FILLER_1_1566 ();
 sg13g2_decap_8 FILLER_1_1579 ();
 sg13g2_decap_8 FILLER_1_1586 ();
 sg13g2_decap_8 FILLER_1_1593 ();
 sg13g2_decap_8 FILLER_1_1600 ();
 sg13g2_decap_8 FILLER_1_1607 ();
 sg13g2_decap_8 FILLER_1_1614 ();
 sg13g2_decap_8 FILLER_1_1621 ();
 sg13g2_decap_8 FILLER_1_1628 ();
 sg13g2_decap_8 FILLER_1_1635 ();
 sg13g2_decap_8 FILLER_1_1642 ();
 sg13g2_decap_8 FILLER_1_1649 ();
 sg13g2_decap_8 FILLER_1_1656 ();
 sg13g2_decap_8 FILLER_1_1663 ();
 sg13g2_decap_8 FILLER_1_1670 ();
 sg13g2_decap_8 FILLER_1_1677 ();
 sg13g2_decap_8 FILLER_1_1684 ();
 sg13g2_decap_8 FILLER_1_1691 ();
 sg13g2_decap_8 FILLER_1_1698 ();
 sg13g2_decap_8 FILLER_1_1705 ();
 sg13g2_decap_8 FILLER_1_1712 ();
 sg13g2_decap_8 FILLER_1_1719 ();
 sg13g2_decap_8 FILLER_1_1726 ();
 sg13g2_decap_8 FILLER_1_1733 ();
 sg13g2_decap_8 FILLER_1_1740 ();
 sg13g2_decap_8 FILLER_1_1747 ();
 sg13g2_decap_8 FILLER_1_1754 ();
 sg13g2_decap_8 FILLER_1_1761 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_4 ();
 sg13g2_decap_4 FILLER_2_49 ();
 sg13g2_fill_2 FILLER_2_53 ();
 sg13g2_fill_2 FILLER_2_76 ();
 sg13g2_decap_8 FILLER_2_87 ();
 sg13g2_fill_1 FILLER_2_94 ();
 sg13g2_decap_8 FILLER_2_115 ();
 sg13g2_fill_1 FILLER_2_122 ();
 sg13g2_fill_1 FILLER_2_128 ();
 sg13g2_decap_4 FILLER_2_134 ();
 sg13g2_fill_2 FILLER_2_138 ();
 sg13g2_decap_4 FILLER_2_160 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_fill_2 FILLER_2_216 ();
 sg13g2_fill_1 FILLER_2_218 ();
 sg13g2_decap_8 FILLER_2_236 ();
 sg13g2_decap_8 FILLER_2_243 ();
 sg13g2_decap_4 FILLER_2_250 ();
 sg13g2_fill_2 FILLER_2_274 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_4 FILLER_2_287 ();
 sg13g2_fill_2 FILLER_2_311 ();
 sg13g2_fill_2 FILLER_2_318 ();
 sg13g2_fill_1 FILLER_2_320 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_decap_4 FILLER_2_332 ();
 sg13g2_decap_8 FILLER_2_352 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_4 FILLER_2_377 ();
 sg13g2_fill_2 FILLER_2_416 ();
 sg13g2_fill_2 FILLER_2_441 ();
 sg13g2_fill_2 FILLER_2_452 ();
 sg13g2_fill_1 FILLER_2_454 ();
 sg13g2_fill_2 FILLER_2_460 ();
 sg13g2_fill_1 FILLER_2_462 ();
 sg13g2_fill_1 FILLER_2_499 ();
 sg13g2_decap_4 FILLER_2_518 ();
 sg13g2_fill_2 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_fill_2 FILLER_2_536 ();
 sg13g2_fill_1 FILLER_2_538 ();
 sg13g2_fill_2 FILLER_2_696 ();
 sg13g2_fill_1 FILLER_2_698 ();
 sg13g2_decap_4 FILLER_2_780 ();
 sg13g2_decap_4 FILLER_2_860 ();
 sg13g2_fill_1 FILLER_2_864 ();
 sg13g2_decap_4 FILLER_2_878 ();
 sg13g2_fill_2 FILLER_2_882 ();
 sg13g2_fill_2 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_899 ();
 sg13g2_fill_2 FILLER_2_906 ();
 sg13g2_decap_4 FILLER_2_943 ();
 sg13g2_fill_2 FILLER_2_947 ();
 sg13g2_fill_2 FILLER_2_980 ();
 sg13g2_fill_1 FILLER_2_982 ();
 sg13g2_decap_4 FILLER_2_992 ();
 sg13g2_fill_2 FILLER_2_996 ();
 sg13g2_fill_2 FILLER_2_1073 ();
 sg13g2_fill_1 FILLER_2_1075 ();
 sg13g2_decap_8 FILLER_2_1116 ();
 sg13g2_decap_4 FILLER_2_1123 ();
 sg13g2_decap_8 FILLER_2_1131 ();
 sg13g2_decap_4 FILLER_2_1138 ();
 sg13g2_decap_8 FILLER_2_1223 ();
 sg13g2_fill_1 FILLER_2_1239 ();
 sg13g2_fill_2 FILLER_2_1262 ();
 sg13g2_fill_1 FILLER_2_1264 ();
 sg13g2_fill_2 FILLER_2_1292 ();
 sg13g2_decap_8 FILLER_2_1386 ();
 sg13g2_fill_2 FILLER_2_1393 ();
 sg13g2_decap_8 FILLER_2_1462 ();
 sg13g2_decap_8 FILLER_2_1469 ();
 sg13g2_fill_1 FILLER_2_1476 ();
 sg13g2_decap_4 FILLER_2_1481 ();
 sg13g2_fill_1 FILLER_2_1485 ();
 sg13g2_fill_2 FILLER_2_1490 ();
 sg13g2_fill_1 FILLER_2_1492 ();
 sg13g2_fill_1 FILLER_2_1520 ();
 sg13g2_fill_1 FILLER_2_1525 ();
 sg13g2_decap_8 FILLER_2_1535 ();
 sg13g2_fill_1 FILLER_2_1542 ();
 sg13g2_decap_8 FILLER_2_1606 ();
 sg13g2_decap_8 FILLER_2_1613 ();
 sg13g2_decap_8 FILLER_2_1620 ();
 sg13g2_decap_8 FILLER_2_1627 ();
 sg13g2_decap_8 FILLER_2_1634 ();
 sg13g2_decap_8 FILLER_2_1641 ();
 sg13g2_decap_8 FILLER_2_1648 ();
 sg13g2_decap_8 FILLER_2_1655 ();
 sg13g2_decap_8 FILLER_2_1662 ();
 sg13g2_decap_8 FILLER_2_1669 ();
 sg13g2_decap_8 FILLER_2_1676 ();
 sg13g2_decap_8 FILLER_2_1683 ();
 sg13g2_decap_8 FILLER_2_1690 ();
 sg13g2_decap_8 FILLER_2_1697 ();
 sg13g2_decap_8 FILLER_2_1704 ();
 sg13g2_decap_8 FILLER_2_1711 ();
 sg13g2_decap_8 FILLER_2_1718 ();
 sg13g2_decap_8 FILLER_2_1725 ();
 sg13g2_decap_8 FILLER_2_1732 ();
 sg13g2_decap_8 FILLER_2_1739 ();
 sg13g2_decap_8 FILLER_2_1746 ();
 sg13g2_decap_8 FILLER_2_1753 ();
 sg13g2_decap_8 FILLER_2_1760 ();
 sg13g2_fill_1 FILLER_2_1767 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_fill_2 FILLER_3_32 ();
 sg13g2_fill_1 FILLER_3_34 ();
 sg13g2_decap_8 FILLER_3_43 ();
 sg13g2_decap_4 FILLER_3_50 ();
 sg13g2_decap_8 FILLER_3_66 ();
 sg13g2_decap_4 FILLER_3_93 ();
 sg13g2_fill_2 FILLER_3_119 ();
 sg13g2_fill_2 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_162 ();
 sg13g2_decap_8 FILLER_3_169 ();
 sg13g2_decap_4 FILLER_3_176 ();
 sg13g2_fill_1 FILLER_3_180 ();
 sg13g2_decap_8 FILLER_3_206 ();
 sg13g2_decap_4 FILLER_3_213 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_fill_2 FILLER_3_230 ();
 sg13g2_fill_1 FILLER_3_232 ();
 sg13g2_fill_2 FILLER_3_245 ();
 sg13g2_fill_1 FILLER_3_259 ();
 sg13g2_decap_4 FILLER_3_269 ();
 sg13g2_fill_2 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_348 ();
 sg13g2_decap_4 FILLER_3_355 ();
 sg13g2_fill_2 FILLER_3_426 ();
 sg13g2_fill_2 FILLER_3_442 ();
 sg13g2_fill_2 FILLER_3_502 ();
 sg13g2_fill_2 FILLER_3_509 ();
 sg13g2_fill_1 FILLER_3_511 ();
 sg13g2_fill_2 FILLER_3_534 ();
 sg13g2_fill_1 FILLER_3_544 ();
 sg13g2_fill_1 FILLER_3_599 ();
 sg13g2_fill_1 FILLER_3_614 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_fill_1 FILLER_3_652 ();
 sg13g2_decap_4 FILLER_3_657 ();
 sg13g2_decap_4 FILLER_3_687 ();
 sg13g2_fill_1 FILLER_3_691 ();
 sg13g2_fill_2 FILLER_3_710 ();
 sg13g2_fill_1 FILLER_3_712 ();
 sg13g2_fill_1 FILLER_3_726 ();
 sg13g2_decap_8 FILLER_3_822 ();
 sg13g2_decap_8 FILLER_3_855 ();
 sg13g2_fill_1 FILLER_3_862 ();
 sg13g2_decap_4 FILLER_3_957 ();
 sg13g2_decap_4 FILLER_3_970 ();
 sg13g2_fill_1 FILLER_3_1001 ();
 sg13g2_fill_2 FILLER_3_1094 ();
 sg13g2_fill_1 FILLER_3_1096 ();
 sg13g2_fill_2 FILLER_3_1101 ();
 sg13g2_decap_8 FILLER_3_1161 ();
 sg13g2_decap_8 FILLER_3_1168 ();
 sg13g2_fill_2 FILLER_3_1175 ();
 sg13g2_fill_1 FILLER_3_1177 ();
 sg13g2_fill_2 FILLER_3_1191 ();
 sg13g2_fill_1 FILLER_3_1193 ();
 sg13g2_fill_2 FILLER_3_1224 ();
 sg13g2_fill_2 FILLER_3_1297 ();
 sg13g2_fill_2 FILLER_3_1335 ();
 sg13g2_decap_8 FILLER_3_1373 ();
 sg13g2_fill_1 FILLER_3_1380 ();
 sg13g2_decap_8 FILLER_3_1394 ();
 sg13g2_fill_2 FILLER_3_1401 ();
 sg13g2_fill_1 FILLER_3_1403 ();
 sg13g2_decap_4 FILLER_3_1417 ();
 sg13g2_fill_1 FILLER_3_1421 ();
 sg13g2_fill_2 FILLER_3_1466 ();
 sg13g2_fill_1 FILLER_3_1495 ();
 sg13g2_decap_8 FILLER_3_1509 ();
 sg13g2_fill_1 FILLER_3_1543 ();
 sg13g2_decap_4 FILLER_3_1566 ();
 sg13g2_fill_2 FILLER_3_1570 ();
 sg13g2_decap_8 FILLER_3_1643 ();
 sg13g2_fill_1 FILLER_3_1650 ();
 sg13g2_decap_8 FILLER_3_1660 ();
 sg13g2_decap_8 FILLER_3_1667 ();
 sg13g2_decap_8 FILLER_3_1674 ();
 sg13g2_decap_8 FILLER_3_1681 ();
 sg13g2_decap_8 FILLER_3_1688 ();
 sg13g2_decap_8 FILLER_3_1695 ();
 sg13g2_decap_8 FILLER_3_1702 ();
 sg13g2_decap_8 FILLER_3_1709 ();
 sg13g2_decap_8 FILLER_3_1716 ();
 sg13g2_decap_8 FILLER_3_1723 ();
 sg13g2_decap_8 FILLER_3_1730 ();
 sg13g2_decap_8 FILLER_3_1737 ();
 sg13g2_decap_8 FILLER_3_1744 ();
 sg13g2_decap_8 FILLER_3_1751 ();
 sg13g2_decap_8 FILLER_3_1758 ();
 sg13g2_fill_2 FILLER_3_1765 ();
 sg13g2_fill_1 FILLER_3_1767 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_24 ();
 sg13g2_fill_1 FILLER_4_31 ();
 sg13g2_fill_2 FILLER_4_58 ();
 sg13g2_fill_1 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_66 ();
 sg13g2_decap_4 FILLER_4_73 ();
 sg13g2_fill_1 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_fill_2 FILLER_4_95 ();
 sg13g2_fill_1 FILLER_4_97 ();
 sg13g2_decap_8 FILLER_4_118 ();
 sg13g2_fill_2 FILLER_4_125 ();
 sg13g2_fill_1 FILLER_4_127 ();
 sg13g2_decap_4 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_162 ();
 sg13g2_decap_4 FILLER_4_169 ();
 sg13g2_fill_1 FILLER_4_173 ();
 sg13g2_fill_1 FILLER_4_187 ();
 sg13g2_fill_2 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_202 ();
 sg13g2_decap_8 FILLER_4_220 ();
 sg13g2_fill_2 FILLER_4_240 ();
 sg13g2_fill_1 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_fill_2 FILLER_4_267 ();
 sg13g2_fill_1 FILLER_4_269 ();
 sg13g2_fill_2 FILLER_4_294 ();
 sg13g2_fill_1 FILLER_4_296 ();
 sg13g2_decap_4 FILLER_4_301 ();
 sg13g2_fill_2 FILLER_4_309 ();
 sg13g2_decap_8 FILLER_4_323 ();
 sg13g2_fill_2 FILLER_4_330 ();
 sg13g2_fill_1 FILLER_4_332 ();
 sg13g2_decap_4 FILLER_4_359 ();
 sg13g2_fill_2 FILLER_4_363 ();
 sg13g2_fill_2 FILLER_4_392 ();
 sg13g2_fill_1 FILLER_4_394 ();
 sg13g2_fill_2 FILLER_4_422 ();
 sg13g2_decap_4 FILLER_4_438 ();
 sg13g2_fill_2 FILLER_4_452 ();
 sg13g2_fill_2 FILLER_4_465 ();
 sg13g2_fill_1 FILLER_4_467 ();
 sg13g2_fill_1 FILLER_4_477 ();
 sg13g2_fill_2 FILLER_4_492 ();
 sg13g2_decap_4 FILLER_4_516 ();
 sg13g2_fill_1 FILLER_4_540 ();
 sg13g2_fill_1 FILLER_4_554 ();
 sg13g2_decap_8 FILLER_4_564 ();
 sg13g2_fill_2 FILLER_4_617 ();
 sg13g2_fill_1 FILLER_4_619 ();
 sg13g2_fill_1 FILLER_4_728 ();
 sg13g2_fill_2 FILLER_4_778 ();
 sg13g2_fill_1 FILLER_4_784 ();
 sg13g2_fill_2 FILLER_4_811 ();
 sg13g2_fill_1 FILLER_4_813 ();
 sg13g2_fill_2 FILLER_4_842 ();
 sg13g2_fill_1 FILLER_4_844 ();
 sg13g2_decap_4 FILLER_4_881 ();
 sg13g2_fill_1 FILLER_4_1060 ();
 sg13g2_decap_8 FILLER_4_1106 ();
 sg13g2_decap_4 FILLER_4_1113 ();
 sg13g2_fill_1 FILLER_4_1117 ();
 sg13g2_decap_8 FILLER_4_1122 ();
 sg13g2_decap_4 FILLER_4_1146 ();
 sg13g2_fill_1 FILLER_4_1150 ();
 sg13g2_fill_1 FILLER_4_1281 ();
 sg13g2_decap_8 FILLER_4_1309 ();
 sg13g2_decap_8 FILLER_4_1316 ();
 sg13g2_fill_2 FILLER_4_1323 ();
 sg13g2_fill_2 FILLER_4_1352 ();
 sg13g2_fill_1 FILLER_4_1444 ();
 sg13g2_decap_4 FILLER_4_1489 ();
 sg13g2_fill_2 FILLER_4_1493 ();
 sg13g2_decap_4 FILLER_4_1629 ();
 sg13g2_fill_1 FILLER_4_1633 ();
 sg13g2_decap_8 FILLER_4_1661 ();
 sg13g2_decap_8 FILLER_4_1668 ();
 sg13g2_decap_8 FILLER_4_1675 ();
 sg13g2_decap_8 FILLER_4_1682 ();
 sg13g2_decap_8 FILLER_4_1689 ();
 sg13g2_decap_8 FILLER_4_1696 ();
 sg13g2_decap_8 FILLER_4_1703 ();
 sg13g2_decap_8 FILLER_4_1710 ();
 sg13g2_decap_8 FILLER_4_1717 ();
 sg13g2_decap_8 FILLER_4_1724 ();
 sg13g2_decap_8 FILLER_4_1731 ();
 sg13g2_decap_8 FILLER_4_1738 ();
 sg13g2_decap_8 FILLER_4_1745 ();
 sg13g2_decap_8 FILLER_4_1752 ();
 sg13g2_decap_8 FILLER_4_1759 ();
 sg13g2_fill_2 FILLER_4_1766 ();
 sg13g2_fill_2 FILLER_5_41 ();
 sg13g2_fill_1 FILLER_5_63 ();
 sg13g2_fill_2 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_74 ();
 sg13g2_fill_2 FILLER_5_94 ();
 sg13g2_decap_4 FILLER_5_104 ();
 sg13g2_decap_4 FILLER_5_112 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_130 ();
 sg13g2_decap_4 FILLER_5_139 ();
 sg13g2_fill_2 FILLER_5_143 ();
 sg13g2_fill_1 FILLER_5_149 ();
 sg13g2_decap_4 FILLER_5_163 ();
 sg13g2_fill_2 FILLER_5_167 ();
 sg13g2_decap_8 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_5_188 ();
 sg13g2_decap_4 FILLER_5_195 ();
 sg13g2_fill_2 FILLER_5_215 ();
 sg13g2_fill_1 FILLER_5_217 ();
 sg13g2_fill_2 FILLER_5_230 ();
 sg13g2_fill_1 FILLER_5_232 ();
 sg13g2_fill_2 FILLER_5_246 ();
 sg13g2_fill_1 FILLER_5_248 ();
 sg13g2_decap_8 FILLER_5_253 ();
 sg13g2_decap_8 FILLER_5_260 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_fill_2 FILLER_5_298 ();
 sg13g2_fill_2 FILLER_5_327 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_4 FILLER_5_364 ();
 sg13g2_fill_2 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_fill_2 FILLER_5_381 ();
 sg13g2_fill_1 FILLER_5_383 ();
 sg13g2_fill_2 FILLER_5_453 ();
 sg13g2_fill_2 FILLER_5_486 ();
 sg13g2_fill_1 FILLER_5_488 ();
 sg13g2_fill_2 FILLER_5_521 ();
 sg13g2_fill_1 FILLER_5_523 ();
 sg13g2_fill_1 FILLER_5_534 ();
 sg13g2_decap_4 FILLER_5_563 ();
 sg13g2_fill_2 FILLER_5_567 ();
 sg13g2_fill_2 FILLER_5_591 ();
 sg13g2_fill_1 FILLER_5_607 ();
 sg13g2_fill_2 FILLER_5_644 ();
 sg13g2_fill_2 FILLER_5_659 ();
 sg13g2_decap_8 FILLER_5_688 ();
 sg13g2_fill_2 FILLER_5_708 ();
 sg13g2_fill_2 FILLER_5_714 ();
 sg13g2_fill_2 FILLER_5_765 ();
 sg13g2_decap_8 FILLER_5_825 ();
 sg13g2_fill_2 FILLER_5_832 ();
 sg13g2_fill_1 FILLER_5_834 ();
 sg13g2_fill_2 FILLER_5_866 ();
 sg13g2_decap_4 FILLER_5_885 ();
 sg13g2_fill_1 FILLER_5_889 ();
 sg13g2_decap_4 FILLER_5_907 ();
 sg13g2_fill_1 FILLER_5_911 ();
 sg13g2_decap_4 FILLER_5_938 ();
 sg13g2_fill_2 FILLER_5_942 ();
 sg13g2_decap_4 FILLER_5_957 ();
 sg13g2_fill_1 FILLER_5_961 ();
 sg13g2_fill_1 FILLER_5_984 ();
 sg13g2_fill_1 FILLER_5_1021 ();
 sg13g2_fill_1 FILLER_5_1049 ();
 sg13g2_fill_2 FILLER_5_1077 ();
 sg13g2_fill_1 FILLER_5_1089 ();
 sg13g2_decap_4 FILLER_5_1180 ();
 sg13g2_fill_1 FILLER_5_1184 ();
 sg13g2_decap_8 FILLER_5_1189 ();
 sg13g2_decap_4 FILLER_5_1205 ();
 sg13g2_fill_1 FILLER_5_1272 ();
 sg13g2_fill_1 FILLER_5_1290 ();
 sg13g2_fill_2 FILLER_5_1309 ();
 sg13g2_decap_4 FILLER_5_1324 ();
 sg13g2_fill_2 FILLER_5_1328 ();
 sg13g2_decap_4 FILLER_5_1334 ();
 sg13g2_fill_1 FILLER_5_1338 ();
 sg13g2_fill_1 FILLER_5_1352 ();
 sg13g2_fill_1 FILLER_5_1392 ();
 sg13g2_fill_1 FILLER_5_1406 ();
 sg13g2_fill_2 FILLER_5_1443 ();
 sg13g2_fill_1 FILLER_5_1445 ();
 sg13g2_fill_2 FILLER_5_1513 ();
 sg13g2_decap_4 FILLER_5_1554 ();
 sg13g2_fill_2 FILLER_5_1558 ();
 sg13g2_decap_4 FILLER_5_1635 ();
 sg13g2_decap_8 FILLER_5_1643 ();
 sg13g2_decap_8 FILLER_5_1650 ();
 sg13g2_decap_8 FILLER_5_1657 ();
 sg13g2_decap_8 FILLER_5_1664 ();
 sg13g2_decap_8 FILLER_5_1671 ();
 sg13g2_decap_8 FILLER_5_1678 ();
 sg13g2_decap_8 FILLER_5_1685 ();
 sg13g2_decap_8 FILLER_5_1692 ();
 sg13g2_decap_8 FILLER_5_1699 ();
 sg13g2_decap_8 FILLER_5_1706 ();
 sg13g2_decap_8 FILLER_5_1713 ();
 sg13g2_decap_8 FILLER_5_1720 ();
 sg13g2_decap_8 FILLER_5_1727 ();
 sg13g2_decap_8 FILLER_5_1734 ();
 sg13g2_decap_8 FILLER_5_1741 ();
 sg13g2_decap_8 FILLER_5_1748 ();
 sg13g2_decap_8 FILLER_5_1755 ();
 sg13g2_decap_4 FILLER_5_1762 ();
 sg13g2_fill_2 FILLER_5_1766 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_22 ();
 sg13g2_decap_8 FILLER_6_29 ();
 sg13g2_decap_4 FILLER_6_48 ();
 sg13g2_fill_1 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_69 ();
 sg13g2_decap_4 FILLER_6_76 ();
 sg13g2_fill_1 FILLER_6_80 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_4 FILLER_6_139 ();
 sg13g2_fill_1 FILLER_6_143 ();
 sg13g2_fill_1 FILLER_6_148 ();
 sg13g2_decap_4 FILLER_6_165 ();
 sg13g2_decap_4 FILLER_6_198 ();
 sg13g2_fill_1 FILLER_6_202 ();
 sg13g2_decap_8 FILLER_6_220 ();
 sg13g2_fill_1 FILLER_6_285 ();
 sg13g2_decap_4 FILLER_6_291 ();
 sg13g2_fill_1 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_300 ();
 sg13g2_decap_8 FILLER_6_307 ();
 sg13g2_decap_8 FILLER_6_314 ();
 sg13g2_decap_4 FILLER_6_321 ();
 sg13g2_decap_8 FILLER_6_355 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_fill_2 FILLER_6_369 ();
 sg13g2_fill_1 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_376 ();
 sg13g2_decap_4 FILLER_6_383 ();
 sg13g2_fill_1 FILLER_6_387 ();
 sg13g2_decap_4 FILLER_6_400 ();
 sg13g2_fill_1 FILLER_6_404 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_fill_2 FILLER_6_440 ();
 sg13g2_fill_2 FILLER_6_447 ();
 sg13g2_fill_1 FILLER_6_459 ();
 sg13g2_fill_2 FILLER_6_464 ();
 sg13g2_fill_1 FILLER_6_466 ();
 sg13g2_decap_4 FILLER_6_476 ();
 sg13g2_fill_2 FILLER_6_484 ();
 sg13g2_fill_2 FILLER_6_491 ();
 sg13g2_fill_1 FILLER_6_493 ();
 sg13g2_fill_1 FILLER_6_499 ();
 sg13g2_fill_2 FILLER_6_504 ();
 sg13g2_fill_1 FILLER_6_506 ();
 sg13g2_decap_8 FILLER_6_516 ();
 sg13g2_fill_1 FILLER_6_527 ();
 sg13g2_decap_4 FILLER_6_533 ();
 sg13g2_fill_2 FILLER_6_537 ();
 sg13g2_decap_8 FILLER_6_556 ();
 sg13g2_fill_2 FILLER_6_563 ();
 sg13g2_fill_2 FILLER_6_597 ();
 sg13g2_fill_2 FILLER_6_613 ();
 sg13g2_fill_1 FILLER_6_615 ();
 sg13g2_fill_1 FILLER_6_652 ();
 sg13g2_fill_2 FILLER_6_657 ();
 sg13g2_fill_1 FILLER_6_659 ();
 sg13g2_fill_2 FILLER_6_677 ();
 sg13g2_fill_1 FILLER_6_679 ();
 sg13g2_fill_1 FILLER_6_728 ();
 sg13g2_fill_2 FILLER_6_765 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_fill_1 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_803 ();
 sg13g2_fill_2 FILLER_6_810 ();
 sg13g2_fill_1 FILLER_6_812 ();
 sg13g2_fill_1 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_845 ();
 sg13g2_fill_2 FILLER_6_852 ();
 sg13g2_fill_1 FILLER_6_1049 ();
 sg13g2_fill_2 FILLER_6_1059 ();
 sg13g2_decap_4 FILLER_6_1111 ();
 sg13g2_fill_2 FILLER_6_1115 ();
 sg13g2_fill_1 FILLER_6_1126 ();
 sg13g2_fill_1 FILLER_6_1140 ();
 sg13g2_decap_8 FILLER_6_1173 ();
 sg13g2_fill_2 FILLER_6_1208 ();
 sg13g2_fill_2 FILLER_6_1218 ();
 sg13g2_fill_2 FILLER_6_1229 ();
 sg13g2_fill_1 FILLER_6_1231 ();
 sg13g2_fill_1 FILLER_6_1258 ();
 sg13g2_decap_4 FILLER_6_1263 ();
 sg13g2_decap_4 FILLER_6_1311 ();
 sg13g2_fill_1 FILLER_6_1342 ();
 sg13g2_fill_1 FILLER_6_1441 ();
 sg13g2_decap_4 FILLER_6_1481 ();
 sg13g2_fill_2 FILLER_6_1485 ();
 sg13g2_fill_2 FILLER_6_1577 ();
 sg13g2_fill_1 FILLER_6_1618 ();
 sg13g2_decap_8 FILLER_6_1647 ();
 sg13g2_decap_4 FILLER_6_1654 ();
 sg13g2_fill_2 FILLER_6_1658 ();
 sg13g2_decap_8 FILLER_6_1673 ();
 sg13g2_decap_8 FILLER_6_1680 ();
 sg13g2_decap_8 FILLER_6_1687 ();
 sg13g2_decap_8 FILLER_6_1694 ();
 sg13g2_decap_8 FILLER_6_1701 ();
 sg13g2_decap_8 FILLER_6_1708 ();
 sg13g2_decap_8 FILLER_6_1715 ();
 sg13g2_decap_8 FILLER_6_1722 ();
 sg13g2_decap_8 FILLER_6_1729 ();
 sg13g2_decap_8 FILLER_6_1736 ();
 sg13g2_decap_8 FILLER_6_1743 ();
 sg13g2_decap_8 FILLER_6_1750 ();
 sg13g2_decap_8 FILLER_6_1757 ();
 sg13g2_decap_4 FILLER_6_1764 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_2 ();
 sg13g2_decap_4 FILLER_7_30 ();
 sg13g2_fill_1 FILLER_7_34 ();
 sg13g2_decap_4 FILLER_7_39 ();
 sg13g2_fill_1 FILLER_7_48 ();
 sg13g2_fill_2 FILLER_7_57 ();
 sg13g2_decap_4 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_4 FILLER_7_91 ();
 sg13g2_fill_1 FILLER_7_95 ();
 sg13g2_decap_8 FILLER_7_109 ();
 sg13g2_decap_4 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_144 ();
 sg13g2_fill_1 FILLER_7_146 ();
 sg13g2_fill_2 FILLER_7_167 ();
 sg13g2_fill_2 FILLER_7_174 ();
 sg13g2_fill_1 FILLER_7_176 ();
 sg13g2_fill_2 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_204 ();
 sg13g2_decap_4 FILLER_7_211 ();
 sg13g2_fill_1 FILLER_7_215 ();
 sg13g2_decap_4 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_246 ();
 sg13g2_decap_8 FILLER_7_253 ();
 sg13g2_decap_4 FILLER_7_260 ();
 sg13g2_decap_4 FILLER_7_268 ();
 sg13g2_fill_2 FILLER_7_289 ();
 sg13g2_decap_4 FILLER_7_346 ();
 sg13g2_fill_2 FILLER_7_350 ();
 sg13g2_fill_2 FILLER_7_365 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_fill_2 FILLER_7_452 ();
 sg13g2_decap_4 FILLER_7_464 ();
 sg13g2_fill_1 FILLER_7_468 ();
 sg13g2_fill_1 FILLER_7_515 ();
 sg13g2_decap_8 FILLER_7_562 ();
 sg13g2_fill_2 FILLER_7_569 ();
 sg13g2_fill_1 FILLER_7_575 ();
 sg13g2_fill_1 FILLER_7_585 ();
 sg13g2_decap_4 FILLER_7_590 ();
 sg13g2_fill_2 FILLER_7_611 ();
 sg13g2_fill_1 FILLER_7_613 ();
 sg13g2_fill_2 FILLER_7_633 ();
 sg13g2_fill_1 FILLER_7_680 ();
 sg13g2_fill_2 FILLER_7_694 ();
 sg13g2_fill_2 FILLER_7_741 ();
 sg13g2_fill_1 FILLER_7_743 ();
 sg13g2_fill_2 FILLER_7_811 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_fill_1 FILLER_7_833 ();
 sg13g2_fill_1 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_899 ();
 sg13g2_decap_8 FILLER_7_906 ();
 sg13g2_decap_8 FILLER_7_926 ();
 sg13g2_decap_8 FILLER_7_933 ();
 sg13g2_fill_2 FILLER_7_940 ();
 sg13g2_decap_8 FILLER_7_959 ();
 sg13g2_fill_1 FILLER_7_966 ();
 sg13g2_fill_1 FILLER_7_984 ();
 sg13g2_fill_2 FILLER_7_1007 ();
 sg13g2_fill_1 FILLER_7_1009 ();
 sg13g2_decap_4 FILLER_7_1051 ();
 sg13g2_fill_2 FILLER_7_1073 ();
 sg13g2_fill_1 FILLER_7_1075 ();
 sg13g2_fill_2 FILLER_7_1117 ();
 sg13g2_fill_2 FILLER_7_1129 ();
 sg13g2_fill_2 FILLER_7_1158 ();
 sg13g2_fill_1 FILLER_7_1160 ();
 sg13g2_decap_8 FILLER_7_1192 ();
 sg13g2_decap_4 FILLER_7_1199 ();
 sg13g2_fill_2 FILLER_7_1203 ();
 sg13g2_decap_8 FILLER_7_1233 ();
 sg13g2_fill_1 FILLER_7_1240 ();
 sg13g2_decap_4 FILLER_7_1245 ();
 sg13g2_fill_1 FILLER_7_1249 ();
 sg13g2_decap_8 FILLER_7_1287 ();
 sg13g2_decap_4 FILLER_7_1294 ();
 sg13g2_fill_2 FILLER_7_1298 ();
 sg13g2_fill_2 FILLER_7_1391 ();
 sg13g2_fill_1 FILLER_7_1393 ();
 sg13g2_fill_1 FILLER_7_1430 ();
 sg13g2_decap_4 FILLER_7_1537 ();
 sg13g2_fill_1 FILLER_7_1541 ();
 sg13g2_decap_8 FILLER_7_1546 ();
 sg13g2_decap_8 FILLER_7_1553 ();
 sg13g2_decap_4 FILLER_7_1560 ();
 sg13g2_fill_1 FILLER_7_1564 ();
 sg13g2_fill_2 FILLER_7_1569 ();
 sg13g2_fill_1 FILLER_7_1571 ();
 sg13g2_fill_1 FILLER_7_1599 ();
 sg13g2_fill_1 FILLER_7_1627 ();
 sg13g2_decap_8 FILLER_7_1691 ();
 sg13g2_decap_4 FILLER_7_1698 ();
 sg13g2_fill_2 FILLER_7_1702 ();
 sg13g2_decap_8 FILLER_7_1708 ();
 sg13g2_decap_8 FILLER_7_1715 ();
 sg13g2_decap_8 FILLER_7_1722 ();
 sg13g2_decap_8 FILLER_7_1729 ();
 sg13g2_decap_8 FILLER_7_1736 ();
 sg13g2_decap_8 FILLER_7_1743 ();
 sg13g2_decap_8 FILLER_7_1750 ();
 sg13g2_decap_8 FILLER_7_1757 ();
 sg13g2_decap_4 FILLER_7_1764 ();
 sg13g2_decap_4 FILLER_8_0 ();
 sg13g2_fill_2 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_19 ();
 sg13g2_decap_4 FILLER_8_26 ();
 sg13g2_fill_1 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_47 ();
 sg13g2_fill_1 FILLER_8_54 ();
 sg13g2_decap_8 FILLER_8_68 ();
 sg13g2_fill_2 FILLER_8_75 ();
 sg13g2_decap_4 FILLER_8_93 ();
 sg13g2_decap_8 FILLER_8_101 ();
 sg13g2_decap_8 FILLER_8_108 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_decap_8 FILLER_8_121 ();
 sg13g2_fill_2 FILLER_8_128 ();
 sg13g2_decap_4 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_187 ();
 sg13g2_fill_1 FILLER_8_201 ();
 sg13g2_decap_4 FILLER_8_240 ();
 sg13g2_fill_2 FILLER_8_244 ();
 sg13g2_decap_8 FILLER_8_250 ();
 sg13g2_decap_8 FILLER_8_257 ();
 sg13g2_decap_8 FILLER_8_293 ();
 sg13g2_decap_8 FILLER_8_300 ();
 sg13g2_fill_2 FILLER_8_307 ();
 sg13g2_fill_1 FILLER_8_309 ();
 sg13g2_fill_1 FILLER_8_337 ();
 sg13g2_decap_8 FILLER_8_358 ();
 sg13g2_fill_2 FILLER_8_365 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_fill_2 FILLER_8_378 ();
 sg13g2_fill_1 FILLER_8_380 ();
 sg13g2_decap_4 FILLER_8_410 ();
 sg13g2_fill_1 FILLER_8_414 ();
 sg13g2_fill_1 FILLER_8_419 ();
 sg13g2_decap_8 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_431 ();
 sg13g2_fill_1 FILLER_8_433 ();
 sg13g2_decap_8 FILLER_8_439 ();
 sg13g2_fill_2 FILLER_8_451 ();
 sg13g2_fill_1 FILLER_8_473 ();
 sg13g2_decap_8 FILLER_8_510 ();
 sg13g2_decap_8 FILLER_8_517 ();
 sg13g2_fill_2 FILLER_8_530 ();
 sg13g2_decap_8 FILLER_8_599 ();
 sg13g2_fill_1 FILLER_8_606 ();
 sg13g2_fill_2 FILLER_8_621 ();
 sg13g2_fill_2 FILLER_8_630 ();
 sg13g2_fill_1 FILLER_8_659 ();
 sg13g2_fill_2 FILLER_8_772 ();
 sg13g2_fill_2 FILLER_8_796 ();
 sg13g2_fill_1 FILLER_8_798 ();
 sg13g2_fill_1 FILLER_8_826 ();
 sg13g2_decap_4 FILLER_8_831 ();
 sg13g2_fill_2 FILLER_8_835 ();
 sg13g2_decap_4 FILLER_8_1025 ();
 sg13g2_fill_2 FILLER_8_1060 ();
 sg13g2_decap_8 FILLER_8_1099 ();
 sg13g2_fill_2 FILLER_8_1106 ();
 sg13g2_fill_2 FILLER_8_1127 ();
 sg13g2_fill_2 FILLER_8_1143 ();
 sg13g2_decap_8 FILLER_8_1210 ();
 sg13g2_decap_4 FILLER_8_1217 ();
 sg13g2_decap_8 FILLER_8_1225 ();
 sg13g2_decap_4 FILLER_8_1232 ();
 sg13g2_fill_2 FILLER_8_1273 ();
 sg13g2_fill_1 FILLER_8_1275 ();
 sg13g2_decap_8 FILLER_8_1322 ();
 sg13g2_fill_2 FILLER_8_1342 ();
 sg13g2_fill_2 FILLER_8_1411 ();
 sg13g2_fill_1 FILLER_8_1413 ();
 sg13g2_decap_8 FILLER_8_1458 ();
 sg13g2_fill_2 FILLER_8_1465 ();
 sg13g2_fill_1 FILLER_8_1467 ();
 sg13g2_fill_1 FILLER_8_1491 ();
 sg13g2_decap_4 FILLER_8_1529 ();
 sg13g2_decap_4 FILLER_8_1581 ();
 sg13g2_fill_1 FILLER_8_1585 ();
 sg13g2_fill_2 FILLER_8_1599 ();
 sg13g2_fill_1 FILLER_8_1623 ();
 sg13g2_decap_4 FILLER_8_1649 ();
 sg13g2_fill_2 FILLER_8_1653 ();
 sg13g2_decap_8 FILLER_8_1668 ();
 sg13g2_fill_1 FILLER_8_1675 ();
 sg13g2_decap_8 FILLER_8_1712 ();
 sg13g2_decap_8 FILLER_8_1719 ();
 sg13g2_decap_8 FILLER_8_1726 ();
 sg13g2_decap_8 FILLER_8_1733 ();
 sg13g2_decap_8 FILLER_8_1740 ();
 sg13g2_decap_8 FILLER_8_1747 ();
 sg13g2_decap_8 FILLER_8_1754 ();
 sg13g2_decap_8 FILLER_8_1761 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_decap_4 FILLER_9_31 ();
 sg13g2_fill_2 FILLER_9_48 ();
 sg13g2_fill_1 FILLER_9_50 ();
 sg13g2_decap_4 FILLER_9_71 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_fill_2 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_167 ();
 sg13g2_fill_1 FILLER_9_221 ();
 sg13g2_fill_1 FILLER_9_281 ();
 sg13g2_fill_2 FILLER_9_294 ();
 sg13g2_fill_1 FILLER_9_296 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_fill_2 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_353 ();
 sg13g2_fill_2 FILLER_9_360 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_fill_2 FILLER_9_430 ();
 sg13g2_fill_1 FILLER_9_436 ();
 sg13g2_fill_2 FILLER_9_449 ();
 sg13g2_fill_2 FILLER_9_479 ();
 sg13g2_fill_2 FILLER_9_564 ();
 sg13g2_fill_1 FILLER_9_566 ();
 sg13g2_fill_2 FILLER_9_580 ();
 sg13g2_fill_1 FILLER_9_582 ();
 sg13g2_fill_2 FILLER_9_592 ();
 sg13g2_fill_1 FILLER_9_594 ();
 sg13g2_fill_2 FILLER_9_601 ();
 sg13g2_fill_1 FILLER_9_603 ();
 sg13g2_fill_1 FILLER_9_615 ();
 sg13g2_fill_2 FILLER_9_674 ();
 sg13g2_fill_2 FILLER_9_681 ();
 sg13g2_fill_2 FILLER_9_704 ();
 sg13g2_fill_1 FILLER_9_719 ();
 sg13g2_fill_2 FILLER_9_814 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_fill_1 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_decap_8 FILLER_9_914 ();
 sg13g2_decap_8 FILLER_9_930 ();
 sg13g2_fill_2 FILLER_9_937 ();
 sg13g2_fill_1 FILLER_9_939 ();
 sg13g2_decap_4 FILLER_9_962 ();
 sg13g2_fill_1 FILLER_9_966 ();
 sg13g2_fill_1 FILLER_9_1025 ();
 sg13g2_decap_4 FILLER_9_1047 ();
 sg13g2_fill_2 FILLER_9_1082 ();
 sg13g2_fill_1 FILLER_9_1084 ();
 sg13g2_fill_2 FILLER_9_1095 ();
 sg13g2_decap_8 FILLER_9_1139 ();
 sg13g2_fill_2 FILLER_9_1146 ();
 sg13g2_fill_2 FILLER_9_1198 ();
 sg13g2_fill_1 FILLER_9_1200 ();
 sg13g2_decap_4 FILLER_9_1211 ();
 sg13g2_fill_1 FILLER_9_1215 ();
 sg13g2_fill_2 FILLER_9_1261 ();
 sg13g2_fill_2 FILLER_9_1299 ();
 sg13g2_fill_1 FILLER_9_1301 ();
 sg13g2_fill_2 FILLER_9_1329 ();
 sg13g2_decap_4 FILLER_9_1392 ();
 sg13g2_fill_2 FILLER_9_1409 ();
 sg13g2_fill_1 FILLER_9_1411 ();
 sg13g2_fill_1 FILLER_9_1433 ();
 sg13g2_decap_8 FILLER_9_1465 ();
 sg13g2_fill_1 FILLER_9_1472 ();
 sg13g2_fill_1 FILLER_9_1527 ();
 sg13g2_decap_4 FILLER_9_1555 ();
 sg13g2_fill_2 FILLER_9_1676 ();
 sg13g2_fill_1 FILLER_9_1678 ();
 sg13g2_decap_8 FILLER_9_1692 ();
 sg13g2_decap_8 FILLER_9_1726 ();
 sg13g2_decap_8 FILLER_9_1733 ();
 sg13g2_decap_8 FILLER_9_1740 ();
 sg13g2_decap_8 FILLER_9_1747 ();
 sg13g2_decap_8 FILLER_9_1754 ();
 sg13g2_decap_8 FILLER_9_1761 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_4 FILLER_10_56 ();
 sg13g2_fill_1 FILLER_10_60 ();
 sg13g2_decap_4 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_79 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_4 FILLER_10_98 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_113 ();
 sg13g2_fill_2 FILLER_10_120 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_194 ();
 sg13g2_decap_8 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_291 ();
 sg13g2_fill_2 FILLER_10_323 ();
 sg13g2_decap_4 FILLER_10_352 ();
 sg13g2_fill_2 FILLER_10_356 ();
 sg13g2_decap_4 FILLER_10_371 ();
 sg13g2_fill_1 FILLER_10_375 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_10_422 ();
 sg13g2_decap_8 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_10_436 ();
 sg13g2_fill_2 FILLER_10_443 ();
 sg13g2_fill_2 FILLER_10_450 ();
 sg13g2_fill_1 FILLER_10_460 ();
 sg13g2_decap_8 FILLER_10_467 ();
 sg13g2_decap_8 FILLER_10_474 ();
 sg13g2_decap_8 FILLER_10_481 ();
 sg13g2_fill_2 FILLER_10_488 ();
 sg13g2_fill_2 FILLER_10_506 ();
 sg13g2_fill_1 FILLER_10_508 ();
 sg13g2_fill_2 FILLER_10_517 ();
 sg13g2_fill_1 FILLER_10_580 ();
 sg13g2_fill_1 FILLER_10_603 ();
 sg13g2_fill_1 FILLER_10_615 ();
 sg13g2_decap_4 FILLER_10_620 ();
 sg13g2_fill_1 FILLER_10_624 ();
 sg13g2_decap_8 FILLER_10_642 ();
 sg13g2_decap_4 FILLER_10_649 ();
 sg13g2_fill_2 FILLER_10_667 ();
 sg13g2_fill_2 FILLER_10_746 ();
 sg13g2_fill_1 FILLER_10_748 ();
 sg13g2_fill_1 FILLER_10_775 ();
 sg13g2_fill_2 FILLER_10_834 ();
 sg13g2_fill_1 FILLER_10_836 ();
 sg13g2_decap_8 FILLER_10_859 ();
 sg13g2_fill_1 FILLER_10_866 ();
 sg13g2_fill_1 FILLER_10_975 ();
 sg13g2_decap_4 FILLER_10_994 ();
 sg13g2_decap_8 FILLER_10_1100 ();
 sg13g2_decap_4 FILLER_10_1111 ();
 sg13g2_fill_2 FILLER_10_1115 ();
 sg13g2_decap_4 FILLER_10_1127 ();
 sg13g2_decap_8 FILLER_10_1140 ();
 sg13g2_decap_8 FILLER_10_1147 ();
 sg13g2_fill_2 FILLER_10_1154 ();
 sg13g2_fill_1 FILLER_10_1156 ();
 sg13g2_decap_8 FILLER_10_1170 ();
 sg13g2_decap_4 FILLER_10_1177 ();
 sg13g2_fill_1 FILLER_10_1181 ();
 sg13g2_decap_8 FILLER_10_1206 ();
 sg13g2_decap_8 FILLER_10_1213 ();
 sg13g2_decap_8 FILLER_10_1220 ();
 sg13g2_decap_8 FILLER_10_1227 ();
 sg13g2_decap_8 FILLER_10_1234 ();
 sg13g2_decap_4 FILLER_10_1241 ();
 sg13g2_fill_2 FILLER_10_1245 ();
 sg13g2_fill_1 FILLER_10_1279 ();
 sg13g2_decap_8 FILLER_10_1299 ();
 sg13g2_fill_1 FILLER_10_1306 ();
 sg13g2_decap_8 FILLER_10_1311 ();
 sg13g2_decap_4 FILLER_10_1318 ();
 sg13g2_decap_8 FILLER_10_1326 ();
 sg13g2_fill_2 FILLER_10_1333 ();
 sg13g2_fill_1 FILLER_10_1335 ();
 sg13g2_decap_8 FILLER_10_1340 ();
 sg13g2_fill_1 FILLER_10_1347 ();
 sg13g2_decap_4 FILLER_10_1385 ();
 sg13g2_fill_2 FILLER_10_1474 ();
 sg13g2_fill_1 FILLER_10_1476 ();
 sg13g2_fill_2 FILLER_10_1517 ();
 sg13g2_fill_1 FILLER_10_1523 ();
 sg13g2_decap_8 FILLER_10_1528 ();
 sg13g2_fill_2 FILLER_10_1535 ();
 sg13g2_fill_2 FILLER_10_1573 ();
 sg13g2_fill_1 FILLER_10_1575 ();
 sg13g2_fill_1 FILLER_10_1621 ();
 sg13g2_fill_2 FILLER_10_1649 ();
 sg13g2_fill_1 FILLER_10_1655 ();
 sg13g2_decap_8 FILLER_10_1711 ();
 sg13g2_decap_8 FILLER_10_1718 ();
 sg13g2_decap_8 FILLER_10_1725 ();
 sg13g2_decap_8 FILLER_10_1732 ();
 sg13g2_decap_8 FILLER_10_1739 ();
 sg13g2_decap_8 FILLER_10_1746 ();
 sg13g2_decap_8 FILLER_10_1753 ();
 sg13g2_decap_8 FILLER_10_1760 ();
 sg13g2_fill_1 FILLER_10_1767 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_28 ();
 sg13g2_fill_1 FILLER_11_54 ();
 sg13g2_decap_8 FILLER_11_80 ();
 sg13g2_fill_2 FILLER_11_87 ();
 sg13g2_fill_2 FILLER_11_94 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_fill_2 FILLER_11_114 ();
 sg13g2_fill_1 FILLER_11_116 ();
 sg13g2_fill_2 FILLER_11_144 ();
 sg13g2_fill_2 FILLER_11_159 ();
 sg13g2_fill_1 FILLER_11_161 ();
 sg13g2_decap_4 FILLER_11_178 ();
 sg13g2_fill_2 FILLER_11_211 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_255 ();
 sg13g2_decap_8 FILLER_11_274 ();
 sg13g2_decap_8 FILLER_11_281 ();
 sg13g2_decap_8 FILLER_11_288 ();
 sg13g2_decap_8 FILLER_11_295 ();
 sg13g2_fill_2 FILLER_11_302 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_decap_4 FILLER_11_309 ();
 sg13g2_fill_2 FILLER_11_313 ();
 sg13g2_decap_4 FILLER_11_355 ();
 sg13g2_fill_1 FILLER_11_359 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_fill_1 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_414 ();
 sg13g2_fill_2 FILLER_11_421 ();
 sg13g2_fill_1 FILLER_11_435 ();
 sg13g2_decap_4 FILLER_11_447 ();
 sg13g2_fill_1 FILLER_11_451 ();
 sg13g2_decap_4 FILLER_11_497 ();
 sg13g2_fill_1 FILLER_11_501 ();
 sg13g2_fill_2 FILLER_11_507 ();
 sg13g2_fill_2 FILLER_11_515 ();
 sg13g2_fill_1 FILLER_11_543 ();
 sg13g2_fill_2 FILLER_11_558 ();
 sg13g2_fill_1 FILLER_11_560 ();
 sg13g2_fill_1 FILLER_11_601 ();
 sg13g2_decap_4 FILLER_11_638 ();
 sg13g2_fill_1 FILLER_11_642 ();
 sg13g2_fill_1 FILLER_11_675 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_fill_1 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_fill_2 FILLER_11_725 ();
 sg13g2_fill_2 FILLER_11_754 ();
 sg13g2_fill_2 FILLER_11_792 ();
 sg13g2_decap_8 FILLER_11_853 ();
 sg13g2_decap_4 FILLER_11_860 ();
 sg13g2_fill_1 FILLER_11_864 ();
 sg13g2_decap_8 FILLER_11_869 ();
 sg13g2_fill_1 FILLER_11_880 ();
 sg13g2_decap_8 FILLER_11_890 ();
 sg13g2_decap_8 FILLER_11_897 ();
 sg13g2_decap_8 FILLER_11_904 ();
 sg13g2_decap_4 FILLER_11_911 ();
 sg13g2_fill_2 FILLER_11_946 ();
 sg13g2_fill_1 FILLER_11_948 ();
 sg13g2_decap_8 FILLER_11_1143 ();
 sg13g2_decap_4 FILLER_11_1150 ();
 sg13g2_fill_2 FILLER_11_1154 ();
 sg13g2_decap_8 FILLER_11_1167 ();
 sg13g2_decap_8 FILLER_11_1174 ();
 sg13g2_decap_4 FILLER_11_1181 ();
 sg13g2_decap_8 FILLER_11_1191 ();
 sg13g2_decap_8 FILLER_11_1198 ();
 sg13g2_decap_4 FILLER_11_1205 ();
 sg13g2_decap_4 FILLER_11_1215 ();
 sg13g2_fill_1 FILLER_11_1219 ();
 sg13g2_decap_8 FILLER_11_1226 ();
 sg13g2_fill_1 FILLER_11_1233 ();
 sg13g2_decap_8 FILLER_11_1240 ();
 sg13g2_decap_8 FILLER_11_1247 ();
 sg13g2_decap_4 FILLER_11_1254 ();
 sg13g2_fill_2 FILLER_11_1290 ();
 sg13g2_fill_1 FILLER_11_1292 ();
 sg13g2_fill_1 FILLER_11_1348 ();
 sg13g2_fill_2 FILLER_11_1359 ();
 sg13g2_fill_1 FILLER_11_1392 ();
 sg13g2_fill_2 FILLER_11_1436 ();
 sg13g2_fill_2 FILLER_11_1456 ();
 sg13g2_fill_1 FILLER_11_1458 ();
 sg13g2_fill_1 FILLER_11_1513 ();
 sg13g2_decap_4 FILLER_11_1550 ();
 sg13g2_fill_2 FILLER_11_1554 ();
 sg13g2_fill_2 FILLER_11_1584 ();
 sg13g2_fill_1 FILLER_11_1586 ();
 sg13g2_fill_2 FILLER_11_1596 ();
 sg13g2_fill_1 FILLER_11_1598 ();
 sg13g2_fill_1 FILLER_11_1608 ();
 sg13g2_fill_1 FILLER_11_1677 ();
 sg13g2_fill_2 FILLER_11_1691 ();
 sg13g2_decap_8 FILLER_11_1720 ();
 sg13g2_decap_8 FILLER_11_1727 ();
 sg13g2_decap_8 FILLER_11_1734 ();
 sg13g2_decap_8 FILLER_11_1741 ();
 sg13g2_decap_8 FILLER_11_1748 ();
 sg13g2_decap_8 FILLER_11_1755 ();
 sg13g2_decap_4 FILLER_11_1762 ();
 sg13g2_fill_2 FILLER_11_1766 ();
 sg13g2_decap_4 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_4 ();
 sg13g2_fill_1 FILLER_12_19 ();
 sg13g2_fill_1 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_4 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_122 ();
 sg13g2_fill_2 FILLER_12_129 ();
 sg13g2_decap_8 FILLER_12_157 ();
 sg13g2_fill_2 FILLER_12_174 ();
 sg13g2_fill_1 FILLER_12_176 ();
 sg13g2_fill_2 FILLER_12_200 ();
 sg13g2_fill_1 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_232 ();
 sg13g2_decap_4 FILLER_12_275 ();
 sg13g2_decap_8 FILLER_12_292 ();
 sg13g2_fill_1 FILLER_12_299 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_fill_2 FILLER_12_344 ();
 sg13g2_fill_2 FILLER_12_351 ();
 sg13g2_fill_1 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_fill_1 FILLER_12_371 ();
 sg13g2_fill_2 FILLER_12_400 ();
 sg13g2_decap_8 FILLER_12_430 ();
 sg13g2_decap_4 FILLER_12_437 ();
 sg13g2_fill_1 FILLER_12_441 ();
 sg13g2_decap_8 FILLER_12_446 ();
 sg13g2_decap_8 FILLER_12_453 ();
 sg13g2_decap_8 FILLER_12_460 ();
 sg13g2_fill_2 FILLER_12_467 ();
 sg13g2_fill_2 FILLER_12_487 ();
 sg13g2_fill_2 FILLER_12_511 ();
 sg13g2_fill_1 FILLER_12_522 ();
 sg13g2_fill_2 FILLER_12_549 ();
 sg13g2_fill_1 FILLER_12_551 ();
 sg13g2_fill_2 FILLER_12_576 ();
 sg13g2_fill_1 FILLER_12_590 ();
 sg13g2_fill_1 FILLER_12_608 ();
 sg13g2_decap_8 FILLER_12_617 ();
 sg13g2_decap_8 FILLER_12_624 ();
 sg13g2_decap_4 FILLER_12_631 ();
 sg13g2_fill_2 FILLER_12_635 ();
 sg13g2_decap_4 FILLER_12_645 ();
 sg13g2_decap_8 FILLER_12_653 ();
 sg13g2_fill_2 FILLER_12_660 ();
 sg13g2_fill_2 FILLER_12_672 ();
 sg13g2_fill_1 FILLER_12_785 ();
 sg13g2_fill_1 FILLER_12_817 ();
 sg13g2_decap_8 FILLER_12_908 ();
 sg13g2_decap_4 FILLER_12_915 ();
 sg13g2_fill_1 FILLER_12_919 ();
 sg13g2_decap_4 FILLER_12_941 ();
 sg13g2_fill_2 FILLER_12_945 ();
 sg13g2_decap_4 FILLER_12_960 ();
 sg13g2_decap_4 FILLER_12_991 ();
 sg13g2_fill_2 FILLER_12_995 ();
 sg13g2_fill_1 FILLER_12_1023 ();
 sg13g2_decap_4 FILLER_12_1083 ();
 sg13g2_fill_1 FILLER_12_1087 ();
 sg13g2_decap_8 FILLER_12_1098 ();
 sg13g2_fill_2 FILLER_12_1105 ();
 sg13g2_decap_8 FILLER_12_1116 ();
 sg13g2_decap_8 FILLER_12_1123 ();
 sg13g2_decap_8 FILLER_12_1130 ();
 sg13g2_fill_2 FILLER_12_1137 ();
 sg13g2_decap_8 FILLER_12_1145 ();
 sg13g2_decap_8 FILLER_12_1152 ();
 sg13g2_decap_8 FILLER_12_1159 ();
 sg13g2_decap_8 FILLER_12_1166 ();
 sg13g2_fill_1 FILLER_12_1173 ();
 sg13g2_fill_1 FILLER_12_1180 ();
 sg13g2_decap_8 FILLER_12_1186 ();
 sg13g2_fill_2 FILLER_12_1193 ();
 sg13g2_decap_8 FILLER_12_1201 ();
 sg13g2_fill_2 FILLER_12_1220 ();
 sg13g2_decap_8 FILLER_12_1228 ();
 sg13g2_decap_8 FILLER_12_1235 ();
 sg13g2_decap_8 FILLER_12_1242 ();
 sg13g2_decap_8 FILLER_12_1249 ();
 sg13g2_decap_4 FILLER_12_1256 ();
 sg13g2_fill_1 FILLER_12_1260 ();
 sg13g2_fill_1 FILLER_12_1298 ();
 sg13g2_decap_8 FILLER_12_1318 ();
 sg13g2_decap_8 FILLER_12_1325 ();
 sg13g2_fill_1 FILLER_12_1332 ();
 sg13g2_decap_4 FILLER_12_1374 ();
 sg13g2_fill_1 FILLER_12_1378 ();
 sg13g2_fill_2 FILLER_12_1388 ();
 sg13g2_fill_2 FILLER_12_1417 ();
 sg13g2_fill_2 FILLER_12_1446 ();
 sg13g2_fill_2 FILLER_12_1484 ();
 sg13g2_fill_1 FILLER_12_1486 ();
 sg13g2_fill_2 FILLER_12_1525 ();
 sg13g2_fill_1 FILLER_12_1527 ();
 sg13g2_fill_1 FILLER_12_1541 ();
 sg13g2_fill_1 FILLER_12_1546 ();
 sg13g2_decap_8 FILLER_12_1569 ();
 sg13g2_fill_2 FILLER_12_1611 ();
 sg13g2_fill_1 FILLER_12_1613 ();
 sg13g2_fill_1 FILLER_12_1627 ();
 sg13g2_fill_1 FILLER_12_1645 ();
 sg13g2_decap_8 FILLER_12_1731 ();
 sg13g2_fill_2 FILLER_12_1765 ();
 sg13g2_fill_1 FILLER_12_1767 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_26 ();
 sg13g2_decap_8 FILLER_13_33 ();
 sg13g2_decap_4 FILLER_13_40 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_4 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_4 FILLER_13_147 ();
 sg13g2_decap_4 FILLER_13_177 ();
 sg13g2_fill_2 FILLER_13_181 ();
 sg13g2_fill_1 FILLER_13_196 ();
 sg13g2_decap_4 FILLER_13_202 ();
 sg13g2_decap_8 FILLER_13_211 ();
 sg13g2_fill_2 FILLER_13_223 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_decap_8 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_344 ();
 sg13g2_fill_1 FILLER_13_346 ();
 sg13g2_decap_4 FILLER_13_351 ();
 sg13g2_fill_1 FILLER_13_355 ();
 sg13g2_fill_2 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_376 ();
 sg13g2_decap_8 FILLER_13_381 ();
 sg13g2_fill_2 FILLER_13_388 ();
 sg13g2_fill_1 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_421 ();
 sg13g2_decap_4 FILLER_13_428 ();
 sg13g2_fill_2 FILLER_13_486 ();
 sg13g2_fill_1 FILLER_13_488 ();
 sg13g2_fill_1 FILLER_13_510 ();
 sg13g2_fill_2 FILLER_13_516 ();
 sg13g2_fill_1 FILLER_13_518 ();
 sg13g2_fill_2 FILLER_13_529 ();
 sg13g2_fill_1 FILLER_13_531 ();
 sg13g2_fill_1 FILLER_13_545 ();
 sg13g2_decap_8 FILLER_13_551 ();
 sg13g2_decap_4 FILLER_13_558 ();
 sg13g2_fill_2 FILLER_13_600 ();
 sg13g2_fill_1 FILLER_13_602 ();
 sg13g2_decap_4 FILLER_13_630 ();
 sg13g2_fill_1 FILLER_13_661 ();
 sg13g2_decap_4 FILLER_13_666 ();
 sg13g2_fill_2 FILLER_13_670 ();
 sg13g2_decap_4 FILLER_13_675 ();
 sg13g2_decap_8 FILLER_13_706 ();
 sg13g2_decap_4 FILLER_13_713 ();
 sg13g2_fill_1 FILLER_13_717 ();
 sg13g2_decap_4 FILLER_13_721 ();
 sg13g2_fill_1 FILLER_13_725 ();
 sg13g2_fill_2 FILLER_13_730 ();
 sg13g2_decap_8 FILLER_13_736 ();
 sg13g2_fill_2 FILLER_13_743 ();
 sg13g2_fill_1 FILLER_13_745 ();
 sg13g2_fill_2 FILLER_13_763 ();
 sg13g2_fill_2 FILLER_13_801 ();
 sg13g2_fill_1 FILLER_13_857 ();
 sg13g2_decap_8 FILLER_13_871 ();
 sg13g2_decap_8 FILLER_13_878 ();
 sg13g2_fill_1 FILLER_13_885 ();
 sg13g2_decap_4 FILLER_13_890 ();
 sg13g2_fill_2 FILLER_13_894 ();
 sg13g2_fill_2 FILLER_13_977 ();
 sg13g2_fill_1 FILLER_13_979 ();
 sg13g2_decap_4 FILLER_13_1038 ();
 sg13g2_fill_1 FILLER_13_1042 ();
 sg13g2_decap_8 FILLER_13_1107 ();
 sg13g2_fill_1 FILLER_13_1114 ();
 sg13g2_fill_1 FILLER_13_1126 ();
 sg13g2_fill_2 FILLER_13_1133 ();
 sg13g2_decap_8 FILLER_13_1141 ();
 sg13g2_decap_4 FILLER_13_1148 ();
 sg13g2_fill_2 FILLER_13_1152 ();
 sg13g2_decap_8 FILLER_13_1160 ();
 sg13g2_decap_8 FILLER_13_1167 ();
 sg13g2_decap_8 FILLER_13_1174 ();
 sg13g2_decap_8 FILLER_13_1186 ();
 sg13g2_decap_8 FILLER_13_1193 ();
 sg13g2_decap_8 FILLER_13_1200 ();
 sg13g2_fill_1 FILLER_13_1207 ();
 sg13g2_decap_4 FILLER_13_1219 ();
 sg13g2_fill_1 FILLER_13_1223 ();
 sg13g2_decap_4 FILLER_13_1230 ();
 sg13g2_decap_4 FILLER_13_1240 ();
 sg13g2_decap_8 FILLER_13_1248 ();
 sg13g2_decap_8 FILLER_13_1255 ();
 sg13g2_decap_4 FILLER_13_1262 ();
 sg13g2_decap_4 FILLER_13_1270 ();
 sg13g2_fill_1 FILLER_13_1291 ();
 sg13g2_fill_2 FILLER_13_1306 ();
 sg13g2_fill_1 FILLER_13_1308 ();
 sg13g2_decap_8 FILLER_13_1313 ();
 sg13g2_decap_4 FILLER_13_1320 ();
 sg13g2_fill_1 FILLER_13_1324 ();
 sg13g2_fill_2 FILLER_13_1342 ();
 sg13g2_decap_4 FILLER_13_1353 ();
 sg13g2_fill_2 FILLER_13_1402 ();
 sg13g2_fill_1 FILLER_13_1404 ();
 sg13g2_fill_2 FILLER_13_1441 ();
 sg13g2_fill_1 FILLER_13_1443 ();
 sg13g2_fill_2 FILLER_13_1466 ();
 sg13g2_fill_2 FILLER_13_1513 ();
 sg13g2_fill_1 FILLER_13_1515 ();
 sg13g2_fill_1 FILLER_13_1553 ();
 sg13g2_decap_4 FILLER_13_1567 ();
 sg13g2_fill_1 FILLER_13_1571 ();
 sg13g2_fill_2 FILLER_13_1680 ();
 sg13g2_decap_8 FILLER_13_1686 ();
 sg13g2_decap_4 FILLER_13_1693 ();
 sg13g2_fill_1 FILLER_13_1697 ();
 sg13g2_decap_8 FILLER_13_1755 ();
 sg13g2_decap_4 FILLER_13_1762 ();
 sg13g2_fill_2 FILLER_13_1766 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_4 FILLER_14_25 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_1 FILLER_14_152 ();
 sg13g2_fill_2 FILLER_14_157 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_decap_8 FILLER_14_170 ();
 sg13g2_decap_4 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_decap_4 FILLER_14_196 ();
 sg13g2_fill_2 FILLER_14_200 ();
 sg13g2_decap_4 FILLER_14_219 ();
 sg13g2_decap_8 FILLER_14_246 ();
 sg13g2_fill_2 FILLER_14_253 ();
 sg13g2_decap_8 FILLER_14_269 ();
 sg13g2_decap_4 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_280 ();
 sg13g2_fill_2 FILLER_14_295 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_fill_1 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_330 ();
 sg13g2_fill_1 FILLER_14_337 ();
 sg13g2_decap_4 FILLER_14_364 ();
 sg13g2_fill_1 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_4 FILLER_14_400 ();
 sg13g2_fill_1 FILLER_14_404 ();
 sg13g2_decap_4 FILLER_14_410 ();
 sg13g2_fill_1 FILLER_14_435 ();
 sg13g2_fill_2 FILLER_14_471 ();
 sg13g2_fill_2 FILLER_14_497 ();
 sg13g2_fill_1 FILLER_14_499 ();
 sg13g2_decap_8 FILLER_14_597 ();
 sg13g2_decap_8 FILLER_14_604 ();
 sg13g2_fill_1 FILLER_14_639 ();
 sg13g2_decap_4 FILLER_14_749 ();
 sg13g2_fill_1 FILLER_14_753 ();
 sg13g2_fill_2 FILLER_14_763 ();
 sg13g2_decap_4 FILLER_14_786 ();
 sg13g2_fill_1 FILLER_14_790 ();
 sg13g2_decap_8 FILLER_14_795 ();
 sg13g2_decap_4 FILLER_14_802 ();
 sg13g2_fill_2 FILLER_14_806 ();
 sg13g2_decap_8 FILLER_14_821 ();
 sg13g2_fill_2 FILLER_14_828 ();
 sg13g2_fill_2 FILLER_14_843 ();
 sg13g2_fill_2 FILLER_14_911 ();
 sg13g2_fill_2 FILLER_14_926 ();
 sg13g2_fill_1 FILLER_14_928 ();
 sg13g2_fill_2 FILLER_14_969 ();
 sg13g2_decap_4 FILLER_14_980 ();
 sg13g2_decap_8 FILLER_14_997 ();
 sg13g2_fill_1 FILLER_14_1030 ();
 sg13g2_fill_2 FILLER_14_1040 ();
 sg13g2_fill_1 FILLER_14_1056 ();
 sg13g2_fill_2 FILLER_14_1067 ();
 sg13g2_fill_1 FILLER_14_1069 ();
 sg13g2_decap_8 FILLER_14_1093 ();
 sg13g2_decap_8 FILLER_14_1100 ();
 sg13g2_decap_8 FILLER_14_1107 ();
 sg13g2_fill_1 FILLER_14_1114 ();
 sg13g2_decap_8 FILLER_14_1121 ();
 sg13g2_decap_8 FILLER_14_1128 ();
 sg13g2_decap_8 FILLER_14_1135 ();
 sg13g2_decap_8 FILLER_14_1142 ();
 sg13g2_fill_2 FILLER_14_1149 ();
 sg13g2_fill_1 FILLER_14_1151 ();
 sg13g2_fill_2 FILLER_14_1158 ();
 sg13g2_decap_8 FILLER_14_1166 ();
 sg13g2_decap_4 FILLER_14_1173 ();
 sg13g2_fill_2 FILLER_14_1177 ();
 sg13g2_fill_1 FILLER_14_1185 ();
 sg13g2_fill_2 FILLER_14_1192 ();
 sg13g2_fill_1 FILLER_14_1194 ();
 sg13g2_decap_8 FILLER_14_1201 ();
 sg13g2_decap_8 FILLER_14_1208 ();
 sg13g2_decap_8 FILLER_14_1215 ();
 sg13g2_fill_2 FILLER_14_1222 ();
 sg13g2_fill_1 FILLER_14_1241 ();
 sg13g2_decap_4 FILLER_14_1254 ();
 sg13g2_fill_2 FILLER_14_1258 ();
 sg13g2_decap_8 FILLER_14_1266 ();
 sg13g2_decap_4 FILLER_14_1273 ();
 sg13g2_fill_1 FILLER_14_1277 ();
 sg13g2_fill_2 FILLER_14_1423 ();
 sg13g2_fill_1 FILLER_14_1425 ();
 sg13g2_fill_1 FILLER_14_1526 ();
 sg13g2_fill_1 FILLER_14_1594 ();
 sg13g2_decap_8 FILLER_14_1692 ();
 sg13g2_fill_2 FILLER_14_1699 ();
 sg13g2_fill_1 FILLER_14_1701 ();
 sg13g2_decap_8 FILLER_14_1733 ();
 sg13g2_decap_4 FILLER_14_1740 ();
 sg13g2_fill_2 FILLER_14_1744 ();
 sg13g2_decap_8 FILLER_14_1750 ();
 sg13g2_decap_8 FILLER_14_1757 ();
 sg13g2_decap_4 FILLER_14_1764 ();
 sg13g2_fill_2 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_30 ();
 sg13g2_fill_1 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_90 ();
 sg13g2_fill_2 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_120 ();
 sg13g2_fill_1 FILLER_15_122 ();
 sg13g2_decap_4 FILLER_15_138 ();
 sg13g2_fill_1 FILLER_15_142 ();
 sg13g2_fill_1 FILLER_15_153 ();
 sg13g2_fill_2 FILLER_15_175 ();
 sg13g2_fill_2 FILLER_15_182 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_decap_8 FILLER_15_247 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_decap_4 FILLER_15_274 ();
 sg13g2_fill_1 FILLER_15_291 ();
 sg13g2_fill_1 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_fill_2 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_370 ();
 sg13g2_fill_2 FILLER_15_377 ();
 sg13g2_fill_1 FILLER_15_379 ();
 sg13g2_decap_4 FILLER_15_384 ();
 sg13g2_fill_2 FILLER_15_388 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_15_421 ();
 sg13g2_fill_1 FILLER_15_423 ();
 sg13g2_decap_8 FILLER_15_427 ();
 sg13g2_decap_4 FILLER_15_438 ();
 sg13g2_fill_1 FILLER_15_442 ();
 sg13g2_fill_2 FILLER_15_448 ();
 sg13g2_fill_2 FILLER_15_468 ();
 sg13g2_fill_1 FILLER_15_470 ();
 sg13g2_decap_4 FILLER_15_475 ();
 sg13g2_fill_2 FILLER_15_483 ();
 sg13g2_decap_4 FILLER_15_494 ();
 sg13g2_decap_8 FILLER_15_511 ();
 sg13g2_fill_2 FILLER_15_518 ();
 sg13g2_fill_1 FILLER_15_520 ();
 sg13g2_fill_2 FILLER_15_526 ();
 sg13g2_decap_8 FILLER_15_537 ();
 sg13g2_fill_2 FILLER_15_544 ();
 sg13g2_fill_1 FILLER_15_546 ();
 sg13g2_decap_4 FILLER_15_560 ();
 sg13g2_fill_1 FILLER_15_564 ();
 sg13g2_decap_4 FILLER_15_575 ();
 sg13g2_fill_2 FILLER_15_579 ();
 sg13g2_decap_8 FILLER_15_594 ();
 sg13g2_decap_8 FILLER_15_601 ();
 sg13g2_decap_8 FILLER_15_608 ();
 sg13g2_fill_2 FILLER_15_615 ();
 sg13g2_fill_2 FILLER_15_652 ();
 sg13g2_fill_1 FILLER_15_654 ();
 sg13g2_fill_2 FILLER_15_673 ();
 sg13g2_decap_4 FILLER_15_688 ();
 sg13g2_fill_1 FILLER_15_692 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_fill_2 FILLER_15_741 ();
 sg13g2_fill_1 FILLER_15_748 ();
 sg13g2_decap_8 FILLER_15_763 ();
 sg13g2_decap_4 FILLER_15_770 ();
 sg13g2_decap_8 FILLER_15_784 ();
 sg13g2_fill_1 FILLER_15_791 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_4 FILLER_15_809 ();
 sg13g2_fill_1 FILLER_15_818 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_4 FILLER_15_835 ();
 sg13g2_fill_1 FILLER_15_839 ();
 sg13g2_fill_1 FILLER_15_846 ();
 sg13g2_decap_8 FILLER_15_854 ();
 sg13g2_decap_8 FILLER_15_861 ();
 sg13g2_decap_8 FILLER_15_868 ();
 sg13g2_decap_8 FILLER_15_875 ();
 sg13g2_fill_2 FILLER_15_882 ();
 sg13g2_decap_4 FILLER_15_947 ();
 sg13g2_fill_1 FILLER_15_951 ();
 sg13g2_decap_4 FILLER_15_965 ();
 sg13g2_decap_4 FILLER_15_973 ();
 sg13g2_fill_2 FILLER_15_977 ();
 sg13g2_fill_2 FILLER_15_983 ();
 sg13g2_fill_1 FILLER_15_985 ();
 sg13g2_fill_2 FILLER_15_993 ();
 sg13g2_fill_1 FILLER_15_995 ();
 sg13g2_decap_4 FILLER_15_1012 ();
 sg13g2_fill_2 FILLER_15_1016 ();
 sg13g2_fill_1 FILLER_15_1025 ();
 sg13g2_fill_2 FILLER_15_1039 ();
 sg13g2_fill_1 FILLER_15_1041 ();
 sg13g2_fill_1 FILLER_15_1069 ();
 sg13g2_decap_8 FILLER_15_1088 ();
 sg13g2_decap_8 FILLER_15_1095 ();
 sg13g2_fill_2 FILLER_15_1102 ();
 sg13g2_fill_1 FILLER_15_1104 ();
 sg13g2_decap_8 FILLER_15_1113 ();
 sg13g2_decap_8 FILLER_15_1120 ();
 sg13g2_decap_8 FILLER_15_1127 ();
 sg13g2_decap_8 FILLER_15_1140 ();
 sg13g2_decap_8 FILLER_15_1147 ();
 sg13g2_decap_4 FILLER_15_1154 ();
 sg13g2_fill_1 FILLER_15_1158 ();
 sg13g2_decap_8 FILLER_15_1170 ();
 sg13g2_decap_4 FILLER_15_1177 ();
 sg13g2_decap_8 FILLER_15_1187 ();
 sg13g2_decap_8 FILLER_15_1194 ();
 sg13g2_fill_2 FILLER_15_1201 ();
 sg13g2_decap_8 FILLER_15_1209 ();
 sg13g2_decap_8 FILLER_15_1216 ();
 sg13g2_decap_4 FILLER_15_1223 ();
 sg13g2_fill_1 FILLER_15_1227 ();
 sg13g2_decap_8 FILLER_15_1234 ();
 sg13g2_decap_8 FILLER_15_1241 ();
 sg13g2_decap_8 FILLER_15_1248 ();
 sg13g2_decap_8 FILLER_15_1255 ();
 sg13g2_decap_8 FILLER_15_1262 ();
 sg13g2_decap_8 FILLER_15_1269 ();
 sg13g2_decap_8 FILLER_15_1276 ();
 sg13g2_fill_2 FILLER_15_1283 ();
 sg13g2_decap_8 FILLER_15_1317 ();
 sg13g2_decap_8 FILLER_15_1324 ();
 sg13g2_fill_2 FILLER_15_1331 ();
 sg13g2_fill_1 FILLER_15_1333 ();
 sg13g2_decap_4 FILLER_15_1347 ();
 sg13g2_fill_2 FILLER_15_1351 ();
 sg13g2_fill_2 FILLER_15_1429 ();
 sg13g2_fill_1 FILLER_15_1431 ();
 sg13g2_fill_2 FILLER_15_1459 ();
 sg13g2_fill_1 FILLER_15_1461 ();
 sg13g2_fill_1 FILLER_15_1504 ();
 sg13g2_fill_2 FILLER_15_1509 ();
 sg13g2_fill_1 FILLER_15_1520 ();
 sg13g2_fill_2 FILLER_15_1525 ();
 sg13g2_fill_1 FILLER_15_1527 ();
 sg13g2_decap_4 FILLER_15_1564 ();
 sg13g2_fill_2 FILLER_15_1568 ();
 sg13g2_fill_2 FILLER_15_1658 ();
 sg13g2_fill_1 FILLER_15_1660 ();
 sg13g2_fill_1 FILLER_15_1724 ();
 sg13g2_fill_2 FILLER_15_1738 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_fill_1 FILLER_16_70 ();
 sg13g2_decap_4 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_4 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_decap_4 FILLER_16_150 ();
 sg13g2_fill_1 FILLER_16_154 ();
 sg13g2_decap_4 FILLER_16_170 ();
 sg13g2_fill_1 FILLER_16_191 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_fill_2 FILLER_16_232 ();
 sg13g2_fill_1 FILLER_16_234 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_4 FILLER_16_266 ();
 sg13g2_fill_1 FILLER_16_270 ();
 sg13g2_fill_2 FILLER_16_297 ();
 sg13g2_decap_8 FILLER_16_311 ();
 sg13g2_fill_2 FILLER_16_318 ();
 sg13g2_fill_1 FILLER_16_320 ();
 sg13g2_decap_4 FILLER_16_331 ();
 sg13g2_fill_2 FILLER_16_335 ();
 sg13g2_decap_4 FILLER_16_373 ();
 sg13g2_fill_2 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_4 FILLER_16_398 ();
 sg13g2_fill_2 FILLER_16_420 ();
 sg13g2_fill_1 FILLER_16_444 ();
 sg13g2_fill_2 FILLER_16_459 ();
 sg13g2_fill_1 FILLER_16_461 ();
 sg13g2_fill_1 FILLER_16_475 ();
 sg13g2_decap_4 FILLER_16_495 ();
 sg13g2_fill_1 FILLER_16_517 ();
 sg13g2_fill_2 FILLER_16_524 ();
 sg13g2_fill_2 FILLER_16_540 ();
 sg13g2_decap_4 FILLER_16_637 ();
 sg13g2_fill_1 FILLER_16_674 ();
 sg13g2_fill_1 FILLER_16_685 ();
 sg13g2_decap_4 FILLER_16_714 ();
 sg13g2_fill_2 FILLER_16_718 ();
 sg13g2_fill_1 FILLER_16_737 ();
 sg13g2_fill_2 FILLER_16_768 ();
 sg13g2_fill_1 FILLER_16_770 ();
 sg13g2_fill_1 FILLER_16_796 ();
 sg13g2_decap_4 FILLER_16_801 ();
 sg13g2_fill_2 FILLER_16_815 ();
 sg13g2_fill_1 FILLER_16_836 ();
 sg13g2_fill_1 FILLER_16_855 ();
 sg13g2_fill_2 FILLER_16_867 ();
 sg13g2_fill_2 FILLER_16_877 ();
 sg13g2_fill_2 FILLER_16_885 ();
 sg13g2_decap_8 FILLER_16_892 ();
 sg13g2_decap_4 FILLER_16_899 ();
 sg13g2_fill_2 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_918 ();
 sg13g2_decap_8 FILLER_16_925 ();
 sg13g2_decap_4 FILLER_16_932 ();
 sg13g2_fill_2 FILLER_16_936 ();
 sg13g2_decap_4 FILLER_16_942 ();
 sg13g2_fill_1 FILLER_16_946 ();
 sg13g2_fill_2 FILLER_16_1002 ();
 sg13g2_fill_2 FILLER_16_1014 ();
 sg13g2_fill_1 FILLER_16_1016 ();
 sg13g2_fill_1 FILLER_16_1058 ();
 sg13g2_fill_2 FILLER_16_1064 ();
 sg13g2_fill_1 FILLER_16_1066 ();
 sg13g2_decap_8 FILLER_16_1087 ();
 sg13g2_decap_8 FILLER_16_1094 ();
 sg13g2_decap_8 FILLER_16_1101 ();
 sg13g2_decap_8 FILLER_16_1108 ();
 sg13g2_decap_8 FILLER_16_1115 ();
 sg13g2_decap_4 FILLER_16_1122 ();
 sg13g2_fill_1 FILLER_16_1126 ();
 sg13g2_decap_8 FILLER_16_1133 ();
 sg13g2_decap_8 FILLER_16_1140 ();
 sg13g2_decap_4 FILLER_16_1147 ();
 sg13g2_fill_2 FILLER_16_1151 ();
 sg13g2_decap_8 FILLER_16_1159 ();
 sg13g2_decap_8 FILLER_16_1166 ();
 sg13g2_decap_8 FILLER_16_1173 ();
 sg13g2_decap_4 FILLER_16_1194 ();
 sg13g2_fill_1 FILLER_16_1198 ();
 sg13g2_fill_2 FILLER_16_1211 ();
 sg13g2_fill_2 FILLER_16_1217 ();
 sg13g2_fill_2 FILLER_16_1224 ();
 sg13g2_decap_8 FILLER_16_1244 ();
 sg13g2_decap_8 FILLER_16_1251 ();
 sg13g2_decap_4 FILLER_16_1258 ();
 sg13g2_decap_8 FILLER_16_1268 ();
 sg13g2_decap_8 FILLER_16_1275 ();
 sg13g2_fill_2 FILLER_16_1282 ();
 sg13g2_decap_8 FILLER_16_1441 ();
 sg13g2_fill_1 FILLER_16_1448 ();
 sg13g2_fill_2 FILLER_16_1471 ();
 sg13g2_fill_1 FILLER_16_1473 ();
 sg13g2_fill_2 FILLER_16_1483 ();
 sg13g2_fill_2 FILLER_16_1495 ();
 sg13g2_fill_1 FILLER_16_1497 ();
 sg13g2_fill_1 FILLER_16_1553 ();
 sg13g2_fill_1 FILLER_16_1626 ();
 sg13g2_fill_2 FILLER_16_1681 ();
 sg13g2_fill_1 FILLER_16_1683 ();
 sg13g2_fill_2 FILLER_16_1756 ();
 sg13g2_fill_1 FILLER_16_1758 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_59 ();
 sg13g2_decap_8 FILLER_17_73 ();
 sg13g2_decap_8 FILLER_17_80 ();
 sg13g2_decap_8 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_fill_1 FILLER_17_96 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_4 FILLER_17_129 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_176 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_222 ();
 sg13g2_fill_2 FILLER_17_238 ();
 sg13g2_fill_1 FILLER_17_240 ();
 sg13g2_decap_8 FILLER_17_255 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_297 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_decap_8 FILLER_17_313 ();
 sg13g2_fill_2 FILLER_17_320 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_fill_2 FILLER_17_354 ();
 sg13g2_fill_1 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_fill_2 FILLER_17_368 ();
 sg13g2_decap_4 FILLER_17_391 ();
 sg13g2_fill_1 FILLER_17_400 ();
 sg13g2_fill_1 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_17_416 ();
 sg13g2_decap_8 FILLER_17_423 ();
 sg13g2_fill_2 FILLER_17_430 ();
 sg13g2_fill_1 FILLER_17_432 ();
 sg13g2_decap_8 FILLER_17_447 ();
 sg13g2_decap_8 FILLER_17_454 ();
 sg13g2_fill_2 FILLER_17_461 ();
 sg13g2_decap_4 FILLER_17_467 ();
 sg13g2_fill_1 FILLER_17_471 ();
 sg13g2_decap_8 FILLER_17_481 ();
 sg13g2_fill_2 FILLER_17_488 ();
 sg13g2_decap_8 FILLER_17_527 ();
 sg13g2_fill_2 FILLER_17_534 ();
 sg13g2_fill_1 FILLER_17_536 ();
 sg13g2_fill_1 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_551 ();
 sg13g2_decap_8 FILLER_17_558 ();
 sg13g2_fill_2 FILLER_17_565 ();
 sg13g2_fill_1 FILLER_17_571 ();
 sg13g2_decap_8 FILLER_17_578 ();
 sg13g2_fill_1 FILLER_17_585 ();
 sg13g2_decap_4 FILLER_17_603 ();
 sg13g2_fill_1 FILLER_17_624 ();
 sg13g2_fill_2 FILLER_17_629 ();
 sg13g2_decap_8 FILLER_17_640 ();
 sg13g2_decap_4 FILLER_17_647 ();
 sg13g2_fill_2 FILLER_17_655 ();
 sg13g2_fill_1 FILLER_17_657 ();
 sg13g2_fill_2 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_678 ();
 sg13g2_fill_2 FILLER_17_685 ();
 sg13g2_fill_2 FILLER_17_717 ();
 sg13g2_decap_4 FILLER_17_728 ();
 sg13g2_fill_1 FILLER_17_732 ();
 sg13g2_decap_4 FILLER_17_743 ();
 sg13g2_decap_8 FILLER_17_766 ();
 sg13g2_decap_8 FILLER_17_773 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_fill_2 FILLER_17_798 ();
 sg13g2_fill_1 FILLER_17_800 ();
 sg13g2_decap_4 FILLER_17_807 ();
 sg13g2_fill_1 FILLER_17_811 ();
 sg13g2_fill_1 FILLER_17_821 ();
 sg13g2_fill_2 FILLER_17_827 ();
 sg13g2_fill_1 FILLER_17_829 ();
 sg13g2_fill_2 FILLER_17_836 ();
 sg13g2_decap_4 FILLER_17_851 ();
 sg13g2_fill_1 FILLER_17_855 ();
 sg13g2_fill_2 FILLER_17_876 ();
 sg13g2_fill_2 FILLER_17_897 ();
 sg13g2_decap_8 FILLER_17_954 ();
 sg13g2_fill_2 FILLER_17_961 ();
 sg13g2_decap_8 FILLER_17_967 ();
 sg13g2_fill_2 FILLER_17_974 ();
 sg13g2_fill_1 FILLER_17_976 ();
 sg13g2_fill_2 FILLER_17_1000 ();
 sg13g2_fill_2 FILLER_17_1026 ();
 sg13g2_decap_8 FILLER_17_1032 ();
 sg13g2_decap_4 FILLER_17_1039 ();
 sg13g2_fill_2 FILLER_17_1043 ();
 sg13g2_fill_1 FILLER_17_1072 ();
 sg13g2_decap_8 FILLER_17_1085 ();
 sg13g2_decap_8 FILLER_17_1092 ();
 sg13g2_decap_4 FILLER_17_1099 ();
 sg13g2_fill_1 FILLER_17_1124 ();
 sg13g2_decap_4 FILLER_17_1143 ();
 sg13g2_fill_2 FILLER_17_1147 ();
 sg13g2_decap_8 FILLER_17_1155 ();
 sg13g2_fill_2 FILLER_17_1162 ();
 sg13g2_fill_1 FILLER_17_1164 ();
 sg13g2_decap_4 FILLER_17_1173 ();
 sg13g2_fill_2 FILLER_17_1177 ();
 sg13g2_decap_8 FILLER_17_1191 ();
 sg13g2_fill_2 FILLER_17_1198 ();
 sg13g2_decap_8 FILLER_17_1206 ();
 sg13g2_decap_8 FILLER_17_1213 ();
 sg13g2_decap_8 FILLER_17_1220 ();
 sg13g2_decap_4 FILLER_17_1227 ();
 sg13g2_fill_1 FILLER_17_1231 ();
 sg13g2_decap_4 FILLER_17_1237 ();
 sg13g2_fill_2 FILLER_17_1241 ();
 sg13g2_decap_8 FILLER_17_1249 ();
 sg13g2_decap_8 FILLER_17_1256 ();
 sg13g2_fill_1 FILLER_17_1263 ();
 sg13g2_decap_8 FILLER_17_1270 ();
 sg13g2_decap_8 FILLER_17_1277 ();
 sg13g2_decap_4 FILLER_17_1284 ();
 sg13g2_fill_1 FILLER_17_1288 ();
 sg13g2_fill_2 FILLER_17_1339 ();
 sg13g2_fill_1 FILLER_17_1341 ();
 sg13g2_fill_2 FILLER_17_1346 ();
 sg13g2_fill_1 FILLER_17_1367 ();
 sg13g2_fill_2 FILLER_17_1402 ();
 sg13g2_fill_1 FILLER_17_1404 ();
 sg13g2_fill_2 FILLER_17_1435 ();
 sg13g2_decap_8 FILLER_17_1441 ();
 sg13g2_decap_4 FILLER_17_1448 ();
 sg13g2_fill_1 FILLER_17_1452 ();
 sg13g2_fill_1 FILLER_17_1498 ();
 sg13g2_decap_8 FILLER_17_1508 ();
 sg13g2_decap_8 FILLER_17_1515 ();
 sg13g2_decap_4 FILLER_17_1522 ();
 sg13g2_fill_1 FILLER_17_1526 ();
 sg13g2_decap_8 FILLER_17_1544 ();
 sg13g2_decap_8 FILLER_17_1551 ();
 sg13g2_fill_1 FILLER_17_1558 ();
 sg13g2_decap_8 FILLER_17_1563 ();
 sg13g2_decap_8 FILLER_17_1570 ();
 sg13g2_fill_2 FILLER_17_1577 ();
 sg13g2_fill_2 FILLER_17_1583 ();
 sg13g2_fill_2 FILLER_17_1651 ();
 sg13g2_fill_2 FILLER_17_1675 ();
 sg13g2_fill_1 FILLER_17_1677 ();
 sg13g2_fill_1 FILLER_17_1714 ();
 sg13g2_fill_2 FILLER_17_1724 ();
 sg13g2_fill_1 FILLER_17_1726 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_30 ();
 sg13g2_fill_1 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_72 ();
 sg13g2_decap_4 FILLER_18_101 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_4 FILLER_18_175 ();
 sg13g2_fill_1 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_197 ();
 sg13g2_decap_8 FILLER_18_204 ();
 sg13g2_decap_4 FILLER_18_211 ();
 sg13g2_fill_2 FILLER_18_215 ();
 sg13g2_decap_4 FILLER_18_222 ();
 sg13g2_fill_2 FILLER_18_226 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_2 FILLER_18_248 ();
 sg13g2_decap_8 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_261 ();
 sg13g2_decap_4 FILLER_18_289 ();
 sg13g2_fill_1 FILLER_18_293 ();
 sg13g2_decap_8 FILLER_18_304 ();
 sg13g2_decap_8 FILLER_18_311 ();
 sg13g2_fill_2 FILLER_18_318 ();
 sg13g2_fill_1 FILLER_18_320 ();
 sg13g2_fill_2 FILLER_18_325 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_decap_4 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_365 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_fill_2 FILLER_18_379 ();
 sg13g2_fill_1 FILLER_18_381 ();
 sg13g2_fill_2 FILLER_18_385 ();
 sg13g2_fill_2 FILLER_18_392 ();
 sg13g2_fill_1 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_409 ();
 sg13g2_fill_1 FILLER_18_416 ();
 sg13g2_decap_8 FILLER_18_432 ();
 sg13g2_decap_8 FILLER_18_439 ();
 sg13g2_decap_4 FILLER_18_446 ();
 sg13g2_fill_2 FILLER_18_450 ();
 sg13g2_decap_4 FILLER_18_465 ();
 sg13g2_fill_2 FILLER_18_469 ();
 sg13g2_decap_4 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_542 ();
 sg13g2_fill_2 FILLER_18_549 ();
 sg13g2_fill_1 FILLER_18_551 ();
 sg13g2_fill_1 FILLER_18_580 ();
 sg13g2_fill_2 FILLER_18_586 ();
 sg13g2_fill_1 FILLER_18_588 ();
 sg13g2_fill_1 FILLER_18_616 ();
 sg13g2_fill_2 FILLER_18_651 ();
 sg13g2_fill_1 FILLER_18_721 ();
 sg13g2_fill_1 FILLER_18_738 ();
 sg13g2_fill_2 FILLER_18_752 ();
 sg13g2_decap_4 FILLER_18_758 ();
 sg13g2_fill_1 FILLER_18_784 ();
 sg13g2_fill_2 FILLER_18_799 ();
 sg13g2_decap_8 FILLER_18_806 ();
 sg13g2_decap_8 FILLER_18_813 ();
 sg13g2_fill_2 FILLER_18_820 ();
 sg13g2_fill_1 FILLER_18_822 ();
 sg13g2_decap_8 FILLER_18_832 ();
 sg13g2_fill_1 FILLER_18_839 ();
 sg13g2_decap_4 FILLER_18_850 ();
 sg13g2_fill_1 FILLER_18_863 ();
 sg13g2_fill_2 FILLER_18_870 ();
 sg13g2_decap_4 FILLER_18_882 ();
 sg13g2_fill_1 FILLER_18_886 ();
 sg13g2_decap_8 FILLER_18_913 ();
 sg13g2_fill_2 FILLER_18_920 ();
 sg13g2_fill_2 FILLER_18_935 ();
 sg13g2_fill_1 FILLER_18_937 ();
 sg13g2_fill_2 FILLER_18_956 ();
 sg13g2_fill_1 FILLER_18_999 ();
 sg13g2_decap_4 FILLER_18_1019 ();
 sg13g2_fill_1 FILLER_18_1051 ();
 sg13g2_decap_4 FILLER_18_1081 ();
 sg13g2_fill_2 FILLER_18_1085 ();
 sg13g2_fill_2 FILLER_18_1092 ();
 sg13g2_fill_1 FILLER_18_1094 ();
 sg13g2_decap_4 FILLER_18_1121 ();
 sg13g2_fill_2 FILLER_18_1143 ();
 sg13g2_decap_8 FILLER_18_1163 ();
 sg13g2_decap_8 FILLER_18_1170 ();
 sg13g2_decap_4 FILLER_18_1177 ();
 sg13g2_fill_2 FILLER_18_1181 ();
 sg13g2_decap_4 FILLER_18_1189 ();
 sg13g2_decap_8 FILLER_18_1217 ();
 sg13g2_decap_8 FILLER_18_1224 ();
 sg13g2_decap_4 FILLER_18_1231 ();
 sg13g2_fill_2 FILLER_18_1235 ();
 sg13g2_decap_8 FILLER_18_1243 ();
 sg13g2_decap_8 FILLER_18_1250 ();
 sg13g2_decap_8 FILLER_18_1263 ();
 sg13g2_decap_8 FILLER_18_1270 ();
 sg13g2_decap_4 FILLER_18_1277 ();
 sg13g2_fill_2 FILLER_18_1281 ();
 sg13g2_decap_8 FILLER_18_1311 ();
 sg13g2_decap_8 FILLER_18_1318 ();
 sg13g2_decap_8 FILLER_18_1325 ();
 sg13g2_decap_4 FILLER_18_1332 ();
 sg13g2_fill_1 FILLER_18_1336 ();
 sg13g2_fill_2 FILLER_18_1369 ();
 sg13g2_fill_2 FILLER_18_1420 ();
 sg13g2_fill_1 FILLER_18_1422 ();
 sg13g2_fill_2 FILLER_18_1477 ();
 sg13g2_fill_1 FILLER_18_1479 ();
 sg13g2_decap_8 FILLER_18_1543 ();
 sg13g2_fill_2 FILLER_18_1563 ();
 sg13g2_fill_1 FILLER_18_1565 ();
 sg13g2_fill_1 FILLER_18_1602 ();
 sg13g2_decap_4 FILLER_18_1702 ();
 sg13g2_decap_4 FILLER_18_1764 ();
 sg13g2_fill_1 FILLER_19_28 ();
 sg13g2_fill_2 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_decap_4 FILLER_19_103 ();
 sg13g2_decap_8 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_8 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_132 ();
 sg13g2_fill_2 FILLER_19_148 ();
 sg13g2_fill_1 FILLER_19_150 ();
 sg13g2_fill_2 FILLER_19_159 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_4 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_204 ();
 sg13g2_decap_4 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_271 ();
 sg13g2_decap_4 FILLER_19_312 ();
 sg13g2_fill_2 FILLER_19_335 ();
 sg13g2_fill_2 FILLER_19_355 ();
 sg13g2_fill_1 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_373 ();
 sg13g2_fill_2 FILLER_19_380 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_fill_2 FILLER_19_417 ();
 sg13g2_fill_1 FILLER_19_419 ();
 sg13g2_decap_8 FILLER_19_433 ();
 sg13g2_decap_8 FILLER_19_440 ();
 sg13g2_decap_4 FILLER_19_447 ();
 sg13g2_decap_4 FILLER_19_461 ();
 sg13g2_fill_1 FILLER_19_465 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_4 FILLER_19_490 ();
 sg13g2_fill_2 FILLER_19_494 ();
 sg13g2_fill_2 FILLER_19_508 ();
 sg13g2_fill_1 FILLER_19_510 ();
 sg13g2_decap_8 FILLER_19_535 ();
 sg13g2_fill_1 FILLER_19_545 ();
 sg13g2_decap_8 FILLER_19_572 ();
 sg13g2_decap_8 FILLER_19_579 ();
 sg13g2_decap_8 FILLER_19_586 ();
 sg13g2_fill_2 FILLER_19_593 ();
 sg13g2_fill_2 FILLER_19_638 ();
 sg13g2_fill_2 FILLER_19_654 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_fill_2 FILLER_19_676 ();
 sg13g2_fill_2 FILLER_19_683 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_fill_2 FILLER_19_697 ();
 sg13g2_fill_1 FILLER_19_699 ();
 sg13g2_fill_1 FILLER_19_705 ();
 sg13g2_decap_8 FILLER_19_712 ();
 sg13g2_decap_4 FILLER_19_719 ();
 sg13g2_fill_1 FILLER_19_743 ();
 sg13g2_decap_8 FILLER_19_752 ();
 sg13g2_decap_8 FILLER_19_759 ();
 sg13g2_decap_8 FILLER_19_766 ();
 sg13g2_fill_1 FILLER_19_773 ();
 sg13g2_fill_1 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_fill_1 FILLER_19_827 ();
 sg13g2_fill_2 FILLER_19_850 ();
 sg13g2_fill_1 FILLER_19_858 ();
 sg13g2_decap_8 FILLER_19_872 ();
 sg13g2_decap_8 FILLER_19_879 ();
 sg13g2_decap_4 FILLER_19_886 ();
 sg13g2_fill_2 FILLER_19_890 ();
 sg13g2_fill_1 FILLER_19_913 ();
 sg13g2_fill_2 FILLER_19_930 ();
 sg13g2_fill_2 FILLER_19_945 ();
 sg13g2_fill_1 FILLER_19_947 ();
 sg13g2_fill_2 FILLER_19_958 ();
 sg13g2_fill_2 FILLER_19_987 ();
 sg13g2_fill_1 FILLER_19_989 ();
 sg13g2_fill_2 FILLER_19_999 ();
 sg13g2_fill_2 FILLER_19_1025 ();
 sg13g2_decap_8 FILLER_19_1031 ();
 sg13g2_fill_2 FILLER_19_1042 ();
 sg13g2_fill_1 FILLER_19_1044 ();
 sg13g2_decap_8 FILLER_19_1075 ();
 sg13g2_fill_1 FILLER_19_1097 ();
 sg13g2_decap_8 FILLER_19_1106 ();
 sg13g2_fill_1 FILLER_19_1113 ();
 sg13g2_decap_4 FILLER_19_1122 ();
 sg13g2_fill_1 FILLER_19_1126 ();
 sg13g2_decap_8 FILLER_19_1133 ();
 sg13g2_decap_8 FILLER_19_1140 ();
 sg13g2_decap_8 FILLER_19_1147 ();
 sg13g2_decap_8 FILLER_19_1154 ();
 sg13g2_decap_8 FILLER_19_1161 ();
 sg13g2_decap_8 FILLER_19_1168 ();
 sg13g2_decap_4 FILLER_19_1175 ();
 sg13g2_fill_2 FILLER_19_1179 ();
 sg13g2_fill_2 FILLER_19_1193 ();
 sg13g2_fill_1 FILLER_19_1195 ();
 sg13g2_fill_2 FILLER_19_1208 ();
 sg13g2_fill_2 FILLER_19_1216 ();
 sg13g2_fill_1 FILLER_19_1218 ();
 sg13g2_fill_2 FILLER_19_1224 ();
 sg13g2_decap_8 FILLER_19_1238 ();
 sg13g2_decap_8 FILLER_19_1245 ();
 sg13g2_decap_8 FILLER_19_1252 ();
 sg13g2_decap_4 FILLER_19_1269 ();
 sg13g2_fill_1 FILLER_19_1273 ();
 sg13g2_decap_8 FILLER_19_1292 ();
 sg13g2_fill_2 FILLER_19_1299 ();
 sg13g2_fill_1 FILLER_19_1301 ();
 sg13g2_decap_4 FILLER_19_1312 ();
 sg13g2_fill_1 FILLER_19_1316 ();
 sg13g2_decap_4 FILLER_19_1321 ();
 sg13g2_fill_1 FILLER_19_1325 ();
 sg13g2_fill_2 FILLER_19_1393 ();
 sg13g2_decap_4 FILLER_19_1463 ();
 sg13g2_fill_2 FILLER_19_1471 ();
 sg13g2_fill_2 FILLER_19_1496 ();
 sg13g2_fill_2 FILLER_19_1520 ();
 sg13g2_fill_1 FILLER_19_1522 ();
 sg13g2_fill_1 FILLER_19_1594 ();
 sg13g2_fill_2 FILLER_19_1604 ();
 sg13g2_fill_2 FILLER_19_1619 ();
 sg13g2_fill_2 FILLER_19_1634 ();
 sg13g2_decap_4 FILLER_19_1645 ();
 sg13g2_fill_1 FILLER_19_1649 ();
 sg13g2_decap_8 FILLER_19_1667 ();
 sg13g2_fill_2 FILLER_19_1674 ();
 sg13g2_fill_1 FILLER_19_1676 ();
 sg13g2_decap_4 FILLER_19_1694 ();
 sg13g2_fill_2 FILLER_19_1698 ();
 sg13g2_fill_2 FILLER_19_1713 ();
 sg13g2_fill_2 FILLER_19_1719 ();
 sg13g2_fill_2 FILLER_19_1766 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_34 ();
 sg13g2_decap_8 FILLER_20_51 ();
 sg13g2_decap_4 FILLER_20_58 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_fill_2 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_fill_1 FILLER_20_118 ();
 sg13g2_fill_2 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_139 ();
 sg13g2_decap_4 FILLER_20_145 ();
 sg13g2_fill_2 FILLER_20_149 ();
 sg13g2_fill_1 FILLER_20_171 ();
 sg13g2_fill_2 FILLER_20_187 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_fill_1 FILLER_20_200 ();
 sg13g2_decap_4 FILLER_20_209 ();
 sg13g2_decap_8 FILLER_20_226 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_4 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_decap_8 FILLER_20_300 ();
 sg13g2_decap_4 FILLER_20_307 ();
 sg13g2_fill_2 FILLER_20_311 ();
 sg13g2_fill_2 FILLER_20_329 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_20_381 ();
 sg13g2_fill_1 FILLER_20_383 ();
 sg13g2_fill_2 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_401 ();
 sg13g2_decap_8 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_20_415 ();
 sg13g2_fill_1 FILLER_20_422 ();
 sg13g2_fill_2 FILLER_20_446 ();
 sg13g2_fill_1 FILLER_20_448 ();
 sg13g2_decap_8 FILLER_20_459 ();
 sg13g2_decap_8 FILLER_20_477 ();
 sg13g2_fill_2 FILLER_20_484 ();
 sg13g2_fill_1 FILLER_20_486 ();
 sg13g2_fill_2 FILLER_20_524 ();
 sg13g2_fill_2 FILLER_20_609 ();
 sg13g2_fill_1 FILLER_20_611 ();
 sg13g2_fill_1 FILLER_20_640 ();
 sg13g2_decap_8 FILLER_20_695 ();
 sg13g2_decap_8 FILLER_20_702 ();
 sg13g2_fill_2 FILLER_20_709 ();
 sg13g2_fill_1 FILLER_20_711 ();
 sg13g2_decap_8 FILLER_20_719 ();
 sg13g2_fill_2 FILLER_20_726 ();
 sg13g2_fill_2 FILLER_20_753 ();
 sg13g2_decap_4 FILLER_20_774 ();
 sg13g2_fill_2 FILLER_20_797 ();
 sg13g2_decap_4 FILLER_20_805 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_fill_1 FILLER_20_841 ();
 sg13g2_decap_8 FILLER_20_846 ();
 sg13g2_fill_2 FILLER_20_853 ();
 sg13g2_fill_1 FILLER_20_855 ();
 sg13g2_decap_8 FILLER_20_860 ();
 sg13g2_fill_1 FILLER_20_867 ();
 sg13g2_decap_4 FILLER_20_873 ();
 sg13g2_fill_2 FILLER_20_895 ();
 sg13g2_fill_1 FILLER_20_897 ();
 sg13g2_decap_4 FILLER_20_909 ();
 sg13g2_fill_2 FILLER_20_913 ();
 sg13g2_decap_8 FILLER_20_918 ();
 sg13g2_decap_8 FILLER_20_925 ();
 sg13g2_fill_1 FILLER_20_932 ();
 sg13g2_decap_4 FILLER_20_965 ();
 sg13g2_fill_1 FILLER_20_969 ();
 sg13g2_fill_1 FILLER_20_998 ();
 sg13g2_fill_2 FILLER_20_1008 ();
 sg13g2_fill_1 FILLER_20_1010 ();
 sg13g2_fill_2 FILLER_20_1024 ();
 sg13g2_fill_1 FILLER_20_1031 ();
 sg13g2_decap_8 FILLER_20_1100 ();
 sg13g2_fill_2 FILLER_20_1107 ();
 sg13g2_fill_1 FILLER_20_1109 ();
 sg13g2_decap_4 FILLER_20_1127 ();
 sg13g2_fill_2 FILLER_20_1131 ();
 sg13g2_decap_8 FILLER_20_1139 ();
 sg13g2_decap_4 FILLER_20_1146 ();
 sg13g2_fill_2 FILLER_20_1150 ();
 sg13g2_decap_8 FILLER_20_1158 ();
 sg13g2_decap_8 FILLER_20_1165 ();
 sg13g2_decap_8 FILLER_20_1172 ();
 sg13g2_fill_2 FILLER_20_1179 ();
 sg13g2_decap_4 FILLER_20_1194 ();
 sg13g2_fill_1 FILLER_20_1198 ();
 sg13g2_decap_8 FILLER_20_1226 ();
 sg13g2_decap_8 FILLER_20_1233 ();
 sg13g2_decap_8 FILLER_20_1240 ();
 sg13g2_decap_4 FILLER_20_1247 ();
 sg13g2_decap_4 FILLER_20_1279 ();
 sg13g2_fill_2 FILLER_20_1311 ();
 sg13g2_fill_2 FILLER_20_1353 ();
 sg13g2_fill_1 FILLER_20_1355 ();
 sg13g2_fill_1 FILLER_20_1391 ();
 sg13g2_decap_8 FILLER_20_1454 ();
 sg13g2_decap_4 FILLER_20_1499 ();
 sg13g2_decap_4 FILLER_20_1588 ();
 sg13g2_decap_4 FILLER_20_1619 ();
 sg13g2_fill_1 FILLER_20_1740 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_54 ();
 sg13g2_fill_1 FILLER_21_56 ();
 sg13g2_fill_2 FILLER_21_77 ();
 sg13g2_fill_1 FILLER_21_79 ();
 sg13g2_decap_8 FILLER_21_107 ();
 sg13g2_decap_8 FILLER_21_114 ();
 sg13g2_fill_2 FILLER_21_121 ();
 sg13g2_decap_8 FILLER_21_141 ();
 sg13g2_decap_4 FILLER_21_148 ();
 sg13g2_fill_1 FILLER_21_155 ();
 sg13g2_decap_8 FILLER_21_169 ();
 sg13g2_decap_4 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_185 ();
 sg13g2_fill_2 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_239 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_2 FILLER_21_265 ();
 sg13g2_decap_4 FILLER_21_271 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_310 ();
 sg13g2_fill_2 FILLER_21_320 ();
 sg13g2_decap_8 FILLER_21_330 ();
 sg13g2_fill_1 FILLER_21_337 ();
 sg13g2_fill_2 FILLER_21_348 ();
 sg13g2_fill_1 FILLER_21_350 ();
 sg13g2_fill_2 FILLER_21_355 ();
 sg13g2_fill_1 FILLER_21_357 ();
 sg13g2_decap_4 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_decap_8 FILLER_21_411 ();
 sg13g2_decap_8 FILLER_21_436 ();
 sg13g2_fill_1 FILLER_21_454 ();
 sg13g2_fill_1 FILLER_21_460 ();
 sg13g2_fill_2 FILLER_21_469 ();
 sg13g2_fill_1 FILLER_21_471 ();
 sg13g2_decap_8 FILLER_21_487 ();
 sg13g2_decap_8 FILLER_21_505 ();
 sg13g2_decap_4 FILLER_21_512 ();
 sg13g2_fill_1 FILLER_21_548 ();
 sg13g2_decap_4 FILLER_21_559 ();
 sg13g2_fill_1 FILLER_21_563 ();
 sg13g2_fill_2 FILLER_21_570 ();
 sg13g2_fill_2 FILLER_21_590 ();
 sg13g2_fill_1 FILLER_21_592 ();
 sg13g2_fill_2 FILLER_21_609 ();
 sg13g2_fill_1 FILLER_21_611 ();
 sg13g2_decap_4 FILLER_21_624 ();
 sg13g2_decap_8 FILLER_21_632 ();
 sg13g2_fill_2 FILLER_21_639 ();
 sg13g2_fill_1 FILLER_21_641 ();
 sg13g2_fill_2 FILLER_21_674 ();
 sg13g2_fill_1 FILLER_21_676 ();
 sg13g2_decap_4 FILLER_21_714 ();
 sg13g2_fill_2 FILLER_21_718 ();
 sg13g2_fill_2 FILLER_21_742 ();
 sg13g2_fill_1 FILLER_21_744 ();
 sg13g2_decap_8 FILLER_21_759 ();
 sg13g2_decap_4 FILLER_21_766 ();
 sg13g2_fill_2 FILLER_21_770 ();
 sg13g2_fill_1 FILLER_21_777 ();
 sg13g2_decap_4 FILLER_21_800 ();
 sg13g2_fill_2 FILLER_21_804 ();
 sg13g2_fill_2 FILLER_21_811 ();
 sg13g2_fill_1 FILLER_21_813 ();
 sg13g2_fill_2 FILLER_21_823 ();
 sg13g2_fill_1 FILLER_21_825 ();
 sg13g2_decap_4 FILLER_21_835 ();
 sg13g2_decap_8 FILLER_21_855 ();
 sg13g2_decap_4 FILLER_21_862 ();
 sg13g2_decap_4 FILLER_21_877 ();
 sg13g2_fill_1 FILLER_21_894 ();
 sg13g2_decap_4 FILLER_21_900 ();
 sg13g2_fill_1 FILLER_21_904 ();
 sg13g2_decap_8 FILLER_21_914 ();
 sg13g2_decap_8 FILLER_21_921 ();
 sg13g2_fill_2 FILLER_21_942 ();
 sg13g2_decap_4 FILLER_21_962 ();
 sg13g2_fill_1 FILLER_21_966 ();
 sg13g2_fill_2 FILLER_21_971 ();
 sg13g2_fill_1 FILLER_21_973 ();
 sg13g2_fill_2 FILLER_21_1013 ();
 sg13g2_fill_2 FILLER_21_1028 ();
 sg13g2_decap_8 FILLER_21_1035 ();
 sg13g2_decap_8 FILLER_21_1042 ();
 sg13g2_fill_2 FILLER_21_1049 ();
 sg13g2_fill_1 FILLER_21_1051 ();
 sg13g2_decap_8 FILLER_21_1078 ();
 sg13g2_fill_2 FILLER_21_1085 ();
 sg13g2_fill_2 FILLER_21_1092 ();
 sg13g2_fill_1 FILLER_21_1094 ();
 sg13g2_decap_8 FILLER_21_1099 ();
 sg13g2_decap_8 FILLER_21_1124 ();
 sg13g2_decap_8 FILLER_21_1131 ();
 sg13g2_decap_8 FILLER_21_1138 ();
 sg13g2_decap_8 FILLER_21_1145 ();
 sg13g2_fill_1 FILLER_21_1152 ();
 sg13g2_fill_1 FILLER_21_1166 ();
 sg13g2_fill_2 FILLER_21_1184 ();
 sg13g2_decap_4 FILLER_21_1195 ();
 sg13g2_fill_2 FILLER_21_1221 ();
 sg13g2_fill_1 FILLER_21_1223 ();
 sg13g2_decap_8 FILLER_21_1230 ();
 sg13g2_decap_8 FILLER_21_1237 ();
 sg13g2_fill_1 FILLER_21_1257 ();
 sg13g2_fill_1 FILLER_21_1262 ();
 sg13g2_decap_4 FILLER_21_1291 ();
 sg13g2_fill_1 FILLER_21_1295 ();
 sg13g2_decap_8 FILLER_21_1309 ();
 sg13g2_fill_1 FILLER_21_1316 ();
 sg13g2_decap_8 FILLER_21_1330 ();
 sg13g2_fill_2 FILLER_21_1337 ();
 sg13g2_fill_1 FILLER_21_1339 ();
 sg13g2_fill_2 FILLER_21_1403 ();
 sg13g2_decap_8 FILLER_21_1446 ();
 sg13g2_fill_2 FILLER_21_1453 ();
 sg13g2_decap_8 FILLER_21_1519 ();
 sg13g2_fill_2 FILLER_21_1526 ();
 sg13g2_fill_1 FILLER_21_1528 ();
 sg13g2_decap_4 FILLER_21_1533 ();
 sg13g2_decap_8 FILLER_21_1541 ();
 sg13g2_fill_2 FILLER_21_1548 ();
 sg13g2_fill_1 FILLER_21_1550 ();
 sg13g2_decap_4 FILLER_21_1645 ();
 sg13g2_fill_1 FILLER_21_1649 ();
 sg13g2_decap_8 FILLER_21_1663 ();
 sg13g2_decap_4 FILLER_21_1670 ();
 sg13g2_fill_1 FILLER_21_1674 ();
 sg13g2_decap_8 FILLER_21_1715 ();
 sg13g2_decap_4 FILLER_21_1722 ();
 sg13g2_decap_8 FILLER_21_1730 ();
 sg13g2_decap_8 FILLER_21_1737 ();
 sg13g2_fill_2 FILLER_21_1744 ();
 sg13g2_decap_8 FILLER_21_1754 ();
 sg13g2_decap_8 FILLER_21_1761 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_4 ();
 sg13g2_fill_1 FILLER_22_33 ();
 sg13g2_decap_4 FILLER_22_44 ();
 sg13g2_fill_1 FILLER_22_48 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_decap_4 FILLER_22_78 ();
 sg13g2_decap_8 FILLER_22_120 ();
 sg13g2_fill_1 FILLER_22_127 ();
 sg13g2_decap_4 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_fill_2 FILLER_22_185 ();
 sg13g2_decap_8 FILLER_22_205 ();
 sg13g2_fill_2 FILLER_22_212 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_8 FILLER_22_234 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_287 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_decap_8 FILLER_22_311 ();
 sg13g2_fill_1 FILLER_22_318 ();
 sg13g2_fill_2 FILLER_22_343 ();
 sg13g2_fill_1 FILLER_22_345 ();
 sg13g2_decap_4 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_387 ();
 sg13g2_decap_4 FILLER_22_417 ();
 sg13g2_fill_1 FILLER_22_421 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_1 FILLER_22_436 ();
 sg13g2_decap_8 FILLER_22_441 ();
 sg13g2_decap_8 FILLER_22_448 ();
 sg13g2_fill_2 FILLER_22_455 ();
 sg13g2_fill_1 FILLER_22_457 ();
 sg13g2_fill_2 FILLER_22_462 ();
 sg13g2_decap_4 FILLER_22_486 ();
 sg13g2_decap_8 FILLER_22_514 ();
 sg13g2_decap_4 FILLER_22_521 ();
 sg13g2_decap_4 FILLER_22_530 ();
 sg13g2_fill_2 FILLER_22_534 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_8 FILLER_22_564 ();
 sg13g2_fill_2 FILLER_22_571 ();
 sg13g2_fill_1 FILLER_22_573 ();
 sg13g2_decap_8 FILLER_22_586 ();
 sg13g2_decap_4 FILLER_22_593 ();
 sg13g2_fill_2 FILLER_22_601 ();
 sg13g2_fill_1 FILLER_22_603 ();
 sg13g2_fill_2 FILLER_22_657 ();
 sg13g2_fill_1 FILLER_22_659 ();
 sg13g2_decap_8 FILLER_22_677 ();
 sg13g2_decap_4 FILLER_22_684 ();
 sg13g2_fill_2 FILLER_22_705 ();
 sg13g2_fill_1 FILLER_22_707 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_fill_2 FILLER_22_739 ();
 sg13g2_fill_1 FILLER_22_741 ();
 sg13g2_decap_4 FILLER_22_746 ();
 sg13g2_fill_2 FILLER_22_750 ();
 sg13g2_fill_1 FILLER_22_757 ();
 sg13g2_decap_4 FILLER_22_776 ();
 sg13g2_fill_1 FILLER_22_780 ();
 sg13g2_decap_8 FILLER_22_800 ();
 sg13g2_fill_2 FILLER_22_835 ();
 sg13g2_fill_1 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_fill_1 FILLER_22_858 ();
 sg13g2_fill_1 FILLER_22_864 ();
 sg13g2_decap_4 FILLER_22_900 ();
 sg13g2_fill_2 FILLER_22_916 ();
 sg13g2_fill_1 FILLER_22_918 ();
 sg13g2_decap_8 FILLER_22_989 ();
 sg13g2_decap_4 FILLER_22_996 ();
 sg13g2_decap_8 FILLER_22_1005 ();
 sg13g2_fill_2 FILLER_22_1012 ();
 sg13g2_fill_1 FILLER_22_1014 ();
 sg13g2_decap_8 FILLER_22_1020 ();
 sg13g2_decap_4 FILLER_22_1027 ();
 sg13g2_fill_1 FILLER_22_1035 ();
 sg13g2_fill_2 FILLER_22_1064 ();
 sg13g2_fill_2 FILLER_22_1122 ();
 sg13g2_fill_1 FILLER_22_1157 ();
 sg13g2_decap_8 FILLER_22_1171 ();
 sg13g2_decap_8 FILLER_22_1178 ();
 sg13g2_decap_8 FILLER_22_1191 ();
 sg13g2_decap_4 FILLER_22_1204 ();
 sg13g2_fill_1 FILLER_22_1208 ();
 sg13g2_decap_8 FILLER_22_1218 ();
 sg13g2_decap_4 FILLER_22_1225 ();
 sg13g2_fill_2 FILLER_22_1229 ();
 sg13g2_decap_8 FILLER_22_1286 ();
 sg13g2_fill_1 FILLER_22_1293 ();
 sg13g2_fill_2 FILLER_22_1348 ();
 sg13g2_fill_1 FILLER_22_1350 ();
 sg13g2_fill_2 FILLER_22_1364 ();
 sg13g2_fill_2 FILLER_22_1437 ();
 sg13g2_decap_4 FILLER_22_1452 ();
 sg13g2_fill_1 FILLER_22_1456 ();
 sg13g2_decap_8 FILLER_22_1525 ();
 sg13g2_fill_2 FILLER_22_1559 ();
 sg13g2_fill_1 FILLER_22_1561 ();
 sg13g2_fill_2 FILLER_22_1624 ();
 sg13g2_fill_1 FILLER_22_1626 ();
 sg13g2_decap_8 FILLER_22_1694 ();
 sg13g2_decap_8 FILLER_22_1728 ();
 sg13g2_decap_8 FILLER_22_1735 ();
 sg13g2_decap_8 FILLER_22_1742 ();
 sg13g2_decap_8 FILLER_22_1749 ();
 sg13g2_decap_8 FILLER_22_1756 ();
 sg13g2_decap_4 FILLER_22_1763 ();
 sg13g2_fill_1 FILLER_22_1767 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_decap_4 FILLER_23_82 ();
 sg13g2_fill_1 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_97 ();
 sg13g2_fill_2 FILLER_23_136 ();
 sg13g2_fill_1 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_229 ();
 sg13g2_fill_2 FILLER_23_273 ();
 sg13g2_fill_1 FILLER_23_275 ();
 sg13g2_fill_1 FILLER_23_303 ();
 sg13g2_fill_1 FILLER_23_313 ();
 sg13g2_fill_2 FILLER_23_324 ();
 sg13g2_fill_1 FILLER_23_326 ();
 sg13g2_decap_4 FILLER_23_337 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_4 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_384 ();
 sg13g2_fill_2 FILLER_23_391 ();
 sg13g2_fill_1 FILLER_23_393 ();
 sg13g2_decap_4 FILLER_23_398 ();
 sg13g2_fill_1 FILLER_23_402 ();
 sg13g2_decap_4 FILLER_23_435 ();
 sg13g2_fill_1 FILLER_23_439 ();
 sg13g2_fill_1 FILLER_23_498 ();
 sg13g2_decap_4 FILLER_23_515 ();
 sg13g2_fill_2 FILLER_23_531 ();
 sg13g2_decap_8 FILLER_23_554 ();
 sg13g2_decap_8 FILLER_23_561 ();
 sg13g2_fill_2 FILLER_23_568 ();
 sg13g2_fill_1 FILLER_23_570 ();
 sg13g2_decap_4 FILLER_23_580 ();
 sg13g2_fill_2 FILLER_23_620 ();
 sg13g2_fill_1 FILLER_23_622 ();
 sg13g2_fill_2 FILLER_23_645 ();
 sg13g2_decap_8 FILLER_23_692 ();
 sg13g2_decap_8 FILLER_23_699 ();
 sg13g2_decap_4 FILLER_23_706 ();
 sg13g2_fill_2 FILLER_23_710 ();
 sg13g2_decap_4 FILLER_23_718 ();
 sg13g2_fill_1 FILLER_23_744 ();
 sg13g2_decap_4 FILLER_23_758 ();
 sg13g2_fill_2 FILLER_23_780 ();
 sg13g2_fill_1 FILLER_23_782 ();
 sg13g2_decap_4 FILLER_23_799 ();
 sg13g2_fill_2 FILLER_23_813 ();
 sg13g2_fill_1 FILLER_23_815 ();
 sg13g2_decap_4 FILLER_23_829 ();
 sg13g2_fill_1 FILLER_23_838 ();
 sg13g2_decap_4 FILLER_23_856 ();
 sg13g2_fill_2 FILLER_23_860 ();
 sg13g2_decap_8 FILLER_23_877 ();
 sg13g2_fill_2 FILLER_23_884 ();
 sg13g2_fill_1 FILLER_23_886 ();
 sg13g2_decap_8 FILLER_23_900 ();
 sg13g2_fill_2 FILLER_23_907 ();
 sg13g2_fill_1 FILLER_23_909 ();
 sg13g2_decap_8 FILLER_23_916 ();
 sg13g2_fill_1 FILLER_23_923 ();
 sg13g2_fill_1 FILLER_23_930 ();
 sg13g2_fill_2 FILLER_23_954 ();
 sg13g2_fill_1 FILLER_23_956 ();
 sg13g2_fill_1 FILLER_23_1053 ();
 sg13g2_decap_8 FILLER_23_1083 ();
 sg13g2_decap_8 FILLER_23_1090 ();
 sg13g2_decap_8 FILLER_23_1097 ();
 sg13g2_fill_1 FILLER_23_1104 ();
 sg13g2_decap_8 FILLER_23_1142 ();
 sg13g2_fill_2 FILLER_23_1157 ();
 sg13g2_decap_8 FILLER_23_1185 ();
 sg13g2_decap_8 FILLER_23_1192 ();
 sg13g2_decap_4 FILLER_23_1203 ();
 sg13g2_fill_1 FILLER_23_1207 ();
 sg13g2_decap_4 FILLER_23_1218 ();
 sg13g2_fill_1 FILLER_23_1222 ();
 sg13g2_fill_1 FILLER_23_1232 ();
 sg13g2_fill_2 FILLER_23_1250 ();
 sg13g2_fill_1 FILLER_23_1252 ();
 sg13g2_fill_2 FILLER_23_1272 ();
 sg13g2_decap_8 FILLER_23_1314 ();
 sg13g2_decap_4 FILLER_23_1321 ();
 sg13g2_fill_1 FILLER_23_1325 ();
 sg13g2_fill_1 FILLER_23_1330 ();
 sg13g2_fill_1 FILLER_23_1411 ();
 sg13g2_fill_1 FILLER_23_1488 ();
 sg13g2_fill_1 FILLER_23_1516 ();
 sg13g2_decap_8 FILLER_23_1521 ();
 sg13g2_fill_2 FILLER_23_1528 ();
 sg13g2_fill_2 FILLER_23_1632 ();
 sg13g2_decap_8 FILLER_23_1651 ();
 sg13g2_fill_1 FILLER_23_1658 ();
 sg13g2_fill_2 FILLER_23_1717 ();
 sg13g2_fill_1 FILLER_23_1719 ();
 sg13g2_decap_8 FILLER_23_1729 ();
 sg13g2_decap_8 FILLER_23_1736 ();
 sg13g2_decap_8 FILLER_23_1743 ();
 sg13g2_decap_8 FILLER_23_1750 ();
 sg13g2_decap_8 FILLER_23_1757 ();
 sg13g2_decap_4 FILLER_23_1764 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_10 ();
 sg13g2_decap_4 FILLER_24_44 ();
 sg13g2_fill_2 FILLER_24_80 ();
 sg13g2_fill_1 FILLER_24_82 ();
 sg13g2_fill_2 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_decap_8 FILLER_24_184 ();
 sg13g2_decap_8 FILLER_24_191 ();
 sg13g2_decap_8 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_decap_4 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_decap_4 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_309 ();
 sg13g2_decap_4 FILLER_24_316 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_329 ();
 sg13g2_decap_8 FILLER_24_336 ();
 sg13g2_decap_8 FILLER_24_343 ();
 sg13g2_decap_4 FILLER_24_350 ();
 sg13g2_fill_1 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_fill_2 FILLER_24_396 ();
 sg13g2_fill_2 FILLER_24_424 ();
 sg13g2_decap_4 FILLER_24_431 ();
 sg13g2_fill_2 FILLER_24_439 ();
 sg13g2_fill_1 FILLER_24_441 ();
 sg13g2_fill_2 FILLER_24_460 ();
 sg13g2_fill_2 FILLER_24_471 ();
 sg13g2_fill_2 FILLER_24_486 ();
 sg13g2_decap_4 FILLER_24_496 ();
 sg13g2_fill_1 FILLER_24_500 ();
 sg13g2_decap_4 FILLER_24_521 ();
 sg13g2_fill_1 FILLER_24_525 ();
 sg13g2_decap_4 FILLER_24_531 ();
 sg13g2_fill_2 FILLER_24_535 ();
 sg13g2_decap_4 FILLER_24_545 ();
 sg13g2_fill_1 FILLER_24_549 ();
 sg13g2_decap_8 FILLER_24_588 ();
 sg13g2_decap_4 FILLER_24_595 ();
 sg13g2_decap_4 FILLER_24_644 ();
 sg13g2_fill_2 FILLER_24_648 ();
 sg13g2_fill_1 FILLER_24_670 ();
 sg13g2_decap_8 FILLER_24_713 ();
 sg13g2_fill_1 FILLER_24_732 ();
 sg13g2_decap_4 FILLER_24_739 ();
 sg13g2_fill_2 FILLER_24_743 ();
 sg13g2_fill_2 FILLER_24_766 ();
 sg13g2_fill_2 FILLER_24_773 ();
 sg13g2_fill_1 FILLER_24_775 ();
 sg13g2_decap_8 FILLER_24_807 ();
 sg13g2_decap_4 FILLER_24_824 ();
 sg13g2_fill_2 FILLER_24_828 ();
 sg13g2_decap_8 FILLER_24_849 ();
 sg13g2_fill_2 FILLER_24_856 ();
 sg13g2_fill_2 FILLER_24_863 ();
 sg13g2_decap_8 FILLER_24_871 ();
 sg13g2_fill_1 FILLER_24_878 ();
 sg13g2_fill_2 FILLER_24_884 ();
 sg13g2_decap_4 FILLER_24_903 ();
 sg13g2_fill_2 FILLER_24_945 ();
 sg13g2_fill_1 FILLER_24_956 ();
 sg13g2_decap_8 FILLER_24_988 ();
 sg13g2_fill_2 FILLER_24_1003 ();
 sg13g2_fill_1 FILLER_24_1005 ();
 sg13g2_decap_8 FILLER_24_1015 ();
 sg13g2_fill_2 FILLER_24_1022 ();
 sg13g2_fill_1 FILLER_24_1024 ();
 sg13g2_fill_1 FILLER_24_1053 ();
 sg13g2_fill_2 FILLER_24_1064 ();
 sg13g2_fill_1 FILLER_24_1066 ();
 sg13g2_fill_1 FILLER_24_1070 ();
 sg13g2_fill_1 FILLER_24_1084 ();
 sg13g2_fill_2 FILLER_24_1104 ();
 sg13g2_fill_1 FILLER_24_1106 ();
 sg13g2_fill_2 FILLER_24_1140 ();
 sg13g2_fill_1 FILLER_24_1142 ();
 sg13g2_fill_2 FILLER_24_1153 ();
 sg13g2_fill_1 FILLER_24_1193 ();
 sg13g2_decap_4 FILLER_24_1231 ();
 sg13g2_fill_1 FILLER_24_1248 ();
 sg13g2_fill_2 FILLER_24_1277 ();
 sg13g2_decap_8 FILLER_24_1287 ();
 sg13g2_decap_8 FILLER_24_1294 ();
 sg13g2_fill_2 FILLER_24_1328 ();
 sg13g2_decap_8 FILLER_24_1339 ();
 sg13g2_fill_2 FILLER_24_1391 ();
 sg13g2_decap_8 FILLER_24_1406 ();
 sg13g2_fill_1 FILLER_24_1413 ();
 sg13g2_fill_2 FILLER_24_1427 ();
 sg13g2_fill_1 FILLER_24_1429 ();
 sg13g2_decap_4 FILLER_24_1506 ();
 sg13g2_fill_2 FILLER_24_1510 ();
 sg13g2_fill_2 FILLER_24_1575 ();
 sg13g2_fill_1 FILLER_24_1577 ();
 sg13g2_fill_1 FILLER_24_1591 ();
 sg13g2_fill_2 FILLER_24_1605 ();
 sg13g2_decap_4 FILLER_24_1611 ();
 sg13g2_fill_1 FILLER_24_1615 ();
 sg13g2_fill_2 FILLER_24_1679 ();
 sg13g2_fill_1 FILLER_24_1681 ();
 sg13g2_decap_8 FILLER_24_1695 ();
 sg13g2_decap_8 FILLER_24_1702 ();
 sg13g2_decap_8 FILLER_24_1709 ();
 sg13g2_decap_8 FILLER_24_1716 ();
 sg13g2_decap_8 FILLER_24_1723 ();
 sg13g2_decap_8 FILLER_24_1730 ();
 sg13g2_decap_8 FILLER_24_1737 ();
 sg13g2_decap_8 FILLER_24_1744 ();
 sg13g2_decap_8 FILLER_24_1751 ();
 sg13g2_decap_8 FILLER_24_1758 ();
 sg13g2_fill_2 FILLER_24_1765 ();
 sg13g2_fill_1 FILLER_24_1767 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_29 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_fill_2 FILLER_25_83 ();
 sg13g2_fill_1 FILLER_25_85 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_fill_1 FILLER_25_174 ();
 sg13g2_decap_4 FILLER_25_203 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_fill_2 FILLER_25_217 ();
 sg13g2_decap_4 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_269 ();
 sg13g2_decap_8 FILLER_25_276 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_352 ();
 sg13g2_fill_2 FILLER_25_359 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_fill_1 FILLER_25_386 ();
 sg13g2_decap_4 FILLER_25_415 ();
 sg13g2_fill_2 FILLER_25_445 ();
 sg13g2_fill_1 FILLER_25_480 ();
 sg13g2_decap_4 FILLER_25_509 ();
 sg13g2_decap_4 FILLER_25_517 ();
 sg13g2_fill_2 FILLER_25_521 ();
 sg13g2_fill_2 FILLER_25_529 ();
 sg13g2_fill_1 FILLER_25_531 ();
 sg13g2_decap_4 FILLER_25_539 ();
 sg13g2_fill_2 FILLER_25_549 ();
 sg13g2_fill_1 FILLER_25_551 ();
 sg13g2_fill_1 FILLER_25_562 ();
 sg13g2_decap_8 FILLER_25_591 ();
 sg13g2_fill_2 FILLER_25_598 ();
 sg13g2_fill_1 FILLER_25_600 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_fill_2 FILLER_25_644 ();
 sg13g2_fill_2 FILLER_25_697 ();
 sg13g2_decap_4 FILLER_25_717 ();
 sg13g2_fill_1 FILLER_25_721 ();
 sg13g2_fill_2 FILLER_25_731 ();
 sg13g2_fill_1 FILLER_25_733 ();
 sg13g2_fill_1 FILLER_25_739 ();
 sg13g2_decap_8 FILLER_25_745 ();
 sg13g2_fill_2 FILLER_25_752 ();
 sg13g2_fill_1 FILLER_25_759 ();
 sg13g2_fill_2 FILLER_25_765 ();
 sg13g2_fill_2 FILLER_25_776 ();
 sg13g2_decap_8 FILLER_25_786 ();
 sg13g2_decap_8 FILLER_25_793 ();
 sg13g2_decap_8 FILLER_25_800 ();
 sg13g2_decap_4 FILLER_25_807 ();
 sg13g2_fill_1 FILLER_25_811 ();
 sg13g2_decap_4 FILLER_25_818 ();
 sg13g2_fill_2 FILLER_25_828 ();
 sg13g2_decap_8 FILLER_25_848 ();
 sg13g2_decap_8 FILLER_25_896 ();
 sg13g2_fill_2 FILLER_25_903 ();
 sg13g2_fill_1 FILLER_25_905 ();
 sg13g2_fill_2 FILLER_25_925 ();
 sg13g2_fill_1 FILLER_25_1037 ();
 sg13g2_fill_1 FILLER_25_1066 ();
 sg13g2_fill_1 FILLER_25_1126 ();
 sg13g2_decap_4 FILLER_25_1176 ();
 sg13g2_fill_2 FILLER_25_1193 ();
 sg13g2_decap_8 FILLER_25_1222 ();
 sg13g2_fill_2 FILLER_25_1261 ();
 sg13g2_fill_2 FILLER_25_1272 ();
 sg13g2_fill_1 FILLER_25_1274 ();
 sg13g2_fill_2 FILLER_25_1284 ();
 sg13g2_fill_1 FILLER_25_1286 ();
 sg13g2_decap_4 FILLER_25_1300 ();
 sg13g2_fill_1 FILLER_25_1304 ();
 sg13g2_fill_1 FILLER_25_1363 ();
 sg13g2_fill_2 FILLER_25_1445 ();
 sg13g2_fill_1 FILLER_25_1447 ();
 sg13g2_decap_8 FILLER_25_1456 ();
 sg13g2_decap_8 FILLER_25_1463 ();
 sg13g2_decap_4 FILLER_25_1470 ();
 sg13g2_decap_4 FILLER_25_1478 ();
 sg13g2_fill_1 FILLER_25_1482 ();
 sg13g2_decap_8 FILLER_25_1500 ();
 sg13g2_fill_1 FILLER_25_1507 ();
 sg13g2_decap_8 FILLER_25_1523 ();
 sg13g2_decap_8 FILLER_25_1530 ();
 sg13g2_decap_4 FILLER_25_1537 ();
 sg13g2_decap_8 FILLER_25_1555 ();
 sg13g2_decap_4 FILLER_25_1562 ();
 sg13g2_fill_1 FILLER_25_1570 ();
 sg13g2_fill_1 FILLER_25_1575 ();
 sg13g2_decap_4 FILLER_25_1589 ();
 sg13g2_fill_1 FILLER_25_1593 ();
 sg13g2_decap_8 FILLER_25_1604 ();
 sg13g2_decap_4 FILLER_25_1611 ();
 sg13g2_fill_1 FILLER_25_1615 ();
 sg13g2_decap_8 FILLER_25_1629 ();
 sg13g2_fill_2 FILLER_25_1636 ();
 sg13g2_fill_1 FILLER_25_1638 ();
 sg13g2_decap_8 FILLER_25_1655 ();
 sg13g2_decap_8 FILLER_25_1662 ();
 sg13g2_fill_1 FILLER_25_1669 ();
 sg13g2_decap_8 FILLER_25_1674 ();
 sg13g2_decap_8 FILLER_25_1681 ();
 sg13g2_decap_8 FILLER_25_1688 ();
 sg13g2_decap_8 FILLER_25_1695 ();
 sg13g2_decap_8 FILLER_25_1702 ();
 sg13g2_decap_8 FILLER_25_1709 ();
 sg13g2_decap_8 FILLER_25_1716 ();
 sg13g2_decap_8 FILLER_25_1723 ();
 sg13g2_decap_8 FILLER_25_1730 ();
 sg13g2_decap_8 FILLER_25_1737 ();
 sg13g2_decap_8 FILLER_25_1744 ();
 sg13g2_decap_8 FILLER_25_1751 ();
 sg13g2_decap_8 FILLER_25_1758 ();
 sg13g2_fill_2 FILLER_25_1765 ();
 sg13g2_fill_1 FILLER_25_1767 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_4 ();
 sg13g2_decap_4 FILLER_26_35 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_89 ();
 sg13g2_fill_2 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_decap_4 FILLER_26_296 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_334 ();
 sg13g2_decap_4 FILLER_26_341 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_decap_8 FILLER_26_352 ();
 sg13g2_decap_4 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_363 ();
 sg13g2_decap_4 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_404 ();
 sg13g2_fill_2 FILLER_26_426 ();
 sg13g2_decap_4 FILLER_26_436 ();
 sg13g2_fill_1 FILLER_26_440 ();
 sg13g2_fill_1 FILLER_26_482 ();
 sg13g2_decap_8 FILLER_26_519 ();
 sg13g2_fill_2 FILLER_26_526 ();
 sg13g2_fill_1 FILLER_26_528 ();
 sg13g2_fill_1 FILLER_26_557 ();
 sg13g2_fill_1 FILLER_26_567 ();
 sg13g2_fill_2 FILLER_26_578 ();
 sg13g2_decap_4 FILLER_26_590 ();
 sg13g2_fill_2 FILLER_26_594 ();
 sg13g2_fill_2 FILLER_26_609 ();
 sg13g2_fill_1 FILLER_26_611 ();
 sg13g2_fill_2 FILLER_26_624 ();
 sg13g2_fill_2 FILLER_26_635 ();
 sg13g2_fill_2 FILLER_26_654 ();
 sg13g2_fill_2 FILLER_26_693 ();
 sg13g2_decap_4 FILLER_26_713 ();
 sg13g2_fill_2 FILLER_26_717 ();
 sg13g2_decap_4 FILLER_26_741 ();
 sg13g2_fill_1 FILLER_26_745 ();
 sg13g2_fill_2 FILLER_26_750 ();
 sg13g2_fill_2 FILLER_26_767 ();
 sg13g2_fill_1 FILLER_26_769 ();
 sg13g2_fill_2 FILLER_26_788 ();
 sg13g2_fill_1 FILLER_26_790 ();
 sg13g2_fill_2 FILLER_26_806 ();
 sg13g2_fill_1 FILLER_26_814 ();
 sg13g2_fill_1 FILLER_26_820 ();
 sg13g2_fill_2 FILLER_26_827 ();
 sg13g2_fill_1 FILLER_26_829 ();
 sg13g2_fill_1 FILLER_26_835 ();
 sg13g2_fill_2 FILLER_26_849 ();
 sg13g2_decap_4 FILLER_26_856 ();
 sg13g2_decap_4 FILLER_26_863 ();
 sg13g2_decap_4 FILLER_26_873 ();
 sg13g2_fill_2 FILLER_26_877 ();
 sg13g2_decap_4 FILLER_26_883 ();
 sg13g2_fill_1 FILLER_26_887 ();
 sg13g2_decap_4 FILLER_26_893 ();
 sg13g2_fill_2 FILLER_26_897 ();
 sg13g2_fill_2 FILLER_26_903 ();
 sg13g2_fill_1 FILLER_26_905 ();
 sg13g2_fill_1 FILLER_26_932 ();
 sg13g2_fill_2 FILLER_26_982 ();
 sg13g2_fill_2 FILLER_26_992 ();
 sg13g2_fill_2 FILLER_26_1002 ();
 sg13g2_fill_1 FILLER_26_1031 ();
 sg13g2_decap_4 FILLER_26_1040 ();
 sg13g2_decap_8 FILLER_26_1048 ();
 sg13g2_decap_4 FILLER_26_1064 ();
 sg13g2_fill_2 FILLER_26_1085 ();
 sg13g2_fill_1 FILLER_26_1100 ();
 sg13g2_decap_4 FILLER_26_1133 ();
 sg13g2_fill_2 FILLER_26_1137 ();
 sg13g2_decap_8 FILLER_26_1208 ();
 sg13g2_fill_1 FILLER_26_1215 ();
 sg13g2_fill_2 FILLER_26_1220 ();
 sg13g2_fill_2 FILLER_26_1231 ();
 sg13g2_fill_1 FILLER_26_1233 ();
 sg13g2_decap_8 FILLER_26_1238 ();
 sg13g2_decap_4 FILLER_26_1245 ();
 sg13g2_fill_2 FILLER_26_1249 ();
 sg13g2_fill_2 FILLER_26_1278 ();
 sg13g2_fill_1 FILLER_26_1280 ();
 sg13g2_decap_8 FILLER_26_1325 ();
 sg13g2_decap_8 FILLER_26_1332 ();
 sg13g2_fill_2 FILLER_26_1378 ();
 sg13g2_decap_8 FILLER_26_1407 ();
 sg13g2_decap_4 FILLER_26_1427 ();
 sg13g2_fill_2 FILLER_26_1431 ();
 sg13g2_decap_8 FILLER_26_1437 ();
 sg13g2_fill_2 FILLER_26_1444 ();
 sg13g2_fill_1 FILLER_26_1446 ();
 sg13g2_decap_4 FILLER_26_1484 ();
 sg13g2_fill_2 FILLER_26_1488 ();
 sg13g2_decap_4 FILLER_26_1500 ();
 sg13g2_fill_1 FILLER_26_1504 ();
 sg13g2_decap_8 FILLER_26_1532 ();
 sg13g2_fill_1 FILLER_26_1557 ();
 sg13g2_decap_8 FILLER_26_1563 ();
 sg13g2_decap_4 FILLER_26_1610 ();
 sg13g2_fill_2 FILLER_26_1633 ();
 sg13g2_fill_1 FILLER_26_1635 ();
 sg13g2_fill_1 FILLER_26_1640 ();
 sg13g2_decap_4 FILLER_26_1656 ();
 sg13g2_decap_8 FILLER_26_1665 ();
 sg13g2_decap_8 FILLER_26_1672 ();
 sg13g2_decap_8 FILLER_26_1679 ();
 sg13g2_decap_8 FILLER_26_1686 ();
 sg13g2_decap_8 FILLER_26_1693 ();
 sg13g2_decap_8 FILLER_26_1700 ();
 sg13g2_decap_8 FILLER_26_1707 ();
 sg13g2_decap_8 FILLER_26_1714 ();
 sg13g2_decap_8 FILLER_26_1721 ();
 sg13g2_decap_8 FILLER_26_1728 ();
 sg13g2_decap_8 FILLER_26_1735 ();
 sg13g2_decap_8 FILLER_26_1742 ();
 sg13g2_decap_8 FILLER_26_1749 ();
 sg13g2_decap_8 FILLER_26_1756 ();
 sg13g2_decap_4 FILLER_26_1763 ();
 sg13g2_fill_1 FILLER_26_1767 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_fill_1 FILLER_27_34 ();
 sg13g2_decap_8 FILLER_27_116 ();
 sg13g2_decap_8 FILLER_27_123 ();
 sg13g2_decap_8 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_137 ();
 sg13g2_fill_1 FILLER_27_205 ();
 sg13g2_fill_2 FILLER_27_214 ();
 sg13g2_fill_1 FILLER_27_216 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_decap_4 FILLER_27_277 ();
 sg13g2_fill_2 FILLER_27_281 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_decap_4 FILLER_27_400 ();
 sg13g2_fill_2 FILLER_27_460 ();
 sg13g2_decap_4 FILLER_27_480 ();
 sg13g2_fill_2 FILLER_27_493 ();
 sg13g2_fill_2 FILLER_27_500 ();
 sg13g2_decap_4 FILLER_27_530 ();
 sg13g2_fill_1 FILLER_27_543 ();
 sg13g2_fill_1 FILLER_27_554 ();
 sg13g2_decap_4 FILLER_27_563 ();
 sg13g2_fill_2 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_587 ();
 sg13g2_fill_2 FILLER_27_594 ();
 sg13g2_fill_1 FILLER_27_624 ();
 sg13g2_fill_2 FILLER_27_629 ();
 sg13g2_fill_1 FILLER_27_631 ();
 sg13g2_decap_4 FILLER_27_678 ();
 sg13g2_fill_1 FILLER_27_682 ();
 sg13g2_fill_1 FILLER_27_715 ();
 sg13g2_fill_1 FILLER_27_750 ();
 sg13g2_fill_1 FILLER_27_762 ();
 sg13g2_decap_4 FILLER_27_772 ();
 sg13g2_decap_8 FILLER_27_788 ();
 sg13g2_decap_4 FILLER_27_829 ();
 sg13g2_fill_1 FILLER_27_833 ();
 sg13g2_decap_4 FILLER_27_860 ();
 sg13g2_fill_2 FILLER_27_963 ();
 sg13g2_fill_1 FILLER_27_965 ();
 sg13g2_fill_1 FILLER_27_1007 ();
 sg13g2_decap_4 FILLER_27_1021 ();
 sg13g2_fill_2 FILLER_27_1025 ();
 sg13g2_decap_8 FILLER_27_1055 ();
 sg13g2_fill_2 FILLER_27_1062 ();
 sg13g2_fill_1 FILLER_27_1064 ();
 sg13g2_fill_2 FILLER_27_1092 ();
 sg13g2_fill_1 FILLER_27_1094 ();
 sg13g2_decap_4 FILLER_27_1122 ();
 sg13g2_fill_1 FILLER_27_1126 ();
 sg13g2_fill_1 FILLER_27_1184 ();
 sg13g2_decap_4 FILLER_27_1194 ();
 sg13g2_decap_8 FILLER_27_1265 ();
 sg13g2_decap_4 FILLER_27_1308 ();
 sg13g2_fill_1 FILLER_27_1339 ();
 sg13g2_fill_2 FILLER_27_1403 ();
 sg13g2_fill_2 FILLER_27_1459 ();
 sg13g2_decap_4 FILLER_27_1481 ();
 sg13g2_fill_2 FILLER_27_1485 ();
 sg13g2_decap_4 FILLER_27_1526 ();
 sg13g2_fill_1 FILLER_27_1530 ();
 sg13g2_fill_2 FILLER_27_1556 ();
 sg13g2_fill_1 FILLER_27_1558 ();
 sg13g2_decap_8 FILLER_27_1591 ();
 sg13g2_decap_8 FILLER_27_1598 ();
 sg13g2_fill_2 FILLER_27_1605 ();
 sg13g2_fill_2 FILLER_27_1646 ();
 sg13g2_fill_1 FILLER_27_1673 ();
 sg13g2_decap_8 FILLER_27_1687 ();
 sg13g2_decap_8 FILLER_27_1694 ();
 sg13g2_decap_8 FILLER_27_1701 ();
 sg13g2_decap_8 FILLER_27_1708 ();
 sg13g2_decap_8 FILLER_27_1715 ();
 sg13g2_decap_8 FILLER_27_1722 ();
 sg13g2_decap_8 FILLER_27_1729 ();
 sg13g2_decap_8 FILLER_27_1736 ();
 sg13g2_decap_8 FILLER_27_1743 ();
 sg13g2_decap_8 FILLER_27_1750 ();
 sg13g2_decap_8 FILLER_27_1757 ();
 sg13g2_decap_4 FILLER_27_1764 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_58 ();
 sg13g2_fill_1 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_71 ();
 sg13g2_fill_1 FILLER_28_88 ();
 sg13g2_fill_2 FILLER_28_121 ();
 sg13g2_fill_2 FILLER_28_167 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_decap_8 FILLER_28_183 ();
 sg13g2_decap_4 FILLER_28_190 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_decap_4 FILLER_28_299 ();
 sg13g2_fill_2 FILLER_28_303 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_4 FILLER_28_317 ();
 sg13g2_decap_4 FILLER_28_329 ();
 sg13g2_fill_2 FILLER_28_333 ();
 sg13g2_fill_1 FILLER_28_358 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_412 ();
 sg13g2_fill_2 FILLER_28_422 ();
 sg13g2_decap_4 FILLER_28_433 ();
 sg13g2_decap_4 FILLER_28_441 ();
 sg13g2_fill_2 FILLER_28_471 ();
 sg13g2_fill_1 FILLER_28_473 ();
 sg13g2_fill_1 FILLER_28_487 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_fill_2 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_558 ();
 sg13g2_fill_2 FILLER_28_575 ();
 sg13g2_decap_8 FILLER_28_587 ();
 sg13g2_decap_4 FILLER_28_594 ();
 sg13g2_fill_2 FILLER_28_615 ();
 sg13g2_fill_2 FILLER_28_675 ();
 sg13g2_decap_4 FILLER_28_714 ();
 sg13g2_fill_1 FILLER_28_718 ();
 sg13g2_fill_1 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_752 ();
 sg13g2_decap_8 FILLER_28_759 ();
 sg13g2_decap_4 FILLER_28_766 ();
 sg13g2_fill_2 FILLER_28_778 ();
 sg13g2_fill_1 FILLER_28_780 ();
 sg13g2_fill_2 FILLER_28_798 ();
 sg13g2_decap_4 FILLER_28_804 ();
 sg13g2_fill_2 FILLER_28_808 ();
 sg13g2_decap_8 FILLER_28_814 ();
 sg13g2_decap_8 FILLER_28_821 ();
 sg13g2_fill_2 FILLER_28_828 ();
 sg13g2_decap_8 FILLER_28_834 ();
 sg13g2_fill_1 FILLER_28_841 ();
 sg13g2_fill_1 FILLER_28_857 ();
 sg13g2_decap_8 FILLER_28_862 ();
 sg13g2_decap_4 FILLER_28_869 ();
 sg13g2_fill_1 FILLER_28_873 ();
 sg13g2_fill_1 FILLER_28_883 ();
 sg13g2_fill_2 FILLER_28_893 ();
 sg13g2_decap_8 FILLER_28_916 ();
 sg13g2_fill_1 FILLER_28_982 ();
 sg13g2_fill_1 FILLER_28_988 ();
 sg13g2_decap_8 FILLER_28_1016 ();
 sg13g2_decap_4 FILLER_28_1023 ();
 sg13g2_fill_2 FILLER_28_1027 ();
 sg13g2_fill_1 FILLER_28_1038 ();
 sg13g2_decap_4 FILLER_28_1066 ();
 sg13g2_fill_1 FILLER_28_1074 ();
 sg13g2_decap_8 FILLER_28_1079 ();
 sg13g2_decap_4 FILLER_28_1086 ();
 sg13g2_fill_2 FILLER_28_1112 ();
 sg13g2_fill_2 FILLER_28_1145 ();
 sg13g2_fill_2 FILLER_28_1183 ();
 sg13g2_decap_8 FILLER_28_1212 ();
 sg13g2_decap_4 FILLER_28_1219 ();
 sg13g2_fill_1 FILLER_28_1223 ();
 sg13g2_fill_2 FILLER_28_1269 ();
 sg13g2_fill_1 FILLER_28_1271 ();
 sg13g2_fill_2 FILLER_28_1289 ();
 sg13g2_fill_1 FILLER_28_1291 ();
 sg13g2_fill_2 FILLER_28_1359 ();
 sg13g2_fill_2 FILLER_28_1383 ();
 sg13g2_fill_2 FILLER_28_1389 ();
 sg13g2_fill_2 FILLER_28_1404 ();
 sg13g2_fill_2 FILLER_28_1423 ();
 sg13g2_fill_1 FILLER_28_1425 ();
 sg13g2_fill_2 FILLER_28_1445 ();
 sg13g2_fill_1 FILLER_28_1447 ();
 sg13g2_decap_8 FILLER_28_1458 ();
 sg13g2_fill_1 FILLER_28_1484 ();
 sg13g2_decap_8 FILLER_28_1489 ();
 sg13g2_fill_2 FILLER_28_1496 ();
 sg13g2_fill_1 FILLER_28_1498 ();
 sg13g2_fill_2 FILLER_28_1503 ();
 sg13g2_fill_1 FILLER_28_1505 ();
 sg13g2_decap_4 FILLER_28_1511 ();
 sg13g2_fill_1 FILLER_28_1515 ();
 sg13g2_decap_8 FILLER_28_1531 ();
 sg13g2_fill_1 FILLER_28_1538 ();
 sg13g2_decap_4 FILLER_28_1549 ();
 sg13g2_decap_8 FILLER_28_1558 ();
 sg13g2_decap_4 FILLER_28_1565 ();
 sg13g2_fill_1 FILLER_28_1569 ();
 sg13g2_decap_8 FILLER_28_1583 ();
 sg13g2_fill_1 FILLER_28_1590 ();
 sg13g2_decap_4 FILLER_28_1601 ();
 sg13g2_fill_1 FILLER_28_1605 ();
 sg13g2_decap_8 FILLER_28_1611 ();
 sg13g2_fill_1 FILLER_28_1618 ();
 sg13g2_fill_1 FILLER_28_1630 ();
 sg13g2_decap_4 FILLER_28_1635 ();
 sg13g2_fill_1 FILLER_28_1660 ();
 sg13g2_decap_4 FILLER_28_1689 ();
 sg13g2_decap_8 FILLER_28_1701 ();
 sg13g2_decap_8 FILLER_28_1708 ();
 sg13g2_decap_8 FILLER_28_1715 ();
 sg13g2_decap_8 FILLER_28_1722 ();
 sg13g2_decap_8 FILLER_28_1729 ();
 sg13g2_decap_8 FILLER_28_1736 ();
 sg13g2_decap_8 FILLER_28_1743 ();
 sg13g2_decap_8 FILLER_28_1750 ();
 sg13g2_decap_8 FILLER_28_1757 ();
 sg13g2_decap_4 FILLER_28_1764 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_107 ();
 sg13g2_fill_2 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_170 ();
 sg13g2_decap_4 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_191 ();
 sg13g2_fill_1 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_218 ();
 sg13g2_decap_8 FILLER_29_260 ();
 sg13g2_fill_2 FILLER_29_267 ();
 sg13g2_fill_1 FILLER_29_286 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_decap_8 FILLER_29_323 ();
 sg13g2_decap_8 FILLER_29_330 ();
 sg13g2_fill_2 FILLER_29_337 ();
 sg13g2_fill_2 FILLER_29_348 ();
 sg13g2_fill_2 FILLER_29_385 ();
 sg13g2_fill_2 FILLER_29_397 ();
 sg13g2_fill_1 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_440 ();
 sg13g2_decap_8 FILLER_29_447 ();
 sg13g2_decap_4 FILLER_29_454 ();
 sg13g2_fill_1 FILLER_29_480 ();
 sg13g2_fill_2 FILLER_29_496 ();
 sg13g2_decap_8 FILLER_29_512 ();
 sg13g2_decap_4 FILLER_29_519 ();
 sg13g2_fill_1 FILLER_29_536 ();
 sg13g2_decap_4 FILLER_29_555 ();
 sg13g2_fill_1 FILLER_29_582 ();
 sg13g2_decap_8 FILLER_29_588 ();
 sg13g2_decap_4 FILLER_29_595 ();
 sg13g2_fill_1 FILLER_29_599 ();
 sg13g2_fill_1 FILLER_29_605 ();
 sg13g2_fill_2 FILLER_29_611 ();
 sg13g2_fill_1 FILLER_29_622 ();
 sg13g2_fill_1 FILLER_29_627 ();
 sg13g2_decap_4 FILLER_29_639 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_fill_2 FILLER_29_704 ();
 sg13g2_fill_1 FILLER_29_706 ();
 sg13g2_fill_1 FILLER_29_719 ();
 sg13g2_fill_1 FILLER_29_753 ();
 sg13g2_decap_4 FILLER_29_759 ();
 sg13g2_fill_1 FILLER_29_763 ();
 sg13g2_decap_4 FILLER_29_795 ();
 sg13g2_fill_1 FILLER_29_799 ();
 sg13g2_fill_2 FILLER_29_809 ();
 sg13g2_fill_2 FILLER_29_883 ();
 sg13g2_fill_2 FILLER_29_903 ();
 sg13g2_fill_1 FILLER_29_905 ();
 sg13g2_fill_1 FILLER_29_919 ();
 sg13g2_fill_2 FILLER_29_981 ();
 sg13g2_fill_1 FILLER_29_983 ();
 sg13g2_decap_4 FILLER_29_1029 ();
 sg13g2_fill_1 FILLER_29_1033 ();
 sg13g2_decap_8 FILLER_29_1055 ();
 sg13g2_decap_8 FILLER_29_1062 ();
 sg13g2_fill_2 FILLER_29_1097 ();
 sg13g2_fill_2 FILLER_29_1166 ();
 sg13g2_fill_1 FILLER_29_1168 ();
 sg13g2_decap_4 FILLER_29_1200 ();
 sg13g2_fill_2 FILLER_29_1204 ();
 sg13g2_fill_2 FILLER_29_1246 ();
 sg13g2_fill_2 FILLER_29_1265 ();
 sg13g2_fill_1 FILLER_29_1343 ();
 sg13g2_fill_1 FILLER_29_1380 ();
 sg13g2_decap_4 FILLER_29_1435 ();
 sg13g2_fill_2 FILLER_29_1439 ();
 sg13g2_fill_2 FILLER_29_1471 ();
 sg13g2_fill_1 FILLER_29_1473 ();
 sg13g2_fill_1 FILLER_29_1509 ();
 sg13g2_fill_1 FILLER_29_1530 ();
 sg13g2_decap_4 FILLER_29_1590 ();
 sg13g2_fill_2 FILLER_29_1594 ();
 sg13g2_fill_2 FILLER_29_1617 ();
 sg13g2_decap_8 FILLER_29_1639 ();
 sg13g2_decap_8 FILLER_29_1646 ();
 sg13g2_decap_8 FILLER_29_1653 ();
 sg13g2_fill_2 FILLER_29_1674 ();
 sg13g2_fill_1 FILLER_29_1676 ();
 sg13g2_fill_1 FILLER_29_1681 ();
 sg13g2_decap_8 FILLER_29_1686 ();
 sg13g2_decap_8 FILLER_29_1693 ();
 sg13g2_decap_8 FILLER_29_1724 ();
 sg13g2_decap_8 FILLER_29_1731 ();
 sg13g2_decap_8 FILLER_29_1738 ();
 sg13g2_decap_8 FILLER_29_1745 ();
 sg13g2_decap_8 FILLER_29_1752 ();
 sg13g2_decap_8 FILLER_29_1759 ();
 sg13g2_fill_2 FILLER_29_1766 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_4 ();
 sg13g2_fill_2 FILLER_30_10 ();
 sg13g2_fill_1 FILLER_30_12 ();
 sg13g2_decap_4 FILLER_30_22 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_56 ();
 sg13g2_fill_2 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_145 ();
 sg13g2_fill_2 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_209 ();
 sg13g2_fill_1 FILLER_30_211 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_260 ();
 sg13g2_decap_4 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_336 ();
 sg13g2_fill_2 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_fill_2 FILLER_30_361 ();
 sg13g2_fill_1 FILLER_30_363 ();
 sg13g2_fill_1 FILLER_30_413 ();
 sg13g2_fill_2 FILLER_30_419 ();
 sg13g2_fill_2 FILLER_30_462 ();
 sg13g2_decap_4 FILLER_30_482 ();
 sg13g2_decap_8 FILLER_30_505 ();
 sg13g2_decap_4 FILLER_30_512 ();
 sg13g2_fill_1 FILLER_30_516 ();
 sg13g2_fill_2 FILLER_30_558 ();
 sg13g2_fill_1 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_566 ();
 sg13g2_fill_1 FILLER_30_591 ();
 sg13g2_fill_1 FILLER_30_629 ();
 sg13g2_fill_2 FILLER_30_646 ();
 sg13g2_decap_4 FILLER_30_652 ();
 sg13g2_fill_1 FILLER_30_656 ();
 sg13g2_decap_4 FILLER_30_669 ();
 sg13g2_fill_1 FILLER_30_673 ();
 sg13g2_fill_2 FILLER_30_715 ();
 sg13g2_fill_1 FILLER_30_717 ();
 sg13g2_fill_2 FILLER_30_732 ();
 sg13g2_fill_1 FILLER_30_734 ();
 sg13g2_fill_1 FILLER_30_755 ();
 sg13g2_fill_2 FILLER_30_761 ();
 sg13g2_fill_1 FILLER_30_763 ();
 sg13g2_decap_4 FILLER_30_780 ();
 sg13g2_fill_2 FILLER_30_788 ();
 sg13g2_fill_1 FILLER_30_790 ();
 sg13g2_fill_2 FILLER_30_837 ();
 sg13g2_fill_2 FILLER_30_887 ();
 sg13g2_fill_2 FILLER_30_966 ();
 sg13g2_fill_1 FILLER_30_1016 ();
 sg13g2_fill_1 FILLER_30_1129 ();
 sg13g2_fill_1 FILLER_30_1139 ();
 sg13g2_fill_1 FILLER_30_1157 ();
 sg13g2_fill_2 FILLER_30_1207 ();
 sg13g2_fill_2 FILLER_30_1222 ();
 sg13g2_fill_2 FILLER_30_1241 ();
 sg13g2_fill_1 FILLER_30_1243 ();
 sg13g2_fill_2 FILLER_30_1361 ();
 sg13g2_decap_4 FILLER_30_1403 ();
 sg13g2_fill_1 FILLER_30_1407 ();
 sg13g2_decap_8 FILLER_30_1432 ();
 sg13g2_decap_8 FILLER_30_1439 ();
 sg13g2_fill_2 FILLER_30_1446 ();
 sg13g2_decap_8 FILLER_30_1471 ();
 sg13g2_decap_4 FILLER_30_1478 ();
 sg13g2_decap_8 FILLER_30_1492 ();
 sg13g2_decap_8 FILLER_30_1499 ();
 sg13g2_decap_8 FILLER_30_1506 ();
 sg13g2_fill_2 FILLER_30_1513 ();
 sg13g2_decap_8 FILLER_30_1529 ();
 sg13g2_fill_2 FILLER_30_1536 ();
 sg13g2_fill_2 FILLER_30_1549 ();
 sg13g2_decap_8 FILLER_30_1557 ();
 sg13g2_decap_4 FILLER_30_1564 ();
 sg13g2_fill_2 FILLER_30_1589 ();
 sg13g2_fill_1 FILLER_30_1605 ();
 sg13g2_decap_8 FILLER_30_1615 ();
 sg13g2_decap_8 FILLER_30_1641 ();
 sg13g2_fill_1 FILLER_30_1648 ();
 sg13g2_decap_8 FILLER_30_1661 ();
 sg13g2_fill_2 FILLER_30_1668 ();
 sg13g2_fill_1 FILLER_30_1676 ();
 sg13g2_decap_8 FILLER_30_1689 ();
 sg13g2_fill_1 FILLER_30_1696 ();
 sg13g2_decap_4 FILLER_30_1710 ();
 sg13g2_fill_2 FILLER_30_1714 ();
 sg13g2_decap_8 FILLER_30_1736 ();
 sg13g2_decap_8 FILLER_30_1743 ();
 sg13g2_decap_8 FILLER_30_1750 ();
 sg13g2_decap_8 FILLER_30_1757 ();
 sg13g2_decap_4 FILLER_30_1764 ();
 sg13g2_fill_1 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_39 ();
 sg13g2_fill_1 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_52 ();
 sg13g2_fill_1 FILLER_31_54 ();
 sg13g2_decap_8 FILLER_31_115 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_4 FILLER_31_133 ();
 sg13g2_fill_2 FILLER_31_137 ();
 sg13g2_decap_8 FILLER_31_167 ();
 sg13g2_fill_1 FILLER_31_174 ();
 sg13g2_decap_4 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_fill_1 FILLER_31_223 ();
 sg13g2_decap_8 FILLER_31_260 ();
 sg13g2_decap_4 FILLER_31_267 ();
 sg13g2_fill_2 FILLER_31_271 ();
 sg13g2_decap_4 FILLER_31_285 ();
 sg13g2_fill_2 FILLER_31_289 ();
 sg13g2_fill_1 FILLER_31_309 ();
 sg13g2_decap_8 FILLER_31_323 ();
 sg13g2_fill_1 FILLER_31_330 ();
 sg13g2_decap_8 FILLER_31_341 ();
 sg13g2_decap_4 FILLER_31_354 ();
 sg13g2_decap_8 FILLER_31_386 ();
 sg13g2_fill_1 FILLER_31_393 ();
 sg13g2_fill_2 FILLER_31_398 ();
 sg13g2_fill_1 FILLER_31_400 ();
 sg13g2_fill_2 FILLER_31_414 ();
 sg13g2_fill_1 FILLER_31_416 ();
 sg13g2_fill_1 FILLER_31_422 ();
 sg13g2_fill_1 FILLER_31_438 ();
 sg13g2_decap_8 FILLER_31_443 ();
 sg13g2_decap_4 FILLER_31_450 ();
 sg13g2_decap_8 FILLER_31_480 ();
 sg13g2_decap_8 FILLER_31_487 ();
 sg13g2_decap_4 FILLER_31_494 ();
 sg13g2_decap_4 FILLER_31_563 ();
 sg13g2_fill_1 FILLER_31_596 ();
 sg13g2_decap_4 FILLER_31_601 ();
 sg13g2_fill_1 FILLER_31_605 ();
 sg13g2_decap_8 FILLER_31_610 ();
 sg13g2_decap_8 FILLER_31_617 ();
 sg13g2_decap_4 FILLER_31_633 ();
 sg13g2_fill_2 FILLER_31_646 ();
 sg13g2_fill_1 FILLER_31_661 ();
 sg13g2_decap_4 FILLER_31_680 ();
 sg13g2_fill_2 FILLER_31_688 ();
 sg13g2_fill_1 FILLER_31_718 ();
 sg13g2_fill_2 FILLER_31_757 ();
 sg13g2_decap_4 FILLER_31_772 ();
 sg13g2_decap_4 FILLER_31_781 ();
 sg13g2_decap_8 FILLER_31_795 ();
 sg13g2_fill_2 FILLER_31_802 ();
 sg13g2_fill_1 FILLER_31_831 ();
 sg13g2_fill_1 FILLER_31_866 ();
 sg13g2_fill_1 FILLER_31_888 ();
 sg13g2_decap_4 FILLER_31_925 ();
 sg13g2_fill_1 FILLER_31_929 ();
 sg13g2_fill_1 FILLER_31_995 ();
 sg13g2_decap_4 FILLER_31_1018 ();
 sg13g2_decap_8 FILLER_31_1026 ();
 sg13g2_decap_4 FILLER_31_1033 ();
 sg13g2_decap_4 FILLER_31_1063 ();
 sg13g2_decap_4 FILLER_31_1085 ();
 sg13g2_fill_1 FILLER_31_1089 ();
 sg13g2_decap_8 FILLER_31_1112 ();
 sg13g2_fill_1 FILLER_31_1119 ();
 sg13g2_fill_2 FILLER_31_1187 ();
 sg13g2_fill_1 FILLER_31_1189 ();
 sg13g2_decap_8 FILLER_31_1245 ();
 sg13g2_fill_2 FILLER_31_1252 ();
 sg13g2_fill_1 FILLER_31_1254 ();
 sg13g2_fill_1 FILLER_31_1268 ();
 sg13g2_fill_2 FILLER_31_1299 ();
 sg13g2_decap_8 FILLER_31_1305 ();
 sg13g2_fill_1 FILLER_31_1312 ();
 sg13g2_decap_4 FILLER_31_1334 ();
 sg13g2_fill_2 FILLER_31_1338 ();
 sg13g2_fill_2 FILLER_31_1357 ();
 sg13g2_decap_4 FILLER_31_1363 ();
 sg13g2_fill_2 FILLER_31_1380 ();
 sg13g2_fill_2 FILLER_31_1395 ();
 sg13g2_fill_1 FILLER_31_1397 ();
 sg13g2_fill_2 FILLER_31_1406 ();
 sg13g2_fill_1 FILLER_31_1408 ();
 sg13g2_fill_1 FILLER_31_1424 ();
 sg13g2_decap_8 FILLER_31_1440 ();
 sg13g2_fill_2 FILLER_31_1447 ();
 sg13g2_fill_1 FILLER_31_1449 ();
 sg13g2_fill_1 FILLER_31_1456 ();
 sg13g2_decap_8 FILLER_31_1477 ();
 sg13g2_fill_2 FILLER_31_1484 ();
 sg13g2_fill_1 FILLER_31_1486 ();
 sg13g2_fill_2 FILLER_31_1537 ();
 sg13g2_decap_8 FILLER_31_1560 ();
 sg13g2_fill_1 FILLER_31_1567 ();
 sg13g2_decap_4 FILLER_31_1589 ();
 sg13g2_fill_1 FILLER_31_1593 ();
 sg13g2_fill_1 FILLER_31_1609 ();
 sg13g2_decap_4 FILLER_31_1615 ();
 sg13g2_fill_1 FILLER_31_1624 ();
 sg13g2_fill_1 FILLER_31_1631 ();
 sg13g2_fill_2 FILLER_31_1643 ();
 sg13g2_fill_2 FILLER_31_1667 ();
 sg13g2_decap_8 FILLER_31_1689 ();
 sg13g2_fill_1 FILLER_31_1696 ();
 sg13g2_decap_8 FILLER_31_1701 ();
 sg13g2_decap_4 FILLER_31_1708 ();
 sg13g2_fill_2 FILLER_31_1712 ();
 sg13g2_decap_8 FILLER_31_1743 ();
 sg13g2_decap_8 FILLER_31_1750 ();
 sg13g2_decap_8 FILLER_31_1757 ();
 sg13g2_decap_4 FILLER_31_1764 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_16 ();
 sg13g2_fill_1 FILLER_32_44 ();
 sg13g2_decap_4 FILLER_32_78 ();
 sg13g2_fill_2 FILLER_32_82 ();
 sg13g2_fill_1 FILLER_32_115 ();
 sg13g2_fill_2 FILLER_32_168 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_fill_1 FILLER_32_176 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_2 FILLER_32_238 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_260 ();
 sg13g2_fill_1 FILLER_32_262 ();
 sg13g2_decap_8 FILLER_32_285 ();
 sg13g2_decap_4 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_296 ();
 sg13g2_decap_4 FILLER_32_321 ();
 sg13g2_fill_2 FILLER_32_338 ();
 sg13g2_decap_4 FILLER_32_346 ();
 sg13g2_decap_4 FILLER_32_364 ();
 sg13g2_fill_1 FILLER_32_368 ();
 sg13g2_fill_1 FILLER_32_374 ();
 sg13g2_decap_8 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_413 ();
 sg13g2_fill_2 FILLER_32_420 ();
 sg13g2_fill_1 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_432 ();
 sg13g2_fill_2 FILLER_32_451 ();
 sg13g2_decap_4 FILLER_32_484 ();
 sg13g2_fill_2 FILLER_32_488 ();
 sg13g2_fill_2 FILLER_32_507 ();
 sg13g2_fill_2 FILLER_32_522 ();
 sg13g2_decap_8 FILLER_32_547 ();
 sg13g2_decap_8 FILLER_32_554 ();
 sg13g2_decap_4 FILLER_32_561 ();
 sg13g2_fill_1 FILLER_32_565 ();
 sg13g2_fill_1 FILLER_32_577 ();
 sg13g2_decap_8 FILLER_32_590 ();
 sg13g2_fill_2 FILLER_32_597 ();
 sg13g2_decap_4 FILLER_32_603 ();
 sg13g2_fill_2 FILLER_32_607 ();
 sg13g2_fill_2 FILLER_32_646 ();
 sg13g2_decap_4 FILLER_32_679 ();
 sg13g2_fill_2 FILLER_32_683 ();
 sg13g2_fill_1 FILLER_32_707 ();
 sg13g2_fill_2 FILLER_32_716 ();
 sg13g2_fill_2 FILLER_32_731 ();
 sg13g2_fill_1 FILLER_32_733 ();
 sg13g2_fill_1 FILLER_32_762 ();
 sg13g2_fill_2 FILLER_32_809 ();
 sg13g2_fill_1 FILLER_32_901 ();
 sg13g2_fill_1 FILLER_32_924 ();
 sg13g2_fill_1 FILLER_32_972 ();
 sg13g2_decap_8 FILLER_32_1014 ();
 sg13g2_decap_4 FILLER_32_1021 ();
 sg13g2_fill_2 FILLER_32_1025 ();
 sg13g2_decap_8 FILLER_32_1031 ();
 sg13g2_fill_2 FILLER_32_1038 ();
 sg13g2_fill_1 FILLER_32_1040 ();
 sg13g2_fill_2 FILLER_32_1069 ();
 sg13g2_fill_1 FILLER_32_1071 ();
 sg13g2_fill_2 FILLER_32_1157 ();
 sg13g2_decap_4 FILLER_32_1185 ();
 sg13g2_fill_2 FILLER_32_1216 ();
 sg13g2_fill_1 FILLER_32_1218 ();
 sg13g2_decap_8 FILLER_32_1223 ();
 sg13g2_decap_4 FILLER_32_1230 ();
 sg13g2_fill_2 FILLER_32_1234 ();
 sg13g2_fill_2 FILLER_32_1398 ();
 sg13g2_fill_1 FILLER_32_1413 ();
 sg13g2_fill_2 FILLER_32_1421 ();
 sg13g2_fill_1 FILLER_32_1423 ();
 sg13g2_decap_8 FILLER_32_1431 ();
 sg13g2_fill_1 FILLER_32_1438 ();
 sg13g2_decap_4 FILLER_32_1444 ();
 sg13g2_fill_2 FILLER_32_1448 ();
 sg13g2_decap_8 FILLER_32_1460 ();
 sg13g2_decap_4 FILLER_32_1484 ();
 sg13g2_fill_1 FILLER_32_1488 ();
 sg13g2_decap_8 FILLER_32_1495 ();
 sg13g2_decap_8 FILLER_32_1502 ();
 sg13g2_decap_8 FILLER_32_1509 ();
 sg13g2_decap_8 FILLER_32_1535 ();
 sg13g2_fill_1 FILLER_32_1542 ();
 sg13g2_decap_8 FILLER_32_1553 ();
 sg13g2_decap_8 FILLER_32_1565 ();
 sg13g2_fill_1 FILLER_32_1572 ();
 sg13g2_decap_8 FILLER_32_1583 ();
 sg13g2_fill_2 FILLER_32_1590 ();
 sg13g2_fill_1 FILLER_32_1592 ();
 sg13g2_fill_2 FILLER_32_1598 ();
 sg13g2_fill_1 FILLER_32_1617 ();
 sg13g2_fill_2 FILLER_32_1623 ();
 sg13g2_fill_2 FILLER_32_1633 ();
 sg13g2_fill_1 FILLER_32_1640 ();
 sg13g2_decap_8 FILLER_32_1645 ();
 sg13g2_decap_4 FILLER_32_1652 ();
 sg13g2_decap_8 FILLER_32_1664 ();
 sg13g2_decap_4 FILLER_32_1675 ();
 sg13g2_decap_4 FILLER_32_1687 ();
 sg13g2_fill_1 FILLER_32_1691 ();
 sg13g2_decap_8 FILLER_32_1709 ();
 sg13g2_decap_4 FILLER_32_1716 ();
 sg13g2_fill_1 FILLER_32_1720 ();
 sg13g2_decap_8 FILLER_32_1741 ();
 sg13g2_decap_8 FILLER_32_1748 ();
 sg13g2_decap_8 FILLER_32_1755 ();
 sg13g2_decap_4 FILLER_32_1762 ();
 sg13g2_fill_2 FILLER_32_1766 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_106 ();
 sg13g2_decap_4 FILLER_33_123 ();
 sg13g2_decap_8 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_142 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_decap_4 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_170 ();
 sg13g2_decap_4 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_183 ();
 sg13g2_decap_8 FILLER_33_192 ();
 sg13g2_fill_2 FILLER_33_199 ();
 sg13g2_fill_1 FILLER_33_201 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_234 ();
 sg13g2_fill_2 FILLER_33_240 ();
 sg13g2_fill_2 FILLER_33_259 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_decap_4 FILLER_33_280 ();
 sg13g2_decap_4 FILLER_33_296 ();
 sg13g2_decap_4 FILLER_33_306 ();
 sg13g2_decap_4 FILLER_33_325 ();
 sg13g2_fill_1 FILLER_33_329 ();
 sg13g2_fill_2 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_377 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_4 FILLER_33_394 ();
 sg13g2_fill_1 FILLER_33_398 ();
 sg13g2_decap_4 FILLER_33_419 ();
 sg13g2_fill_2 FILLER_33_435 ();
 sg13g2_decap_8 FILLER_33_445 ();
 sg13g2_fill_2 FILLER_33_452 ();
 sg13g2_fill_2 FILLER_33_459 ();
 sg13g2_fill_2 FILLER_33_473 ();
 sg13g2_decap_8 FILLER_33_488 ();
 sg13g2_decap_8 FILLER_33_495 ();
 sg13g2_decap_8 FILLER_33_502 ();
 sg13g2_fill_2 FILLER_33_509 ();
 sg13g2_fill_1 FILLER_33_511 ();
 sg13g2_fill_1 FILLER_33_571 ();
 sg13g2_decap_4 FILLER_33_580 ();
 sg13g2_fill_2 FILLER_33_592 ();
 sg13g2_fill_1 FILLER_33_639 ();
 sg13g2_fill_1 FILLER_33_649 ();
 sg13g2_fill_2 FILLER_33_654 ();
 sg13g2_fill_2 FILLER_33_669 ();
 sg13g2_fill_1 FILLER_33_671 ();
 sg13g2_fill_2 FILLER_33_681 ();
 sg13g2_decap_4 FILLER_33_744 ();
 sg13g2_fill_2 FILLER_33_748 ();
 sg13g2_decap_8 FILLER_33_768 ();
 sg13g2_fill_2 FILLER_33_779 ();
 sg13g2_decap_4 FILLER_33_795 ();
 sg13g2_fill_1 FILLER_33_808 ();
 sg13g2_decap_4 FILLER_33_817 ();
 sg13g2_fill_2 FILLER_33_830 ();
 sg13g2_fill_1 FILLER_33_832 ();
 sg13g2_fill_1 FILLER_33_862 ();
 sg13g2_fill_2 FILLER_33_872 ();
 sg13g2_fill_1 FILLER_33_874 ();
 sg13g2_fill_2 FILLER_33_909 ();
 sg13g2_fill_2 FILLER_33_924 ();
 sg13g2_fill_2 FILLER_33_971 ();
 sg13g2_fill_2 FILLER_33_986 ();
 sg13g2_fill_1 FILLER_33_988 ();
 sg13g2_decap_4 FILLER_33_1154 ();
 sg13g2_fill_1 FILLER_33_1158 ();
 sg13g2_fill_2 FILLER_33_1186 ();
 sg13g2_decap_8 FILLER_33_1205 ();
 sg13g2_fill_1 FILLER_33_1240 ();
 sg13g2_fill_2 FILLER_33_1254 ();
 sg13g2_decap_8 FILLER_33_1282 ();
 sg13g2_decap_8 FILLER_33_1289 ();
 sg13g2_decap_4 FILLER_33_1296 ();
 sg13g2_fill_1 FILLER_33_1300 ();
 sg13g2_decap_8 FILLER_33_1321 ();
 sg13g2_decap_8 FILLER_33_1328 ();
 sg13g2_fill_2 FILLER_33_1335 ();
 sg13g2_fill_1 FILLER_33_1342 ();
 sg13g2_decap_8 FILLER_33_1348 ();
 sg13g2_decap_4 FILLER_33_1355 ();
 sg13g2_fill_2 FILLER_33_1364 ();
 sg13g2_fill_1 FILLER_33_1366 ();
 sg13g2_decap_8 FILLER_33_1371 ();
 sg13g2_decap_8 FILLER_33_1378 ();
 sg13g2_decap_8 FILLER_33_1385 ();
 sg13g2_fill_2 FILLER_33_1392 ();
 sg13g2_fill_1 FILLER_33_1394 ();
 sg13g2_fill_2 FILLER_33_1412 ();
 sg13g2_fill_1 FILLER_33_1427 ();
 sg13g2_fill_2 FILLER_33_1432 ();
 sg13g2_fill_2 FILLER_33_1442 ();
 sg13g2_decap_8 FILLER_33_1465 ();
 sg13g2_decap_4 FILLER_33_1472 ();
 sg13g2_fill_1 FILLER_33_1476 ();
 sg13g2_decap_8 FILLER_33_1483 ();
 sg13g2_fill_2 FILLER_33_1500 ();
 sg13g2_decap_4 FILLER_33_1528 ();
 sg13g2_fill_2 FILLER_33_1532 ();
 sg13g2_fill_1 FILLER_33_1544 ();
 sg13g2_fill_2 FILLER_33_1558 ();
 sg13g2_fill_1 FILLER_33_1560 ();
 sg13g2_decap_4 FILLER_33_1581 ();
 sg13g2_decap_4 FILLER_33_1621 ();
 sg13g2_fill_1 FILLER_33_1625 ();
 sg13g2_fill_1 FILLER_33_1638 ();
 sg13g2_decap_4 FILLER_33_1652 ();
 sg13g2_fill_1 FILLER_33_1656 ();
 sg13g2_decap_4 FILLER_33_1673 ();
 sg13g2_decap_4 FILLER_33_1697 ();
 sg13g2_decap_8 FILLER_33_1735 ();
 sg13g2_fill_2 FILLER_33_1742 ();
 sg13g2_fill_1 FILLER_33_1744 ();
 sg13g2_decap_8 FILLER_33_1748 ();
 sg13g2_decap_8 FILLER_33_1755 ();
 sg13g2_decap_4 FILLER_33_1762 ();
 sg13g2_fill_2 FILLER_33_1766 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_29 ();
 sg13g2_fill_1 FILLER_34_31 ();
 sg13g2_decap_8 FILLER_34_59 ();
 sg13g2_fill_2 FILLER_34_66 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_4 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_fill_2 FILLER_34_171 ();
 sg13g2_fill_1 FILLER_34_173 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_254 ();
 sg13g2_fill_2 FILLER_34_290 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_fill_1 FILLER_34_308 ();
 sg13g2_fill_2 FILLER_34_320 ();
 sg13g2_fill_2 FILLER_34_357 ();
 sg13g2_fill_1 FILLER_34_359 ();
 sg13g2_fill_1 FILLER_34_371 ();
 sg13g2_fill_2 FILLER_34_388 ();
 sg13g2_fill_1 FILLER_34_399 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_decap_4 FILLER_34_419 ();
 sg13g2_fill_1 FILLER_34_423 ();
 sg13g2_fill_2 FILLER_34_437 ();
 sg13g2_decap_8 FILLER_34_443 ();
 sg13g2_fill_2 FILLER_34_450 ();
 sg13g2_fill_1 FILLER_34_452 ();
 sg13g2_decap_8 FILLER_34_457 ();
 sg13g2_decap_8 FILLER_34_464 ();
 sg13g2_decap_4 FILLER_34_471 ();
 sg13g2_fill_1 FILLER_34_475 ();
 sg13g2_decap_4 FILLER_34_522 ();
 sg13g2_fill_2 FILLER_34_550 ();
 sg13g2_fill_1 FILLER_34_552 ();
 sg13g2_fill_2 FILLER_34_570 ();
 sg13g2_fill_2 FILLER_34_577 ();
 sg13g2_fill_1 FILLER_34_579 ();
 sg13g2_decap_8 FILLER_34_588 ();
 sg13g2_decap_4 FILLER_34_595 ();
 sg13g2_fill_2 FILLER_34_681 ();
 sg13g2_fill_2 FILLER_34_695 ();
 sg13g2_decap_4 FILLER_34_766 ();
 sg13g2_fill_2 FILLER_34_806 ();
 sg13g2_decap_4 FILLER_34_848 ();
 sg13g2_fill_1 FILLER_34_852 ();
 sg13g2_decap_4 FILLER_34_880 ();
 sg13g2_fill_2 FILLER_34_884 ();
 sg13g2_fill_2 FILLER_34_940 ();
 sg13g2_fill_1 FILLER_34_942 ();
 sg13g2_fill_1 FILLER_34_956 ();
 sg13g2_fill_1 FILLER_34_1002 ();
 sg13g2_fill_2 FILLER_34_1027 ();
 sg13g2_fill_1 FILLER_34_1029 ();
 sg13g2_decap_8 FILLER_34_1034 ();
 sg13g2_decap_8 FILLER_34_1041 ();
 sg13g2_decap_4 FILLER_34_1048 ();
 sg13g2_decap_4 FILLER_34_1069 ();
 sg13g2_fill_1 FILLER_34_1073 ();
 sg13g2_fill_1 FILLER_34_1141 ();
 sg13g2_decap_4 FILLER_34_1209 ();
 sg13g2_fill_1 FILLER_34_1213 ();
 sg13g2_decap_8 FILLER_34_1227 ();
 sg13g2_decap_4 FILLER_34_1234 ();
 sg13g2_fill_2 FILLER_34_1238 ();
 sg13g2_fill_2 FILLER_34_1263 ();
 sg13g2_decap_4 FILLER_34_1308 ();
 sg13g2_fill_1 FILLER_34_1339 ();
 sg13g2_fill_2 FILLER_34_1355 ();
 sg13g2_fill_1 FILLER_34_1357 ();
 sg13g2_decap_8 FILLER_34_1381 ();
 sg13g2_decap_8 FILLER_34_1388 ();
 sg13g2_fill_1 FILLER_34_1395 ();
 sg13g2_decap_4 FILLER_34_1437 ();
 sg13g2_decap_4 FILLER_34_1457 ();
 sg13g2_fill_1 FILLER_34_1484 ();
 sg13g2_decap_8 FILLER_34_1493 ();
 sg13g2_decap_4 FILLER_34_1524 ();
 sg13g2_fill_2 FILLER_34_1549 ();
 sg13g2_fill_2 FILLER_34_1556 ();
 sg13g2_fill_1 FILLER_34_1568 ();
 sg13g2_decap_8 FILLER_34_1579 ();
 sg13g2_decap_8 FILLER_34_1586 ();
 sg13g2_decap_8 FILLER_34_1593 ();
 sg13g2_fill_2 FILLER_34_1600 ();
 sg13g2_fill_2 FILLER_34_1623 ();
 sg13g2_decap_4 FILLER_34_1633 ();
 sg13g2_fill_1 FILLER_34_1637 ();
 sg13g2_decap_8 FILLER_34_1644 ();
 sg13g2_decap_8 FILLER_34_1651 ();
 sg13g2_fill_2 FILLER_34_1658 ();
 sg13g2_decap_8 FILLER_34_1686 ();
 sg13g2_fill_2 FILLER_34_1693 ();
 sg13g2_fill_1 FILLER_34_1695 ();
 sg13g2_decap_8 FILLER_34_1717 ();
 sg13g2_fill_2 FILLER_34_1724 ();
 sg13g2_fill_2 FILLER_34_1729 ();
 sg13g2_fill_2 FILLER_34_1743 ();
 sg13g2_decap_8 FILLER_34_1757 ();
 sg13g2_decap_4 FILLER_34_1764 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_4 ();
 sg13g2_fill_2 FILLER_35_38 ();
 sg13g2_fill_2 FILLER_35_50 ();
 sg13g2_fill_1 FILLER_35_52 ();
 sg13g2_fill_2 FILLER_35_57 ();
 sg13g2_fill_1 FILLER_35_59 ();
 sg13g2_fill_1 FILLER_35_82 ();
 sg13g2_decap_8 FILLER_35_87 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_145 ();
 sg13g2_decap_4 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_156 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_fill_1 FILLER_35_169 ();
 sg13g2_decap_4 FILLER_35_175 ();
 sg13g2_fill_2 FILLER_35_179 ();
 sg13g2_fill_2 FILLER_35_186 ();
 sg13g2_fill_1 FILLER_35_188 ();
 sg13g2_decap_8 FILLER_35_197 ();
 sg13g2_decap_4 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_208 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_decap_4 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_243 ();
 sg13g2_decap_4 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_278 ();
 sg13g2_decap_8 FILLER_35_285 ();
 sg13g2_decap_4 FILLER_35_292 ();
 sg13g2_fill_2 FILLER_35_296 ();
 sg13g2_fill_2 FILLER_35_310 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_fill_2 FILLER_35_340 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_fill_1 FILLER_35_369 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_fill_2 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_405 ();
 sg13g2_fill_1 FILLER_35_407 ();
 sg13g2_fill_2 FILLER_35_426 ();
 sg13g2_fill_1 FILLER_35_428 ();
 sg13g2_fill_1 FILLER_35_433 ();
 sg13g2_fill_2 FILLER_35_439 ();
 sg13g2_fill_1 FILLER_35_441 ();
 sg13g2_fill_1 FILLER_35_476 ();
 sg13g2_decap_4 FILLER_35_494 ();
 sg13g2_fill_1 FILLER_35_498 ();
 sg13g2_decap_8 FILLER_35_503 ();
 sg13g2_fill_1 FILLER_35_523 ();
 sg13g2_fill_1 FILLER_35_541 ();
 sg13g2_fill_2 FILLER_35_567 ();
 sg13g2_fill_1 FILLER_35_645 ();
 sg13g2_fill_2 FILLER_35_672 ();
 sg13g2_fill_2 FILLER_35_718 ();
 sg13g2_fill_1 FILLER_35_720 ();
 sg13g2_fill_1 FILLER_35_734 ();
 sg13g2_fill_2 FILLER_35_748 ();
 sg13g2_fill_1 FILLER_35_750 ();
 sg13g2_fill_2 FILLER_35_787 ();
 sg13g2_decap_4 FILLER_35_800 ();
 sg13g2_fill_1 FILLER_35_804 ();
 sg13g2_fill_1 FILLER_35_866 ();
 sg13g2_decap_8 FILLER_35_889 ();
 sg13g2_fill_2 FILLER_35_896 ();
 sg13g2_fill_1 FILLER_35_945 ();
 sg13g2_fill_2 FILLER_35_959 ();
 sg13g2_fill_1 FILLER_35_961 ();
 sg13g2_decap_8 FILLER_35_979 ();
 sg13g2_fill_1 FILLER_35_994 ();
 sg13g2_fill_2 FILLER_35_1011 ();
 sg13g2_decap_4 FILLER_35_1021 ();
 sg13g2_fill_1 FILLER_35_1096 ();
 sg13g2_fill_2 FILLER_35_1114 ();
 sg13g2_fill_1 FILLER_35_1116 ();
 sg13g2_decap_8 FILLER_35_1183 ();
 sg13g2_fill_1 FILLER_35_1190 ();
 sg13g2_decap_8 FILLER_35_1219 ();
 sg13g2_decap_8 FILLER_35_1226 ();
 sg13g2_decap_4 FILLER_35_1233 ();
 sg13g2_fill_1 FILLER_35_1260 ();
 sg13g2_fill_1 FILLER_35_1270 ();
 sg13g2_fill_2 FILLER_35_1281 ();
 sg13g2_fill_1 FILLER_35_1283 ();
 sg13g2_decap_8 FILLER_35_1294 ();
 sg13g2_decap_4 FILLER_35_1301 ();
 sg13g2_fill_2 FILLER_35_1305 ();
 sg13g2_fill_2 FILLER_35_1317 ();
 sg13g2_fill_1 FILLER_35_1319 ();
 sg13g2_decap_8 FILLER_35_1325 ();
 sg13g2_decap_4 FILLER_35_1332 ();
 sg13g2_decap_8 FILLER_35_1352 ();
 sg13g2_decap_8 FILLER_35_1374 ();
 sg13g2_decap_4 FILLER_35_1381 ();
 sg13g2_fill_1 FILLER_35_1385 ();
 sg13g2_decap_4 FILLER_35_1399 ();
 sg13g2_fill_1 FILLER_35_1403 ();
 sg13g2_fill_2 FILLER_35_1409 ();
 sg13g2_fill_1 FILLER_35_1422 ();
 sg13g2_fill_1 FILLER_35_1444 ();
 sg13g2_fill_1 FILLER_35_1453 ();
 sg13g2_decap_8 FILLER_35_1462 ();
 sg13g2_fill_2 FILLER_35_1469 ();
 sg13g2_fill_1 FILLER_35_1471 ();
 sg13g2_decap_8 FILLER_35_1480 ();
 sg13g2_decap_8 FILLER_35_1487 ();
 sg13g2_fill_1 FILLER_35_1498 ();
 sg13g2_fill_2 FILLER_35_1509 ();
 sg13g2_decap_4 FILLER_35_1516 ();
 sg13g2_fill_2 FILLER_35_1520 ();
 sg13g2_decap_8 FILLER_35_1535 ();
 sg13g2_decap_8 FILLER_35_1542 ();
 sg13g2_decap_8 FILLER_35_1554 ();
 sg13g2_fill_1 FILLER_35_1561 ();
 sg13g2_decap_8 FILLER_35_1580 ();
 sg13g2_decap_8 FILLER_35_1587 ();
 sg13g2_decap_4 FILLER_35_1594 ();
 sg13g2_fill_1 FILLER_35_1598 ();
 sg13g2_fill_2 FILLER_35_1612 ();
 sg13g2_decap_8 FILLER_35_1622 ();
 sg13g2_fill_2 FILLER_35_1629 ();
 sg13g2_fill_1 FILLER_35_1631 ();
 sg13g2_decap_8 FILLER_35_1648 ();
 sg13g2_decap_8 FILLER_35_1673 ();
 sg13g2_fill_2 FILLER_35_1680 ();
 sg13g2_fill_2 FILLER_35_1692 ();
 sg13g2_fill_1 FILLER_35_1694 ();
 sg13g2_decap_8 FILLER_35_1709 ();
 sg13g2_decap_8 FILLER_35_1716 ();
 sg13g2_decap_4 FILLER_35_1723 ();
 sg13g2_fill_2 FILLER_35_1727 ();
 sg13g2_fill_1 FILLER_35_1741 ();
 sg13g2_decap_4 FILLER_35_1763 ();
 sg13g2_fill_1 FILLER_35_1767 ();
 sg13g2_fill_1 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_83 ();
 sg13g2_fill_1 FILLER_36_99 ();
 sg13g2_decap_4 FILLER_36_113 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_decap_4 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_fill_1 FILLER_36_177 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_207 ();
 sg13g2_decap_4 FILLER_36_214 ();
 sg13g2_fill_1 FILLER_36_218 ();
 sg13g2_fill_2 FILLER_36_237 ();
 sg13g2_fill_1 FILLER_36_239 ();
 sg13g2_decap_8 FILLER_36_271 ();
 sg13g2_fill_2 FILLER_36_294 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_decap_8 FILLER_36_328 ();
 sg13g2_decap_8 FILLER_36_335 ();
 sg13g2_decap_4 FILLER_36_342 ();
 sg13g2_fill_1 FILLER_36_352 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_fill_1 FILLER_36_378 ();
 sg13g2_decap_4 FILLER_36_397 ();
 sg13g2_fill_2 FILLER_36_401 ();
 sg13g2_decap_4 FILLER_36_431 ();
 sg13g2_fill_2 FILLER_36_435 ();
 sg13g2_fill_2 FILLER_36_456 ();
 sg13g2_decap_4 FILLER_36_468 ();
 sg13g2_fill_2 FILLER_36_472 ();
 sg13g2_decap_4 FILLER_36_489 ();
 sg13g2_decap_8 FILLER_36_508 ();
 sg13g2_fill_2 FILLER_36_515 ();
 sg13g2_decap_8 FILLER_36_530 ();
 sg13g2_fill_2 FILLER_36_537 ();
 sg13g2_fill_1 FILLER_36_552 ();
 sg13g2_decap_8 FILLER_36_570 ();
 sg13g2_decap_4 FILLER_36_577 ();
 sg13g2_fill_1 FILLER_36_581 ();
 sg13g2_fill_1 FILLER_36_585 ();
 sg13g2_decap_8 FILLER_36_603 ();
 sg13g2_decap_4 FILLER_36_610 ();
 sg13g2_fill_1 FILLER_36_614 ();
 sg13g2_decap_8 FILLER_36_666 ();
 sg13g2_decap_4 FILLER_36_673 ();
 sg13g2_fill_2 FILLER_36_677 ();
 sg13g2_fill_1 FILLER_36_683 ();
 sg13g2_fill_1 FILLER_36_694 ();
 sg13g2_fill_2 FILLER_36_699 ();
 sg13g2_fill_1 FILLER_36_701 ();
 sg13g2_decap_4 FILLER_36_711 ();
 sg13g2_decap_4 FILLER_36_752 ();
 sg13g2_fill_1 FILLER_36_756 ();
 sg13g2_fill_2 FILLER_36_805 ();
 sg13g2_fill_1 FILLER_36_813 ();
 sg13g2_fill_1 FILLER_36_828 ();
 sg13g2_fill_1 FILLER_36_887 ();
 sg13g2_fill_2 FILLER_36_918 ();
 sg13g2_fill_2 FILLER_36_952 ();
 sg13g2_fill_1 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_972 ();
 sg13g2_decap_4 FILLER_36_979 ();
 sg13g2_decap_4 FILLER_36_988 ();
 sg13g2_decap_8 FILLER_36_997 ();
 sg13g2_fill_1 FILLER_36_1004 ();
 sg13g2_fill_1 FILLER_36_1010 ();
 sg13g2_decap_8 FILLER_36_1016 ();
 sg13g2_fill_1 FILLER_36_1023 ();
 sg13g2_decap_8 FILLER_36_1028 ();
 sg13g2_fill_1 FILLER_36_1035 ();
 sg13g2_decap_8 FILLER_36_1040 ();
 sg13g2_decap_4 FILLER_36_1047 ();
 sg13g2_fill_1 FILLER_36_1051 ();
 sg13g2_decap_8 FILLER_36_1065 ();
 sg13g2_decap_4 FILLER_36_1072 ();
 sg13g2_decap_4 FILLER_36_1134 ();
 sg13g2_decap_8 FILLER_36_1201 ();
 sg13g2_decap_8 FILLER_36_1208 ();
 sg13g2_decap_4 FILLER_36_1215 ();
 sg13g2_fill_1 FILLER_36_1219 ();
 sg13g2_fill_1 FILLER_36_1239 ();
 sg13g2_fill_2 FILLER_36_1244 ();
 sg13g2_decap_8 FILLER_36_1254 ();
 sg13g2_decap_4 FILLER_36_1261 ();
 sg13g2_fill_2 FILLER_36_1277 ();
 sg13g2_fill_1 FILLER_36_1279 ();
 sg13g2_decap_8 FILLER_36_1290 ();
 sg13g2_decap_8 FILLER_36_1297 ();
 sg13g2_fill_2 FILLER_36_1304 ();
 sg13g2_fill_1 FILLER_36_1306 ();
 sg13g2_decap_8 FILLER_36_1321 ();
 sg13g2_decap_4 FILLER_36_1350 ();
 sg13g2_fill_2 FILLER_36_1354 ();
 sg13g2_fill_2 FILLER_36_1366 ();
 sg13g2_decap_8 FILLER_36_1383 ();
 sg13g2_decap_8 FILLER_36_1390 ();
 sg13g2_fill_1 FILLER_36_1397 ();
 sg13g2_decap_8 FILLER_36_1406 ();
 sg13g2_fill_2 FILLER_36_1413 ();
 sg13g2_fill_1 FILLER_36_1415 ();
 sg13g2_fill_2 FILLER_36_1434 ();
 sg13g2_decap_8 FILLER_36_1452 ();
 sg13g2_decap_8 FILLER_36_1459 ();
 sg13g2_fill_2 FILLER_36_1466 ();
 sg13g2_decap_4 FILLER_36_1486 ();
 sg13g2_fill_1 FILLER_36_1495 ();
 sg13g2_decap_4 FILLER_36_1508 ();
 sg13g2_fill_2 FILLER_36_1512 ();
 sg13g2_fill_1 FILLER_36_1523 ();
 sg13g2_fill_2 FILLER_36_1545 ();
 sg13g2_fill_1 FILLER_36_1547 ();
 sg13g2_fill_2 FILLER_36_1582 ();
 sg13g2_fill_1 FILLER_36_1584 ();
 sg13g2_decap_8 FILLER_36_1595 ();
 sg13g2_decap_8 FILLER_36_1602 ();
 sg13g2_decap_4 FILLER_36_1609 ();
 sg13g2_fill_1 FILLER_36_1613 ();
 sg13g2_decap_4 FILLER_36_1622 ();
 sg13g2_fill_1 FILLER_36_1626 ();
 sg13g2_fill_1 FILLER_36_1640 ();
 sg13g2_decap_8 FILLER_36_1653 ();
 sg13g2_fill_1 FILLER_36_1660 ();
 sg13g2_fill_2 FILLER_36_1683 ();
 sg13g2_fill_1 FILLER_36_1685 ();
 sg13g2_fill_1 FILLER_36_1691 ();
 sg13g2_decap_8 FILLER_36_1705 ();
 sg13g2_decap_4 FILLER_36_1712 ();
 sg13g2_fill_2 FILLER_36_1716 ();
 sg13g2_fill_2 FILLER_36_1729 ();
 sg13g2_fill_1 FILLER_36_1731 ();
 sg13g2_fill_2 FILLER_36_1737 ();
 sg13g2_decap_8 FILLER_36_1760 ();
 sg13g2_fill_1 FILLER_36_1767 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_7 ();
 sg13g2_fill_2 FILLER_37_37 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_decap_4 FILLER_37_50 ();
 sg13g2_fill_2 FILLER_37_118 ();
 sg13g2_decap_4 FILLER_37_148 ();
 sg13g2_decap_4 FILLER_37_170 ();
 sg13g2_decap_4 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_decap_8 FILLER_37_233 ();
 sg13g2_fill_2 FILLER_37_240 ();
 sg13g2_decap_8 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_decap_4 FILLER_37_277 ();
 sg13g2_fill_1 FILLER_37_285 ();
 sg13g2_fill_2 FILLER_37_291 ();
 sg13g2_decap_4 FILLER_37_313 ();
 sg13g2_fill_2 FILLER_37_317 ();
 sg13g2_decap_4 FILLER_37_323 ();
 sg13g2_decap_8 FILLER_37_346 ();
 sg13g2_fill_2 FILLER_37_353 ();
 sg13g2_fill_1 FILLER_37_355 ();
 sg13g2_fill_2 FILLER_37_384 ();
 sg13g2_fill_1 FILLER_37_386 ();
 sg13g2_decap_4 FILLER_37_399 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_414 ();
 sg13g2_fill_1 FILLER_37_416 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_2 FILLER_37_436 ();
 sg13g2_fill_1 FILLER_37_517 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_4 FILLER_37_570 ();
 sg13g2_fill_1 FILLER_37_574 ();
 sg13g2_fill_2 FILLER_37_592 ();
 sg13g2_fill_1 FILLER_37_594 ();
 sg13g2_fill_1 FILLER_37_599 ();
 sg13g2_fill_1 FILLER_37_611 ();
 sg13g2_fill_2 FILLER_37_659 ();
 sg13g2_fill_1 FILLER_37_661 ();
 sg13g2_decap_8 FILLER_37_716 ();
 sg13g2_fill_2 FILLER_37_723 ();
 sg13g2_fill_1 FILLER_37_738 ();
 sg13g2_fill_2 FILLER_37_757 ();
 sg13g2_decap_4 FILLER_37_781 ();
 sg13g2_fill_2 FILLER_37_785 ();
 sg13g2_fill_2 FILLER_37_802 ();
 sg13g2_fill_2 FILLER_37_829 ();
 sg13g2_fill_1 FILLER_37_831 ();
 sg13g2_decap_4 FILLER_37_845 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_fill_1 FILLER_37_910 ();
 sg13g2_fill_1 FILLER_37_928 ();
 sg13g2_decap_8 FILLER_37_947 ();
 sg13g2_fill_1 FILLER_37_954 ();
 sg13g2_fill_2 FILLER_37_978 ();
 sg13g2_fill_2 FILLER_37_1024 ();
 sg13g2_fill_1 FILLER_37_1026 ();
 sg13g2_fill_2 FILLER_37_1098 ();
 sg13g2_fill_1 FILLER_37_1100 ();
 sg13g2_fill_1 FILLER_37_1123 ();
 sg13g2_fill_2 FILLER_37_1133 ();
 sg13g2_fill_1 FILLER_37_1211 ();
 sg13g2_fill_2 FILLER_37_1234 ();
 sg13g2_fill_2 FILLER_37_1261 ();
 sg13g2_fill_2 FILLER_37_1272 ();
 sg13g2_fill_2 FILLER_37_1278 ();
 sg13g2_decap_4 FILLER_37_1294 ();
 sg13g2_fill_2 FILLER_37_1301 ();
 sg13g2_fill_2 FILLER_37_1313 ();
 sg13g2_decap_4 FILLER_37_1325 ();
 sg13g2_fill_2 FILLER_37_1329 ();
 sg13g2_decap_4 FILLER_37_1349 ();
 sg13g2_decap_8 FILLER_37_1373 ();
 sg13g2_fill_2 FILLER_37_1380 ();
 sg13g2_fill_1 FILLER_37_1382 ();
 sg13g2_fill_2 FILLER_37_1416 ();
 sg13g2_fill_1 FILLER_37_1418 ();
 sg13g2_decap_8 FILLER_37_1424 ();
 sg13g2_decap_4 FILLER_37_1459 ();
 sg13g2_fill_2 FILLER_37_1468 ();
 sg13g2_fill_1 FILLER_37_1470 ();
 sg13g2_fill_2 FILLER_37_1484 ();
 sg13g2_decap_4 FILLER_37_1518 ();
 sg13g2_fill_1 FILLER_37_1539 ();
 sg13g2_fill_2 FILLER_37_1547 ();
 sg13g2_fill_1 FILLER_37_1549 ();
 sg13g2_decap_8 FILLER_37_1555 ();
 sg13g2_fill_2 FILLER_37_1562 ();
 sg13g2_fill_1 FILLER_37_1564 ();
 sg13g2_fill_2 FILLER_37_1583 ();
 sg13g2_fill_1 FILLER_37_1585 ();
 sg13g2_decap_8 FILLER_37_1593 ();
 sg13g2_decap_4 FILLER_37_1600 ();
 sg13g2_fill_2 FILLER_37_1604 ();
 sg13g2_fill_1 FILLER_37_1614 ();
 sg13g2_fill_1 FILLER_37_1629 ();
 sg13g2_fill_2 FILLER_37_1638 ();
 sg13g2_decap_8 FILLER_37_1651 ();
 sg13g2_fill_1 FILLER_37_1658 ();
 sg13g2_fill_2 FILLER_37_1685 ();
 sg13g2_decap_4 FILLER_37_1708 ();
 sg13g2_fill_2 FILLER_37_1712 ();
 sg13g2_fill_1 FILLER_37_1726 ();
 sg13g2_fill_2 FILLER_37_1747 ();
 sg13g2_decap_8 FILLER_37_1761 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_29 ();
 sg13g2_fill_1 FILLER_38_33 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_decap_4 FILLER_38_90 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_fill_2 FILLER_38_117 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_1 FILLER_38_129 ();
 sg13g2_decap_8 FILLER_38_149 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_decap_8 FILLER_38_181 ();
 sg13g2_decap_8 FILLER_38_188 ();
 sg13g2_fill_1 FILLER_38_195 ();
 sg13g2_decap_8 FILLER_38_205 ();
 sg13g2_decap_4 FILLER_38_212 ();
 sg13g2_decap_4 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_249 ();
 sg13g2_fill_2 FILLER_38_256 ();
 sg13g2_fill_1 FILLER_38_258 ();
 sg13g2_fill_1 FILLER_38_267 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_fill_1 FILLER_38_302 ();
 sg13g2_decap_8 FILLER_38_311 ();
 sg13g2_decap_8 FILLER_38_318 ();
 sg13g2_decap_4 FILLER_38_325 ();
 sg13g2_decap_4 FILLER_38_342 ();
 sg13g2_fill_2 FILLER_38_358 ();
 sg13g2_fill_1 FILLER_38_360 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_fill_2 FILLER_38_379 ();
 sg13g2_fill_1 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_412 ();
 sg13g2_decap_4 FILLER_38_419 ();
 sg13g2_decap_4 FILLER_38_458 ();
 sg13g2_fill_1 FILLER_38_462 ();
 sg13g2_fill_2 FILLER_38_489 ();
 sg13g2_fill_1 FILLER_38_491 ();
 sg13g2_fill_1 FILLER_38_511 ();
 sg13g2_decap_4 FILLER_38_534 ();
 sg13g2_decap_8 FILLER_38_550 ();
 sg13g2_fill_1 FILLER_38_557 ();
 sg13g2_decap_8 FILLER_38_571 ();
 sg13g2_fill_1 FILLER_38_578 ();
 sg13g2_fill_1 FILLER_38_592 ();
 sg13g2_decap_4 FILLER_38_658 ();
 sg13g2_fill_1 FILLER_38_662 ();
 sg13g2_fill_1 FILLER_38_677 ();
 sg13g2_fill_1 FILLER_38_687 ();
 sg13g2_fill_1 FILLER_38_706 ();
 sg13g2_fill_1 FILLER_38_738 ();
 sg13g2_decap_8 FILLER_38_835 ();
 sg13g2_decap_4 FILLER_38_858 ();
 sg13g2_fill_1 FILLER_38_862 ();
 sg13g2_fill_1 FILLER_38_914 ();
 sg13g2_decap_4 FILLER_38_947 ();
 sg13g2_fill_2 FILLER_38_951 ();
 sg13g2_decap_8 FILLER_38_966 ();
 sg13g2_fill_2 FILLER_38_973 ();
 sg13g2_fill_1 FILLER_38_975 ();
 sg13g2_fill_2 FILLER_38_997 ();
 sg13g2_fill_1 FILLER_38_1010 ();
 sg13g2_fill_2 FILLER_38_1086 ();
 sg13g2_fill_1 FILLER_38_1088 ();
 sg13g2_decap_4 FILLER_38_1093 ();
 sg13g2_fill_2 FILLER_38_1101 ();
 sg13g2_fill_2 FILLER_38_1125 ();
 sg13g2_fill_1 FILLER_38_1127 ();
 sg13g2_decap_8 FILLER_38_1195 ();
 sg13g2_decap_8 FILLER_38_1202 ();
 sg13g2_decap_8 FILLER_38_1209 ();
 sg13g2_fill_2 FILLER_38_1216 ();
 sg13g2_fill_1 FILLER_38_1218 ();
 sg13g2_decap_8 FILLER_38_1232 ();
 sg13g2_decap_4 FILLER_38_1239 ();
 sg13g2_fill_1 FILLER_38_1243 ();
 sg13g2_decap_8 FILLER_38_1248 ();
 sg13g2_decap_8 FILLER_38_1260 ();
 sg13g2_fill_1 FILLER_38_1267 ();
 sg13g2_fill_1 FILLER_38_1278 ();
 sg13g2_decap_8 FILLER_38_1294 ();
 sg13g2_decap_4 FILLER_38_1301 ();
 sg13g2_fill_2 FILLER_38_1305 ();
 sg13g2_fill_1 FILLER_38_1347 ();
 sg13g2_fill_2 FILLER_38_1358 ();
 sg13g2_fill_1 FILLER_38_1360 ();
 sg13g2_fill_1 FILLER_38_1369 ();
 sg13g2_decap_4 FILLER_38_1378 ();
 sg13g2_fill_2 FILLER_38_1382 ();
 sg13g2_decap_8 FILLER_38_1388 ();
 sg13g2_decap_8 FILLER_38_1395 ();
 sg13g2_fill_1 FILLER_38_1402 ();
 sg13g2_decap_4 FILLER_38_1418 ();
 sg13g2_decap_4 FILLER_38_1439 ();
 sg13g2_fill_2 FILLER_38_1443 ();
 sg13g2_decap_8 FILLER_38_1455 ();
 sg13g2_decap_4 FILLER_38_1462 ();
 sg13g2_fill_1 FILLER_38_1466 ();
 sg13g2_fill_2 FILLER_38_1479 ();
 sg13g2_fill_2 FILLER_38_1485 ();
 sg13g2_fill_1 FILLER_38_1487 ();
 sg13g2_fill_2 FILLER_38_1502 ();
 sg13g2_fill_1 FILLER_38_1504 ();
 sg13g2_fill_2 FILLER_38_1531 ();
 sg13g2_fill_1 FILLER_38_1533 ();
 sg13g2_decap_8 FILLER_38_1544 ();
 sg13g2_fill_1 FILLER_38_1578 ();
 sg13g2_decap_8 FILLER_38_1591 ();
 sg13g2_decap_8 FILLER_38_1598 ();
 sg13g2_fill_2 FILLER_38_1605 ();
 sg13g2_decap_8 FILLER_38_1625 ();
 sg13g2_fill_1 FILLER_38_1635 ();
 sg13g2_decap_8 FILLER_38_1645 ();
 sg13g2_decap_4 FILLER_38_1652 ();
 sg13g2_fill_2 FILLER_38_1656 ();
 sg13g2_fill_2 FILLER_38_1666 ();
 sg13g2_fill_2 FILLER_38_1681 ();
 sg13g2_fill_1 FILLER_38_1683 ();
 sg13g2_decap_8 FILLER_38_1701 ();
 sg13g2_decap_8 FILLER_38_1708 ();
 sg13g2_decap_4 FILLER_38_1715 ();
 sg13g2_decap_4 FILLER_38_1727 ();
 sg13g2_fill_1 FILLER_38_1738 ();
 sg13g2_decap_8 FILLER_38_1754 ();
 sg13g2_decap_8 FILLER_38_1761 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_4 ();
 sg13g2_decap_4 FILLER_39_10 ();
 sg13g2_fill_1 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_44 ();
 sg13g2_decap_8 FILLER_39_55 ();
 sg13g2_fill_2 FILLER_39_89 ();
 sg13g2_fill_1 FILLER_39_100 ();
 sg13g2_decap_8 FILLER_39_114 ();
 sg13g2_fill_2 FILLER_39_121 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_fill_1 FILLER_39_146 ();
 sg13g2_fill_1 FILLER_39_156 ();
 sg13g2_fill_1 FILLER_39_175 ();
 sg13g2_decap_4 FILLER_39_188 ();
 sg13g2_fill_1 FILLER_39_254 ();
 sg13g2_decap_4 FILLER_39_273 ();
 sg13g2_fill_2 FILLER_39_277 ();
 sg13g2_fill_1 FILLER_39_295 ();
 sg13g2_fill_1 FILLER_39_322 ();
 sg13g2_fill_2 FILLER_39_336 ();
 sg13g2_fill_1 FILLER_39_338 ();
 sg13g2_decap_4 FILLER_39_344 ();
 sg13g2_fill_2 FILLER_39_348 ();
 sg13g2_fill_1 FILLER_39_358 ();
 sg13g2_decap_4 FILLER_39_364 ();
 sg13g2_fill_1 FILLER_39_368 ();
 sg13g2_fill_2 FILLER_39_373 ();
 sg13g2_fill_2 FILLER_39_388 ();
 sg13g2_fill_1 FILLER_39_390 ();
 sg13g2_decap_4 FILLER_39_415 ();
 sg13g2_decap_4 FILLER_39_432 ();
 sg13g2_fill_2 FILLER_39_444 ();
 sg13g2_decap_8 FILLER_39_477 ();
 sg13g2_decap_4 FILLER_39_484 ();
 sg13g2_fill_2 FILLER_39_488 ();
 sg13g2_fill_1 FILLER_39_550 ();
 sg13g2_fill_1 FILLER_39_612 ();
 sg13g2_fill_2 FILLER_39_640 ();
 sg13g2_fill_1 FILLER_39_642 ();
 sg13g2_decap_4 FILLER_39_724 ();
 sg13g2_fill_2 FILLER_39_741 ();
 sg13g2_fill_1 FILLER_39_753 ();
 sg13g2_fill_1 FILLER_39_763 ();
 sg13g2_fill_1 FILLER_39_786 ();
 sg13g2_decap_4 FILLER_39_793 ();
 sg13g2_fill_1 FILLER_39_813 ();
 sg13g2_decap_4 FILLER_39_875 ();
 sg13g2_decap_8 FILLER_39_928 ();
 sg13g2_decap_8 FILLER_39_935 ();
 sg13g2_decap_4 FILLER_39_942 ();
 sg13g2_fill_1 FILLER_39_946 ();
 sg13g2_decap_8 FILLER_39_968 ();
 sg13g2_decap_8 FILLER_39_975 ();
 sg13g2_fill_1 FILLER_39_982 ();
 sg13g2_decap_4 FILLER_39_991 ();
 sg13g2_fill_2 FILLER_39_1058 ();
 sg13g2_fill_2 FILLER_39_1145 ();
 sg13g2_fill_1 FILLER_39_1147 ();
 sg13g2_fill_2 FILLER_39_1184 ();
 sg13g2_fill_1 FILLER_39_1186 ();
 sg13g2_decap_4 FILLER_39_1256 ();
 sg13g2_fill_1 FILLER_39_1273 ();
 sg13g2_fill_2 FILLER_39_1289 ();
 sg13g2_decap_8 FILLER_39_1301 ();
 sg13g2_decap_8 FILLER_39_1308 ();
 sg13g2_decap_8 FILLER_39_1315 ();
 sg13g2_fill_2 FILLER_39_1322 ();
 sg13g2_fill_1 FILLER_39_1324 ();
 sg13g2_decap_8 FILLER_39_1342 ();
 sg13g2_decap_8 FILLER_39_1349 ();
 sg13g2_fill_1 FILLER_39_1356 ();
 sg13g2_fill_1 FILLER_39_1366 ();
 sg13g2_fill_1 FILLER_39_1372 ();
 sg13g2_fill_2 FILLER_39_1381 ();
 sg13g2_decap_4 FILLER_39_1400 ();
 sg13g2_fill_2 FILLER_39_1404 ();
 sg13g2_fill_1 FILLER_39_1415 ();
 sg13g2_decap_8 FILLER_39_1424 ();
 sg13g2_fill_1 FILLER_39_1431 ();
 sg13g2_decap_8 FILLER_39_1460 ();
 sg13g2_decap_4 FILLER_39_1467 ();
 sg13g2_fill_2 FILLER_39_1471 ();
 sg13g2_decap_8 FILLER_39_1502 ();
 sg13g2_decap_8 FILLER_39_1509 ();
 sg13g2_decap_8 FILLER_39_1516 ();
 sg13g2_decap_8 FILLER_39_1547 ();
 sg13g2_decap_8 FILLER_39_1554 ();
 sg13g2_decap_4 FILLER_39_1561 ();
 sg13g2_fill_2 FILLER_39_1565 ();
 sg13g2_fill_1 FILLER_39_1591 ();
 sg13g2_decap_8 FILLER_39_1600 ();
 sg13g2_fill_2 FILLER_39_1607 ();
 sg13g2_fill_2 FILLER_39_1628 ();
 sg13g2_decap_8 FILLER_39_1648 ();
 sg13g2_decap_8 FILLER_39_1655 ();
 sg13g2_decap_4 FILLER_39_1662 ();
 sg13g2_fill_1 FILLER_39_1678 ();
 sg13g2_fill_2 FILLER_39_1689 ();
 sg13g2_decap_8 FILLER_39_1706 ();
 sg13g2_decap_8 FILLER_39_1713 ();
 sg13g2_decap_8 FILLER_39_1725 ();
 sg13g2_fill_2 FILLER_39_1736 ();
 sg13g2_fill_1 FILLER_39_1738 ();
 sg13g2_decap_8 FILLER_39_1754 ();
 sg13g2_decap_8 FILLER_39_1761 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_29 ();
 sg13g2_fill_1 FILLER_40_36 ();
 sg13g2_fill_1 FILLER_40_51 ();
 sg13g2_fill_1 FILLER_40_75 ();
 sg13g2_decap_4 FILLER_40_113 ();
 sg13g2_fill_2 FILLER_40_117 ();
 sg13g2_decap_4 FILLER_40_146 ();
 sg13g2_fill_1 FILLER_40_160 ();
 sg13g2_fill_2 FILLER_40_183 ();
 sg13g2_decap_8 FILLER_40_195 ();
 sg13g2_decap_8 FILLER_40_202 ();
 sg13g2_decap_4 FILLER_40_209 ();
 sg13g2_fill_1 FILLER_40_213 ();
 sg13g2_fill_1 FILLER_40_218 ();
 sg13g2_decap_8 FILLER_40_223 ();
 sg13g2_decap_4 FILLER_40_230 ();
 sg13g2_fill_2 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_275 ();
 sg13g2_decap_4 FILLER_40_282 ();
 sg13g2_fill_1 FILLER_40_286 ();
 sg13g2_fill_1 FILLER_40_305 ();
 sg13g2_decap_4 FILLER_40_314 ();
 sg13g2_fill_1 FILLER_40_318 ();
 sg13g2_decap_4 FILLER_40_323 ();
 sg13g2_fill_1 FILLER_40_327 ();
 sg13g2_fill_2 FILLER_40_332 ();
 sg13g2_decap_4 FILLER_40_339 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_389 ();
 sg13g2_fill_1 FILLER_40_401 ();
 sg13g2_fill_1 FILLER_40_415 ();
 sg13g2_fill_2 FILLER_40_421 ();
 sg13g2_fill_1 FILLER_40_423 ();
 sg13g2_decap_8 FILLER_40_428 ();
 sg13g2_fill_2 FILLER_40_448 ();
 sg13g2_fill_1 FILLER_40_450 ();
 sg13g2_decap_8 FILLER_40_479 ();
 sg13g2_decap_8 FILLER_40_486 ();
 sg13g2_fill_1 FILLER_40_493 ();
 sg13g2_decap_8 FILLER_40_523 ();
 sg13g2_decap_8 FILLER_40_530 ();
 sg13g2_decap_8 FILLER_40_537 ();
 sg13g2_fill_1 FILLER_40_544 ();
 sg13g2_decap_8 FILLER_40_569 ();
 sg13g2_decap_4 FILLER_40_576 ();
 sg13g2_decap_4 FILLER_40_585 ();
 sg13g2_fill_2 FILLER_40_589 ();
 sg13g2_fill_1 FILLER_40_654 ();
 sg13g2_fill_2 FILLER_40_676 ();
 sg13g2_fill_1 FILLER_40_678 ();
 sg13g2_decap_4 FILLER_40_698 ();
 sg13g2_fill_1 FILLER_40_736 ();
 sg13g2_fill_1 FILLER_40_755 ();
 sg13g2_fill_1 FILLER_40_783 ();
 sg13g2_fill_2 FILLER_40_806 ();
 sg13g2_fill_2 FILLER_40_826 ();
 sg13g2_fill_1 FILLER_40_828 ();
 sg13g2_fill_2 FILLER_40_841 ();
 sg13g2_fill_2 FILLER_40_898 ();
 sg13g2_fill_1 FILLER_40_900 ();
 sg13g2_decap_8 FILLER_40_931 ();
 sg13g2_decap_4 FILLER_40_938 ();
 sg13g2_decap_8 FILLER_40_969 ();
 sg13g2_decap_8 FILLER_40_976 ();
 sg13g2_fill_2 FILLER_40_997 ();
 sg13g2_fill_1 FILLER_40_999 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_fill_1 FILLER_40_1022 ();
 sg13g2_fill_2 FILLER_40_1027 ();
 sg13g2_decap_8 FILLER_40_1046 ();
 sg13g2_decap_4 FILLER_40_1053 ();
 sg13g2_fill_2 FILLER_40_1057 ();
 sg13g2_fill_1 FILLER_40_1068 ();
 sg13g2_decap_8 FILLER_40_1073 ();
 sg13g2_decap_8 FILLER_40_1080 ();
 sg13g2_fill_2 FILLER_40_1100 ();
 sg13g2_fill_1 FILLER_40_1102 ();
 sg13g2_decap_8 FILLER_40_1161 ();
 sg13g2_fill_2 FILLER_40_1168 ();
 sg13g2_fill_1 FILLER_40_1170 ();
 sg13g2_fill_2 FILLER_40_1179 ();
 sg13g2_fill_1 FILLER_40_1181 ();
 sg13g2_fill_1 FILLER_40_1190 ();
 sg13g2_decap_8 FILLER_40_1204 ();
 sg13g2_decap_8 FILLER_40_1211 ();
 sg13g2_fill_2 FILLER_40_1218 ();
 sg13g2_fill_1 FILLER_40_1220 ();
 sg13g2_fill_2 FILLER_40_1236 ();
 sg13g2_fill_1 FILLER_40_1238 ();
 sg13g2_fill_1 FILLER_40_1272 ();
 sg13g2_decap_8 FILLER_40_1282 ();
 sg13g2_decap_4 FILLER_40_1289 ();
 sg13g2_decap_4 FILLER_40_1313 ();
 sg13g2_fill_1 FILLER_40_1317 ();
 sg13g2_fill_2 FILLER_40_1336 ();
 sg13g2_decap_4 FILLER_40_1346 ();
 sg13g2_fill_1 FILLER_40_1350 ();
 sg13g2_decap_4 FILLER_40_1361 ();
 sg13g2_fill_2 FILLER_40_1369 ();
 sg13g2_fill_1 FILLER_40_1371 ();
 sg13g2_fill_2 FILLER_40_1380 ();
 sg13g2_decap_8 FILLER_40_1387 ();
 sg13g2_decap_4 FILLER_40_1394 ();
 sg13g2_fill_2 FILLER_40_1398 ();
 sg13g2_fill_2 FILLER_40_1432 ();
 sg13g2_fill_1 FILLER_40_1434 ();
 sg13g2_fill_2 FILLER_40_1447 ();
 sg13g2_fill_1 FILLER_40_1449 ();
 sg13g2_decap_8 FILLER_40_1466 ();
 sg13g2_decap_4 FILLER_40_1473 ();
 sg13g2_decap_4 FILLER_40_1498 ();
 sg13g2_fill_1 FILLER_40_1502 ();
 sg13g2_decap_8 FILLER_40_1507 ();
 sg13g2_fill_1 FILLER_40_1514 ();
 sg13g2_fill_2 FILLER_40_1518 ();
 sg13g2_fill_2 FILLER_40_1525 ();
 sg13g2_fill_1 FILLER_40_1527 ();
 sg13g2_fill_2 FILLER_40_1554 ();
 sg13g2_fill_1 FILLER_40_1556 ();
 sg13g2_fill_2 FILLER_40_1564 ();
 sg13g2_decap_4 FILLER_40_1576 ();
 sg13g2_fill_2 FILLER_40_1580 ();
 sg13g2_decap_8 FILLER_40_1586 ();
 sg13g2_fill_2 FILLER_40_1597 ();
 sg13g2_fill_1 FILLER_40_1599 ();
 sg13g2_decap_4 FILLER_40_1612 ();
 sg13g2_decap_8 FILLER_40_1621 ();
 sg13g2_decap_8 FILLER_40_1628 ();
 sg13g2_fill_1 FILLER_40_1635 ();
 sg13g2_decap_8 FILLER_40_1646 ();
 sg13g2_decap_4 FILLER_40_1653 ();
 sg13g2_fill_1 FILLER_40_1657 ();
 sg13g2_decap_8 FILLER_40_1667 ();
 sg13g2_fill_1 FILLER_40_1684 ();
 sg13g2_decap_8 FILLER_40_1709 ();
 sg13g2_decap_8 FILLER_40_1716 ();
 sg13g2_decap_8 FILLER_40_1723 ();
 sg13g2_fill_2 FILLER_40_1730 ();
 sg13g2_decap_4 FILLER_40_1735 ();
 sg13g2_decap_8 FILLER_40_1760 ();
 sg13g2_fill_1 FILLER_40_1767 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_11 ();
 sg13g2_decap_4 FILLER_41_18 ();
 sg13g2_decap_4 FILLER_41_54 ();
 sg13g2_fill_1 FILLER_41_58 ();
 sg13g2_decap_8 FILLER_41_73 ();
 sg13g2_decap_8 FILLER_41_80 ();
 sg13g2_fill_2 FILLER_41_87 ();
 sg13g2_fill_1 FILLER_41_99 ();
 sg13g2_fill_2 FILLER_41_132 ();
 sg13g2_fill_1 FILLER_41_134 ();
 sg13g2_decap_4 FILLER_41_161 ();
 sg13g2_fill_2 FILLER_41_170 ();
 sg13g2_decap_4 FILLER_41_185 ();
 sg13g2_fill_2 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_205 ();
 sg13g2_fill_1 FILLER_41_212 ();
 sg13g2_fill_2 FILLER_41_252 ();
 sg13g2_fill_2 FILLER_41_308 ();
 sg13g2_decap_4 FILLER_41_330 ();
 sg13g2_fill_1 FILLER_41_334 ();
 sg13g2_fill_2 FILLER_41_348 ();
 sg13g2_fill_1 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_358 ();
 sg13g2_decap_8 FILLER_41_365 ();
 sg13g2_decap_4 FILLER_41_372 ();
 sg13g2_fill_1 FILLER_41_376 ();
 sg13g2_fill_2 FILLER_41_471 ();
 sg13g2_fill_1 FILLER_41_473 ();
 sg13g2_fill_2 FILLER_41_483 ();
 sg13g2_fill_1 FILLER_41_499 ();
 sg13g2_fill_2 FILLER_41_505 ();
 sg13g2_fill_1 FILLER_41_507 ();
 sg13g2_decap_4 FILLER_41_531 ();
 sg13g2_fill_2 FILLER_41_535 ();
 sg13g2_decap_4 FILLER_41_541 ();
 sg13g2_fill_2 FILLER_41_545 ();
 sg13g2_fill_2 FILLER_41_615 ();
 sg13g2_fill_1 FILLER_41_617 ();
 sg13g2_fill_1 FILLER_41_658 ();
 sg13g2_fill_1 FILLER_41_668 ();
 sg13g2_decap_8 FILLER_41_683 ();
 sg13g2_fill_1 FILLER_41_690 ();
 sg13g2_decap_8 FILLER_41_704 ();
 sg13g2_fill_2 FILLER_41_732 ();
 sg13g2_fill_2 FILLER_41_747 ();
 sg13g2_fill_1 FILLER_41_749 ();
 sg13g2_decap_4 FILLER_41_777 ();
 sg13g2_fill_1 FILLER_41_781 ();
 sg13g2_fill_2 FILLER_41_785 ();
 sg13g2_fill_2 FILLER_41_808 ();
 sg13g2_fill_1 FILLER_41_840 ();
 sg13g2_decap_4 FILLER_41_863 ();
 sg13g2_decap_4 FILLER_41_905 ();
 sg13g2_fill_2 FILLER_41_909 ();
 sg13g2_decap_4 FILLER_41_932 ();
 sg13g2_fill_2 FILLER_41_936 ();
 sg13g2_decap_4 FILLER_41_947 ();
 sg13g2_fill_1 FILLER_41_951 ();
 sg13g2_fill_1 FILLER_41_959 ();
 sg13g2_fill_1 FILLER_41_1010 ();
 sg13g2_fill_2 FILLER_41_1150 ();
 sg13g2_fill_1 FILLER_41_1216 ();
 sg13g2_decap_8 FILLER_41_1251 ();
 sg13g2_decap_8 FILLER_41_1258 ();
 sg13g2_decap_4 FILLER_41_1265 ();
 sg13g2_fill_1 FILLER_41_1269 ();
 sg13g2_decap_8 FILLER_41_1289 ();
 sg13g2_fill_1 FILLER_41_1296 ();
 sg13g2_fill_2 FILLER_41_1331 ();
 sg13g2_fill_1 FILLER_41_1333 ();
 sg13g2_decap_8 FILLER_41_1390 ();
 sg13g2_decap_8 FILLER_41_1397 ();
 sg13g2_decap_4 FILLER_41_1404 ();
 sg13g2_fill_1 FILLER_41_1418 ();
 sg13g2_decap_8 FILLER_41_1423 ();
 sg13g2_fill_2 FILLER_41_1430 ();
 sg13g2_fill_1 FILLER_41_1432 ();
 sg13g2_fill_2 FILLER_41_1441 ();
 sg13g2_fill_1 FILLER_41_1443 ();
 sg13g2_fill_1 FILLER_41_1449 ();
 sg13g2_fill_2 FILLER_41_1458 ();
 sg13g2_fill_1 FILLER_41_1460 ();
 sg13g2_decap_8 FILLER_41_1485 ();
 sg13g2_fill_2 FILLER_41_1492 ();
 sg13g2_decap_8 FILLER_41_1525 ();
 sg13g2_decap_8 FILLER_41_1532 ();
 sg13g2_fill_2 FILLER_41_1539 ();
 sg13g2_decap_8 FILLER_41_1557 ();
 sg13g2_decap_8 FILLER_41_1564 ();
 sg13g2_decap_4 FILLER_41_1571 ();
 sg13g2_decap_4 FILLER_41_1590 ();
 sg13g2_fill_1 FILLER_41_1604 ();
 sg13g2_decap_8 FILLER_41_1621 ();
 sg13g2_fill_2 FILLER_41_1628 ();
 sg13g2_fill_2 FILLER_41_1634 ();
 sg13g2_fill_2 FILLER_41_1651 ();
 sg13g2_fill_1 FILLER_41_1653 ();
 sg13g2_decap_4 FILLER_41_1675 ();
 sg13g2_decap_4 FILLER_41_1687 ();
 sg13g2_fill_1 FILLER_41_1691 ();
 sg13g2_decap_4 FILLER_41_1703 ();
 sg13g2_decap_8 FILLER_41_1717 ();
 sg13g2_fill_1 FILLER_41_1724 ();
 sg13g2_decap_8 FILLER_41_1742 ();
 sg13g2_decap_8 FILLER_41_1756 ();
 sg13g2_decap_4 FILLER_41_1763 ();
 sg13g2_fill_1 FILLER_41_1767 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_2 ();
 sg13g2_fill_2 FILLER_42_62 ();
 sg13g2_decap_8 FILLER_42_113 ();
 sg13g2_decap_8 FILLER_42_120 ();
 sg13g2_decap_8 FILLER_42_127 ();
 sg13g2_decap_8 FILLER_42_134 ();
 sg13g2_decap_8 FILLER_42_169 ();
 sg13g2_decap_8 FILLER_42_176 ();
 sg13g2_fill_2 FILLER_42_183 ();
 sg13g2_fill_1 FILLER_42_185 ();
 sg13g2_decap_4 FILLER_42_191 ();
 sg13g2_fill_1 FILLER_42_195 ();
 sg13g2_fill_1 FILLER_42_224 ();
 sg13g2_decap_4 FILLER_42_229 ();
 sg13g2_fill_1 FILLER_42_237 ();
 sg13g2_decap_4 FILLER_42_242 ();
 sg13g2_fill_2 FILLER_42_267 ();
 sg13g2_fill_2 FILLER_42_273 ();
 sg13g2_fill_2 FILLER_42_284 ();
 sg13g2_fill_1 FILLER_42_286 ();
 sg13g2_fill_1 FILLER_42_300 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_fill_2 FILLER_42_329 ();
 sg13g2_fill_1 FILLER_42_331 ();
 sg13g2_decap_4 FILLER_42_360 ();
 sg13g2_decap_8 FILLER_42_368 ();
 sg13g2_fill_2 FILLER_42_375 ();
 sg13g2_fill_1 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_390 ();
 sg13g2_decap_8 FILLER_42_397 ();
 sg13g2_decap_4 FILLER_42_404 ();
 sg13g2_fill_1 FILLER_42_408 ();
 sg13g2_decap_4 FILLER_42_414 ();
 sg13g2_decap_8 FILLER_42_422 ();
 sg13g2_decap_4 FILLER_42_429 ();
 sg13g2_fill_2 FILLER_42_433 ();
 sg13g2_fill_2 FILLER_42_463 ();
 sg13g2_decap_4 FILLER_42_560 ();
 sg13g2_fill_2 FILLER_42_564 ();
 sg13g2_fill_1 FILLER_42_592 ();
 sg13g2_fill_2 FILLER_42_627 ();
 sg13g2_fill_1 FILLER_42_629 ();
 sg13g2_fill_1 FILLER_42_635 ();
 sg13g2_decap_8 FILLER_42_703 ();
 sg13g2_fill_1 FILLER_42_710 ();
 sg13g2_fill_2 FILLER_42_735 ();
 sg13g2_fill_2 FILLER_42_759 ();
 sg13g2_decap_4 FILLER_42_791 ();
 sg13g2_fill_2 FILLER_42_798 ();
 sg13g2_fill_1 FILLER_42_800 ();
 sg13g2_fill_2 FILLER_42_872 ();
 sg13g2_decap_8 FILLER_42_878 ();
 sg13g2_decap_8 FILLER_42_898 ();
 sg13g2_fill_2 FILLER_42_905 ();
 sg13g2_fill_1 FILLER_42_907 ();
 sg13g2_decap_8 FILLER_42_952 ();
 sg13g2_fill_2 FILLER_42_999 ();
 sg13g2_decap_8 FILLER_42_1007 ();
 sg13g2_fill_2 FILLER_42_1014 ();
 sg13g2_fill_1 FILLER_42_1016 ();
 sg13g2_fill_1 FILLER_42_1021 ();
 sg13g2_decap_8 FILLER_42_1027 ();
 sg13g2_decap_4 FILLER_42_1034 ();
 sg13g2_fill_1 FILLER_42_1055 ();
 sg13g2_decap_8 FILLER_42_1074 ();
 sg13g2_fill_1 FILLER_42_1081 ();
 sg13g2_decap_4 FILLER_42_1110 ();
 sg13g2_fill_2 FILLER_42_1128 ();
 sg13g2_fill_1 FILLER_42_1156 ();
 sg13g2_fill_2 FILLER_42_1170 ();
 sg13g2_fill_2 FILLER_42_1177 ();
 sg13g2_fill_2 FILLER_42_1201 ();
 sg13g2_fill_1 FILLER_42_1203 ();
 sg13g2_decap_8 FILLER_42_1235 ();
 sg13g2_decap_8 FILLER_42_1242 ();
 sg13g2_fill_2 FILLER_42_1249 ();
 sg13g2_fill_1 FILLER_42_1251 ();
 sg13g2_decap_8 FILLER_42_1300 ();
 sg13g2_fill_2 FILLER_42_1307 ();
 sg13g2_decap_4 FILLER_42_1314 ();
 sg13g2_decap_8 FILLER_42_1328 ();
 sg13g2_fill_2 FILLER_42_1335 ();
 sg13g2_decap_8 FILLER_42_1351 ();
 sg13g2_decap_8 FILLER_42_1358 ();
 sg13g2_decap_4 FILLER_42_1365 ();
 sg13g2_fill_2 FILLER_42_1369 ();
 sg13g2_decap_8 FILLER_42_1377 ();
 sg13g2_decap_8 FILLER_42_1388 ();
 sg13g2_decap_4 FILLER_42_1395 ();
 sg13g2_decap_8 FILLER_42_1431 ();
 sg13g2_decap_8 FILLER_42_1456 ();
 sg13g2_decap_8 FILLER_42_1463 ();
 sg13g2_decap_8 FILLER_42_1470 ();
 sg13g2_fill_2 FILLER_42_1477 ();
 sg13g2_fill_1 FILLER_42_1492 ();
 sg13g2_decap_8 FILLER_42_1514 ();
 sg13g2_decap_4 FILLER_42_1521 ();
 sg13g2_fill_1 FILLER_42_1525 ();
 sg13g2_fill_1 FILLER_42_1531 ();
 sg13g2_fill_1 FILLER_42_1544 ();
 sg13g2_decap_4 FILLER_42_1550 ();
 sg13g2_decap_8 FILLER_42_1572 ();
 sg13g2_fill_2 FILLER_42_1579 ();
 sg13g2_fill_1 FILLER_42_1581 ();
 sg13g2_fill_2 FILLER_42_1591 ();
 sg13g2_decap_8 FILLER_42_1612 ();
 sg13g2_decap_4 FILLER_42_1619 ();
 sg13g2_fill_1 FILLER_42_1623 ();
 sg13g2_decap_8 FILLER_42_1665 ();
 sg13g2_decap_4 FILLER_42_1672 ();
 sg13g2_fill_1 FILLER_42_1676 ();
 sg13g2_decap_8 FILLER_42_1686 ();
 sg13g2_decap_4 FILLER_42_1693 ();
 sg13g2_fill_2 FILLER_42_1697 ();
 sg13g2_fill_1 FILLER_42_1723 ();
 sg13g2_fill_2 FILLER_42_1748 ();
 sg13g2_fill_1 FILLER_42_1750 ();
 sg13g2_decap_4 FILLER_42_1764 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_7 ();
 sg13g2_decap_4 FILLER_43_12 ();
 sg13g2_fill_1 FILLER_43_16 ();
 sg13g2_fill_1 FILLER_43_44 ();
 sg13g2_decap_4 FILLER_43_58 ();
 sg13g2_fill_1 FILLER_43_76 ();
 sg13g2_fill_1 FILLER_43_93 ();
 sg13g2_fill_2 FILLER_43_100 ();
 sg13g2_fill_2 FILLER_43_130 ();
 sg13g2_decap_8 FILLER_43_136 ();
 sg13g2_decap_8 FILLER_43_143 ();
 sg13g2_decap_4 FILLER_43_150 ();
 sg13g2_fill_2 FILLER_43_154 ();
 sg13g2_fill_1 FILLER_43_179 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_decap_8 FILLER_43_215 ();
 sg13g2_decap_4 FILLER_43_222 ();
 sg13g2_fill_2 FILLER_43_226 ();
 sg13g2_fill_2 FILLER_43_270 ();
 sg13g2_fill_1 FILLER_43_320 ();
 sg13g2_decap_4 FILLER_43_353 ();
 sg13g2_fill_2 FILLER_43_357 ();
 sg13g2_decap_4 FILLER_43_392 ();
 sg13g2_decap_4 FILLER_43_400 ();
 sg13g2_fill_1 FILLER_43_404 ();
 sg13g2_fill_1 FILLER_43_418 ();
 sg13g2_fill_2 FILLER_43_446 ();
 sg13g2_fill_2 FILLER_43_456 ();
 sg13g2_fill_1 FILLER_43_458 ();
 sg13g2_fill_1 FILLER_43_469 ();
 sg13g2_fill_2 FILLER_43_492 ();
 sg13g2_fill_1 FILLER_43_494 ();
 sg13g2_fill_1 FILLER_43_515 ();
 sg13g2_fill_2 FILLER_43_521 ();
 sg13g2_decap_8 FILLER_43_527 ();
 sg13g2_fill_1 FILLER_43_534 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_4 FILLER_43_553 ();
 sg13g2_fill_2 FILLER_43_557 ();
 sg13g2_fill_1 FILLER_43_629 ();
 sg13g2_fill_2 FILLER_43_641 ();
 sg13g2_fill_1 FILLER_43_643 ();
 sg13g2_decap_8 FILLER_43_661 ();
 sg13g2_fill_2 FILLER_43_668 ();
 sg13g2_fill_1 FILLER_43_670 ();
 sg13g2_fill_2 FILLER_43_730 ();
 sg13g2_fill_1 FILLER_43_767 ();
 sg13g2_fill_2 FILLER_43_862 ();
 sg13g2_fill_2 FILLER_43_878 ();
 sg13g2_fill_1 FILLER_43_889 ();
 sg13g2_fill_1 FILLER_43_917 ();
 sg13g2_fill_2 FILLER_43_936 ();
 sg13g2_fill_2 FILLER_43_965 ();
 sg13g2_decap_4 FILLER_43_977 ();
 sg13g2_fill_1 FILLER_43_1020 ();
 sg13g2_decap_8 FILLER_43_1030 ();
 sg13g2_fill_2 FILLER_43_1070 ();
 sg13g2_fill_1 FILLER_43_1127 ();
 sg13g2_decap_4 FILLER_43_1164 ();
 sg13g2_fill_2 FILLER_43_1210 ();
 sg13g2_fill_1 FILLER_43_1212 ();
 sg13g2_fill_2 FILLER_43_1239 ();
 sg13g2_fill_1 FILLER_43_1241 ();
 sg13g2_fill_2 FILLER_43_1246 ();
 sg13g2_decap_8 FILLER_43_1260 ();
 sg13g2_decap_4 FILLER_43_1267 ();
 sg13g2_fill_2 FILLER_43_1278 ();
 sg13g2_fill_2 FILLER_43_1294 ();
 sg13g2_fill_2 FILLER_43_1328 ();
 sg13g2_fill_2 FILLER_43_1344 ();
 sg13g2_decap_4 FILLER_43_1354 ();
 sg13g2_fill_2 FILLER_43_1358 ();
 sg13g2_fill_2 FILLER_43_1372 ();
 sg13g2_decap_8 FILLER_43_1387 ();
 sg13g2_decap_4 FILLER_43_1394 ();
 sg13g2_fill_2 FILLER_43_1398 ();
 sg13g2_decap_8 FILLER_43_1408 ();
 sg13g2_decap_8 FILLER_43_1415 ();
 sg13g2_decap_8 FILLER_43_1422 ();
 sg13g2_fill_2 FILLER_43_1429 ();
 sg13g2_fill_1 FILLER_43_1431 ();
 sg13g2_decap_8 FILLER_43_1458 ();
 sg13g2_decap_4 FILLER_43_1465 ();
 sg13g2_fill_1 FILLER_43_1469 ();
 sg13g2_decap_4 FILLER_43_1483 ();
 sg13g2_fill_1 FILLER_43_1487 ();
 sg13g2_fill_2 FILLER_43_1506 ();
 sg13g2_fill_1 FILLER_43_1508 ();
 sg13g2_fill_2 FILLER_43_1514 ();
 sg13g2_decap_4 FILLER_43_1535 ();
 sg13g2_fill_1 FILLER_43_1539 ();
 sg13g2_fill_2 FILLER_43_1553 ();
 sg13g2_fill_1 FILLER_43_1555 ();
 sg13g2_decap_4 FILLER_43_1572 ();
 sg13g2_fill_2 FILLER_43_1576 ();
 sg13g2_fill_1 FILLER_43_1595 ();
 sg13g2_fill_2 FILLER_43_1606 ();
 sg13g2_decap_8 FILLER_43_1616 ();
 sg13g2_decap_4 FILLER_43_1623 ();
 sg13g2_fill_1 FILLER_43_1627 ();
 sg13g2_fill_2 FILLER_43_1631 ();
 sg13g2_fill_1 FILLER_43_1638 ();
 sg13g2_decap_8 FILLER_43_1650 ();
 sg13g2_fill_1 FILLER_43_1657 ();
 sg13g2_decap_4 FILLER_43_1667 ();
 sg13g2_fill_2 FILLER_43_1671 ();
 sg13g2_decap_8 FILLER_43_1693 ();
 sg13g2_fill_1 FILLER_43_1700 ();
 sg13g2_decap_4 FILLER_43_1726 ();
 sg13g2_fill_1 FILLER_43_1730 ();
 sg13g2_decap_4 FILLER_43_1747 ();
 sg13g2_fill_2 FILLER_43_1751 ();
 sg13g2_decap_8 FILLER_43_1758 ();
 sg13g2_fill_2 FILLER_43_1765 ();
 sg13g2_fill_1 FILLER_43_1767 ();
 sg13g2_decap_4 FILLER_44_0 ();
 sg13g2_fill_1 FILLER_44_32 ();
 sg13g2_fill_2 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_57 ();
 sg13g2_decap_8 FILLER_44_112 ();
 sg13g2_decap_4 FILLER_44_119 ();
 sg13g2_fill_1 FILLER_44_154 ();
 sg13g2_decap_8 FILLER_44_245 ();
 sg13g2_fill_2 FILLER_44_252 ();
 sg13g2_fill_2 FILLER_44_274 ();
 sg13g2_fill_1 FILLER_44_276 ();
 sg13g2_fill_2 FILLER_44_281 ();
 sg13g2_fill_1 FILLER_44_296 ();
 sg13g2_decap_4 FILLER_44_315 ();
 sg13g2_fill_2 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_371 ();
 sg13g2_fill_1 FILLER_44_390 ();
 sg13g2_decap_4 FILLER_44_418 ();
 sg13g2_fill_2 FILLER_44_422 ();
 sg13g2_decap_8 FILLER_44_428 ();
 sg13g2_decap_4 FILLER_44_435 ();
 sg13g2_fill_1 FILLER_44_462 ();
 sg13g2_fill_2 FILLER_44_476 ();
 sg13g2_fill_1 FILLER_44_514 ();
 sg13g2_fill_2 FILLER_44_527 ();
 sg13g2_fill_1 FILLER_44_529 ();
 sg13g2_decap_4 FILLER_44_558 ();
 sg13g2_fill_2 FILLER_44_562 ();
 sg13g2_fill_1 FILLER_44_568 ();
 sg13g2_fill_2 FILLER_44_582 ();
 sg13g2_fill_2 FILLER_44_610 ();
 sg13g2_decap_4 FILLER_44_621 ();
 sg13g2_fill_2 FILLER_44_643 ();
 sg13g2_fill_1 FILLER_44_712 ();
 sg13g2_fill_2 FILLER_44_722 ();
 sg13g2_fill_1 FILLER_44_724 ();
 sg13g2_decap_8 FILLER_44_762 ();
 sg13g2_decap_8 FILLER_44_769 ();
 sg13g2_decap_8 FILLER_44_776 ();
 sg13g2_fill_1 FILLER_44_783 ();
 sg13g2_fill_1 FILLER_44_800 ();
 sg13g2_fill_2 FILLER_44_819 ();
 sg13g2_fill_2 FILLER_44_825 ();
 sg13g2_fill_1 FILLER_44_827 ();
 sg13g2_fill_2 FILLER_44_931 ();
 sg13g2_fill_1 FILLER_44_942 ();
 sg13g2_decap_8 FILLER_44_956 ();
 sg13g2_decap_4 FILLER_44_963 ();
 sg13g2_decap_8 FILLER_44_1004 ();
 sg13g2_decap_4 FILLER_44_1011 ();
 sg13g2_fill_2 FILLER_44_1015 ();
 sg13g2_fill_2 FILLER_44_1045 ();
 sg13g2_fill_1 FILLER_44_1047 ();
 sg13g2_fill_2 FILLER_44_1125 ();
 sg13g2_fill_2 FILLER_44_1201 ();
 sg13g2_fill_1 FILLER_44_1203 ();
 sg13g2_fill_2 FILLER_44_1237 ();
 sg13g2_fill_1 FILLER_44_1239 ();
 sg13g2_fill_1 FILLER_44_1264 ();
 sg13g2_fill_2 FILLER_44_1291 ();
 sg13g2_fill_2 FILLER_44_1301 ();
 sg13g2_fill_1 FILLER_44_1317 ();
 sg13g2_decap_8 FILLER_44_1322 ();
 sg13g2_decap_4 FILLER_44_1329 ();
 sg13g2_fill_2 FILLER_44_1333 ();
 sg13g2_decap_8 FILLER_44_1349 ();
 sg13g2_fill_2 FILLER_44_1356 ();
 sg13g2_fill_1 FILLER_44_1358 ();
 sg13g2_decap_8 FILLER_44_1373 ();
 sg13g2_decap_8 FILLER_44_1380 ();
 sg13g2_decap_8 FILLER_44_1387 ();
 sg13g2_fill_2 FILLER_44_1434 ();
 sg13g2_fill_1 FILLER_44_1456 ();
 sg13g2_fill_2 FILLER_44_1470 ();
 sg13g2_fill_1 FILLER_44_1472 ();
 sg13g2_fill_2 FILLER_44_1486 ();
 sg13g2_fill_1 FILLER_44_1488 ();
 sg13g2_decap_8 FILLER_44_1497 ();
 sg13g2_decap_8 FILLER_44_1504 ();
 sg13g2_decap_4 FILLER_44_1511 ();
 sg13g2_fill_1 FILLER_44_1515 ();
 sg13g2_decap_4 FILLER_44_1537 ();
 sg13g2_fill_1 FILLER_44_1541 ();
 sg13g2_decap_8 FILLER_44_1555 ();
 sg13g2_fill_1 FILLER_44_1562 ();
 sg13g2_decap_4 FILLER_44_1569 ();
 sg13g2_fill_1 FILLER_44_1573 ();
 sg13g2_decap_8 FILLER_44_1578 ();
 sg13g2_fill_1 FILLER_44_1585 ();
 sg13g2_fill_2 FILLER_44_1620 ();
 sg13g2_fill_1 FILLER_44_1622 ();
 sg13g2_fill_1 FILLER_44_1630 ();
 sg13g2_fill_2 FILLER_44_1649 ();
 sg13g2_fill_1 FILLER_44_1651 ();
 sg13g2_decap_8 FILLER_44_1672 ();
 sg13g2_fill_1 FILLER_44_1679 ();
 sg13g2_decap_4 FILLER_44_1688 ();
 sg13g2_fill_2 FILLER_44_1692 ();
 sg13g2_fill_2 FILLER_44_1707 ();
 sg13g2_fill_1 FILLER_44_1709 ();
 sg13g2_decap_4 FILLER_44_1719 ();
 sg13g2_fill_2 FILLER_44_1723 ();
 sg13g2_fill_1 FILLER_44_1744 ();
 sg13g2_fill_2 FILLER_44_1766 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_58 ();
 sg13g2_fill_1 FILLER_45_60 ();
 sg13g2_decap_8 FILLER_45_75 ();
 sg13g2_fill_1 FILLER_45_82 ();
 sg13g2_fill_2 FILLER_45_97 ();
 sg13g2_fill_1 FILLER_45_109 ();
 sg13g2_fill_1 FILLER_45_146 ();
 sg13g2_decap_4 FILLER_45_156 ();
 sg13g2_fill_2 FILLER_45_191 ();
 sg13g2_fill_1 FILLER_45_193 ();
 sg13g2_fill_1 FILLER_45_241 ();
 sg13g2_decap_4 FILLER_45_256 ();
 sg13g2_fill_2 FILLER_45_260 ();
 sg13g2_fill_1 FILLER_45_265 ();
 sg13g2_decap_8 FILLER_45_284 ();
 sg13g2_fill_1 FILLER_45_291 ();
 sg13g2_fill_1 FILLER_45_309 ();
 sg13g2_fill_1 FILLER_45_337 ();
 sg13g2_fill_2 FILLER_45_364 ();
 sg13g2_fill_1 FILLER_45_366 ();
 sg13g2_fill_1 FILLER_45_395 ();
 sg13g2_decap_4 FILLER_45_422 ();
 sg13g2_fill_1 FILLER_45_459 ();
 sg13g2_fill_2 FILLER_45_465 ();
 sg13g2_fill_1 FILLER_45_467 ();
 sg13g2_fill_1 FILLER_45_482 ();
 sg13g2_fill_2 FILLER_45_495 ();
 sg13g2_fill_2 FILLER_45_501 ();
 sg13g2_fill_2 FILLER_45_524 ();
 sg13g2_fill_1 FILLER_45_526 ();
 sg13g2_decap_4 FILLER_45_564 ();
 sg13g2_fill_2 FILLER_45_568 ();
 sg13g2_fill_2 FILLER_45_623 ();
 sg13g2_fill_1 FILLER_45_638 ();
 sg13g2_fill_1 FILLER_45_648 ();
 sg13g2_fill_2 FILLER_45_663 ();
 sg13g2_fill_1 FILLER_45_665 ();
 sg13g2_fill_1 FILLER_45_702 ();
 sg13g2_fill_1 FILLER_45_730 ();
 sg13g2_fill_2 FILLER_45_752 ();
 sg13g2_fill_1 FILLER_45_781 ();
 sg13g2_fill_2 FILLER_45_809 ();
 sg13g2_fill_1 FILLER_45_843 ();
 sg13g2_decap_8 FILLER_45_862 ();
 sg13g2_decap_4 FILLER_45_873 ();
 sg13g2_fill_2 FILLER_45_877 ();
 sg13g2_fill_2 FILLER_45_893 ();
 sg13g2_fill_2 FILLER_45_899 ();
 sg13g2_fill_1 FILLER_45_901 ();
 sg13g2_fill_2 FILLER_45_911 ();
 sg13g2_fill_1 FILLER_45_913 ();
 sg13g2_fill_2 FILLER_45_918 ();
 sg13g2_fill_1 FILLER_45_947 ();
 sg13g2_decap_4 FILLER_45_995 ();
 sg13g2_fill_1 FILLER_45_1005 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_fill_2 FILLER_45_1077 ();
 sg13g2_fill_1 FILLER_45_1079 ();
 sg13g2_fill_1 FILLER_45_1090 ();
 sg13g2_fill_1 FILLER_45_1110 ();
 sg13g2_fill_1 FILLER_45_1125 ();
 sg13g2_decap_4 FILLER_45_1158 ();
 sg13g2_fill_2 FILLER_45_1171 ();
 sg13g2_fill_1 FILLER_45_1173 ();
 sg13g2_fill_2 FILLER_45_1196 ();
 sg13g2_fill_1 FILLER_45_1208 ();
 sg13g2_fill_1 FILLER_45_1218 ();
 sg13g2_decap_4 FILLER_45_1242 ();
 sg13g2_fill_2 FILLER_45_1246 ();
 sg13g2_fill_2 FILLER_45_1255 ();
 sg13g2_decap_8 FILLER_45_1260 ();
 sg13g2_decap_4 FILLER_45_1267 ();
 sg13g2_fill_2 FILLER_45_1271 ();
 sg13g2_decap_4 FILLER_45_1291 ();
 sg13g2_fill_1 FILLER_45_1295 ();
 sg13g2_fill_2 FILLER_45_1305 ();
 sg13g2_fill_1 FILLER_45_1312 ();
 sg13g2_decap_8 FILLER_45_1318 ();
 sg13g2_fill_2 FILLER_45_1325 ();
 sg13g2_decap_8 FILLER_45_1331 ();
 sg13g2_decap_8 FILLER_45_1343 ();
 sg13g2_decap_8 FILLER_45_1350 ();
 sg13g2_fill_2 FILLER_45_1357 ();
 sg13g2_decap_8 FILLER_45_1370 ();
 sg13g2_decap_4 FILLER_45_1377 ();
 sg13g2_decap_8 FILLER_45_1413 ();
 sg13g2_fill_1 FILLER_45_1420 ();
 sg13g2_decap_8 FILLER_45_1433 ();
 sg13g2_fill_2 FILLER_45_1449 ();
 sg13g2_fill_1 FILLER_45_1451 ();
 sg13g2_decap_8 FILLER_45_1457 ();
 sg13g2_decap_8 FILLER_45_1464 ();
 sg13g2_fill_2 FILLER_45_1489 ();
 sg13g2_decap_4 FILLER_45_1503 ();
 sg13g2_fill_1 FILLER_45_1507 ();
 sg13g2_decap_4 FILLER_45_1519 ();
 sg13g2_fill_2 FILLER_45_1523 ();
 sg13g2_decap_4 FILLER_45_1535 ();
 sg13g2_fill_2 FILLER_45_1539 ();
 sg13g2_fill_1 FILLER_45_1549 ();
 sg13g2_decap_8 FILLER_45_1562 ();
 sg13g2_decap_8 FILLER_45_1569 ();
 sg13g2_decap_8 FILLER_45_1589 ();
 sg13g2_decap_8 FILLER_45_1596 ();
 sg13g2_decap_4 FILLER_45_1603 ();
 sg13g2_fill_1 FILLER_45_1607 ();
 sg13g2_decap_8 FILLER_45_1614 ();
 sg13g2_decap_4 FILLER_45_1621 ();
 sg13g2_decap_4 FILLER_45_1630 ();
 sg13g2_fill_1 FILLER_45_1638 ();
 sg13g2_decap_4 FILLER_45_1647 ();
 sg13g2_decap_8 FILLER_45_1664 ();
 sg13g2_decap_8 FILLER_45_1671 ();
 sg13g2_fill_2 FILLER_45_1678 ();
 sg13g2_decap_8 FILLER_45_1694 ();
 sg13g2_decap_8 FILLER_45_1724 ();
 sg13g2_fill_2 FILLER_45_1745 ();
 sg13g2_fill_1 FILLER_45_1747 ();
 sg13g2_decap_8 FILLER_45_1756 ();
 sg13g2_decap_4 FILLER_45_1763 ();
 sg13g2_fill_1 FILLER_45_1767 ();
 sg13g2_fill_1 FILLER_46_32 ();
 sg13g2_fill_1 FILLER_46_42 ();
 sg13g2_fill_1 FILLER_46_61 ();
 sg13g2_fill_1 FILLER_46_149 ();
 sg13g2_decap_4 FILLER_46_155 ();
 sg13g2_fill_2 FILLER_46_159 ();
 sg13g2_fill_2 FILLER_46_196 ();
 sg13g2_fill_1 FILLER_46_297 ();
 sg13g2_fill_2 FILLER_46_347 ();
 sg13g2_fill_1 FILLER_46_358 ();
 sg13g2_fill_2 FILLER_46_392 ();
 sg13g2_fill_1 FILLER_46_394 ();
 sg13g2_fill_1 FILLER_46_400 ();
 sg13g2_fill_2 FILLER_46_434 ();
 sg13g2_decap_4 FILLER_46_454 ();
 sg13g2_fill_2 FILLER_46_458 ();
 sg13g2_fill_1 FILLER_46_492 ();
 sg13g2_fill_1 FILLER_46_498 ();
 sg13g2_fill_2 FILLER_46_508 ();
 sg13g2_fill_1 FILLER_46_510 ();
 sg13g2_fill_2 FILLER_46_520 ();
 sg13g2_fill_2 FILLER_46_531 ();
 sg13g2_fill_1 FILLER_46_533 ();
 sg13g2_fill_2 FILLER_46_556 ();
 sg13g2_fill_2 FILLER_46_563 ();
 sg13g2_fill_1 FILLER_46_565 ();
 sg13g2_fill_2 FILLER_46_583 ();
 sg13g2_fill_2 FILLER_46_631 ();
 sg13g2_fill_1 FILLER_46_633 ();
 sg13g2_fill_2 FILLER_46_647 ();
 sg13g2_fill_2 FILLER_46_662 ();
 sg13g2_fill_1 FILLER_46_747 ();
 sg13g2_fill_1 FILLER_46_762 ();
 sg13g2_fill_2 FILLER_46_778 ();
 sg13g2_fill_1 FILLER_46_780 ();
 sg13g2_decap_4 FILLER_46_793 ();
 sg13g2_fill_1 FILLER_46_797 ();
 sg13g2_fill_1 FILLER_46_806 ();
 sg13g2_fill_1 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_939 ();
 sg13g2_fill_1 FILLER_46_972 ();
 sg13g2_fill_2 FILLER_46_979 ();
 sg13g2_fill_1 FILLER_46_981 ();
 sg13g2_decap_8 FILLER_46_991 ();
 sg13g2_decap_8 FILLER_46_998 ();
 sg13g2_fill_1 FILLER_46_1005 ();
 sg13g2_fill_1 FILLER_46_1034 ();
 sg13g2_fill_1 FILLER_46_1048 ();
 sg13g2_fill_2 FILLER_46_1077 ();
 sg13g2_fill_2 FILLER_46_1089 ();
 sg13g2_fill_2 FILLER_46_1101 ();
 sg13g2_fill_1 FILLER_46_1103 ();
 sg13g2_decap_8 FILLER_46_1112 ();
 sg13g2_fill_2 FILLER_46_1119 ();
 sg13g2_decap_4 FILLER_46_1158 ();
 sg13g2_fill_1 FILLER_46_1198 ();
 sg13g2_fill_1 FILLER_46_1239 ();
 sg13g2_decap_8 FILLER_46_1268 ();
 sg13g2_fill_2 FILLER_46_1275 ();
 sg13g2_fill_1 FILLER_46_1277 ();
 sg13g2_fill_2 FILLER_46_1286 ();
 sg13g2_fill_1 FILLER_46_1292 ();
 sg13g2_fill_1 FILLER_46_1327 ();
 sg13g2_fill_2 FILLER_46_1341 ();
 sg13g2_fill_1 FILLER_46_1346 ();
 sg13g2_decap_4 FILLER_46_1350 ();
 sg13g2_fill_2 FILLER_46_1354 ();
 sg13g2_fill_1 FILLER_46_1369 ();
 sg13g2_decap_4 FILLER_46_1394 ();
 sg13g2_fill_1 FILLER_46_1398 ();
 sg13g2_decap_4 FILLER_46_1415 ();
 sg13g2_fill_2 FILLER_46_1419 ();
 sg13g2_fill_2 FILLER_46_1426 ();
 sg13g2_decap_8 FILLER_46_1431 ();
 sg13g2_fill_2 FILLER_46_1438 ();
 sg13g2_decap_8 FILLER_46_1460 ();
 sg13g2_decap_8 FILLER_46_1467 ();
 sg13g2_decap_4 FILLER_46_1474 ();
 sg13g2_fill_1 FILLER_46_1478 ();
 sg13g2_fill_1 FILLER_46_1499 ();
 sg13g2_decap_8 FILLER_46_1513 ();
 sg13g2_fill_2 FILLER_46_1520 ();
 sg13g2_fill_1 FILLER_46_1522 ();
 sg13g2_decap_8 FILLER_46_1541 ();
 sg13g2_fill_1 FILLER_46_1548 ();
 sg13g2_decap_8 FILLER_46_1564 ();
 sg13g2_decap_4 FILLER_46_1571 ();
 sg13g2_fill_1 FILLER_46_1575 ();
 sg13g2_decap_4 FILLER_46_1594 ();
 sg13g2_fill_1 FILLER_46_1598 ();
 sg13g2_decap_8 FILLER_46_1639 ();
 sg13g2_fill_1 FILLER_46_1646 ();
 sg13g2_fill_1 FILLER_46_1673 ();
 sg13g2_fill_2 FILLER_46_1702 ();
 sg13g2_fill_1 FILLER_46_1704 ();
 sg13g2_fill_1 FILLER_46_1714 ();
 sg13g2_fill_2 FILLER_46_1720 ();
 sg13g2_fill_1 FILLER_46_1722 ();
 sg13g2_fill_2 FILLER_46_1737 ();
 sg13g2_fill_1 FILLER_46_1739 ();
 sg13g2_decap_4 FILLER_46_1764 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_7 ();
 sg13g2_fill_1 FILLER_47_48 ();
 sg13g2_fill_2 FILLER_47_69 ();
 sg13g2_decap_4 FILLER_47_75 ();
 sg13g2_fill_1 FILLER_47_79 ();
 sg13g2_fill_1 FILLER_47_197 ();
 sg13g2_decap_8 FILLER_47_234 ();
 sg13g2_decap_4 FILLER_47_241 ();
 sg13g2_fill_2 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_251 ();
 sg13g2_decap_4 FILLER_47_258 ();
 sg13g2_fill_2 FILLER_47_294 ();
 sg13g2_fill_2 FILLER_47_329 ();
 sg13g2_fill_1 FILLER_47_364 ();
 sg13g2_fill_2 FILLER_47_419 ();
 sg13g2_fill_1 FILLER_47_421 ();
 sg13g2_fill_2 FILLER_47_433 ();
 sg13g2_fill_1 FILLER_47_435 ();
 sg13g2_fill_2 FILLER_47_441 ();
 sg13g2_fill_1 FILLER_47_443 ();
 sg13g2_decap_4 FILLER_47_449 ();
 sg13g2_fill_1 FILLER_47_453 ();
 sg13g2_fill_1 FILLER_47_459 ();
 sg13g2_fill_2 FILLER_47_469 ();
 sg13g2_fill_1 FILLER_47_471 ();
 sg13g2_fill_2 FILLER_47_492 ();
 sg13g2_fill_1 FILLER_47_494 ();
 sg13g2_fill_2 FILLER_47_528 ();
 sg13g2_fill_1 FILLER_47_530 ();
 sg13g2_decap_4 FILLER_47_611 ();
 sg13g2_fill_1 FILLER_47_635 ();
 sg13g2_fill_2 FILLER_47_663 ();
 sg13g2_decap_8 FILLER_47_710 ();
 sg13g2_decap_4 FILLER_47_717 ();
 sg13g2_decap_4 FILLER_47_730 ();
 sg13g2_fill_1 FILLER_47_775 ();
 sg13g2_decap_4 FILLER_47_839 ();
 sg13g2_decap_8 FILLER_47_860 ();
 sg13g2_fill_1 FILLER_47_893 ();
 sg13g2_decap_4 FILLER_47_903 ();
 sg13g2_fill_1 FILLER_47_907 ();
 sg13g2_fill_2 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_967 ();
 sg13g2_fill_2 FILLER_47_974 ();
 sg13g2_fill_2 FILLER_47_1028 ();
 sg13g2_fill_1 FILLER_47_1030 ();
 sg13g2_fill_2 FILLER_47_1040 ();
 sg13g2_fill_1 FILLER_47_1042 ();
 sg13g2_fill_1 FILLER_47_1079 ();
 sg13g2_decap_8 FILLER_47_1100 ();
 sg13g2_fill_2 FILLER_47_1127 ();
 sg13g2_decap_4 FILLER_47_1152 ();
 sg13g2_fill_2 FILLER_47_1217 ();
 sg13g2_decap_8 FILLER_47_1266 ();
 sg13g2_fill_1 FILLER_47_1273 ();
 sg13g2_fill_1 FILLER_47_1301 ();
 sg13g2_fill_2 FILLER_47_1346 ();
 sg13g2_decap_8 FILLER_47_1377 ();
 sg13g2_decap_8 FILLER_47_1384 ();
 sg13g2_decap_4 FILLER_47_1391 ();
 sg13g2_fill_2 FILLER_47_1416 ();
 sg13g2_fill_1 FILLER_47_1418 ();
 sg13g2_fill_1 FILLER_47_1424 ();
 sg13g2_decap_4 FILLER_47_1443 ();
 sg13g2_fill_2 FILLER_47_1447 ();
 sg13g2_fill_2 FILLER_47_1453 ();
 sg13g2_fill_1 FILLER_47_1455 ();
 sg13g2_decap_8 FILLER_47_1464 ();
 sg13g2_decap_4 FILLER_47_1471 ();
 sg13g2_fill_1 FILLER_47_1475 ();
 sg13g2_fill_2 FILLER_47_1489 ();
 sg13g2_decap_8 FILLER_47_1496 ();
 sg13g2_decap_4 FILLER_47_1503 ();
 sg13g2_fill_1 FILLER_47_1520 ();
 sg13g2_decap_8 FILLER_47_1537 ();
 sg13g2_decap_4 FILLER_47_1544 ();
 sg13g2_decap_8 FILLER_47_1563 ();
 sg13g2_fill_2 FILLER_47_1570 ();
 sg13g2_fill_1 FILLER_47_1572 ();
 sg13g2_fill_2 FILLER_47_1598 ();
 sg13g2_decap_8 FILLER_47_1617 ();
 sg13g2_decap_8 FILLER_47_1624 ();
 sg13g2_fill_2 FILLER_47_1631 ();
 sg13g2_decap_8 FILLER_47_1637 ();
 sg13g2_fill_2 FILLER_47_1644 ();
 sg13g2_decap_8 FILLER_47_1667 ();
 sg13g2_fill_1 FILLER_47_1689 ();
 sg13g2_decap_8 FILLER_47_1702 ();
 sg13g2_fill_2 FILLER_47_1709 ();
 sg13g2_fill_1 FILLER_47_1716 ();
 sg13g2_decap_8 FILLER_47_1726 ();
 sg13g2_fill_2 FILLER_47_1733 ();
 sg13g2_fill_1 FILLER_47_1746 ();
 sg13g2_decap_8 FILLER_47_1756 ();
 sg13g2_decap_4 FILLER_47_1763 ();
 sg13g2_fill_1 FILLER_47_1767 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_51 ();
 sg13g2_fill_2 FILLER_48_105 ();
 sg13g2_fill_1 FILLER_48_107 ();
 sg13g2_fill_1 FILLER_48_126 ();
 sg13g2_decap_4 FILLER_48_146 ();
 sg13g2_fill_1 FILLER_48_150 ();
 sg13g2_fill_1 FILLER_48_155 ();
 sg13g2_fill_2 FILLER_48_160 ();
 sg13g2_fill_2 FILLER_48_177 ();
 sg13g2_fill_2 FILLER_48_224 ();
 sg13g2_fill_1 FILLER_48_226 ();
 sg13g2_fill_2 FILLER_48_240 ();
 sg13g2_fill_1 FILLER_48_242 ();
 sg13g2_fill_2 FILLER_48_249 ();
 sg13g2_fill_2 FILLER_48_297 ();
 sg13g2_fill_2 FILLER_48_321 ();
 sg13g2_fill_1 FILLER_48_323 ();
 sg13g2_fill_1 FILLER_48_347 ();
 sg13g2_fill_1 FILLER_48_373 ();
 sg13g2_fill_2 FILLER_48_383 ();
 sg13g2_fill_2 FILLER_48_426 ();
 sg13g2_decap_4 FILLER_48_445 ();
 sg13g2_fill_1 FILLER_48_487 ();
 sg13g2_decap_4 FILLER_48_525 ();
 sg13g2_fill_2 FILLER_48_529 ();
 sg13g2_fill_2 FILLER_48_540 ();
 sg13g2_decap_4 FILLER_48_559 ();
 sg13g2_fill_1 FILLER_48_576 ();
 sg13g2_fill_2 FILLER_48_621 ();
 sg13g2_fill_1 FILLER_48_653 ();
 sg13g2_decap_8 FILLER_48_705 ();
 sg13g2_decap_4 FILLER_48_712 ();
 sg13g2_decap_8 FILLER_48_726 ();
 sg13g2_decap_8 FILLER_48_733 ();
 sg13g2_decap_4 FILLER_48_789 ();
 sg13g2_fill_2 FILLER_48_793 ();
 sg13g2_fill_2 FILLER_48_808 ();
 sg13g2_fill_1 FILLER_48_810 ();
 sg13g2_fill_1 FILLER_48_824 ();
 sg13g2_decap_4 FILLER_48_834 ();
 sg13g2_fill_2 FILLER_48_838 ();
 sg13g2_decap_4 FILLER_48_843 ();
 sg13g2_decap_8 FILLER_48_885 ();
 sg13g2_decap_4 FILLER_48_892 ();
 sg13g2_fill_2 FILLER_48_896 ();
 sg13g2_fill_2 FILLER_48_926 ();
 sg13g2_decap_4 FILLER_48_941 ();
 sg13g2_fill_1 FILLER_48_945 ();
 sg13g2_fill_2 FILLER_48_977 ();
 sg13g2_fill_2 FILLER_48_1034 ();
 sg13g2_fill_1 FILLER_48_1079 ();
 sg13g2_fill_1 FILLER_48_1090 ();
 sg13g2_fill_1 FILLER_48_1132 ();
 sg13g2_fill_2 FILLER_48_1138 ();
 sg13g2_fill_1 FILLER_48_1140 ();
 sg13g2_fill_1 FILLER_48_1145 ();
 sg13g2_fill_1 FILLER_48_1156 ();
 sg13g2_decap_8 FILLER_48_1174 ();
 sg13g2_fill_2 FILLER_48_1181 ();
 sg13g2_fill_1 FILLER_48_1183 ();
 sg13g2_decap_4 FILLER_48_1188 ();
 sg13g2_fill_1 FILLER_48_1192 ();
 sg13g2_fill_2 FILLER_48_1222 ();
 sg13g2_fill_1 FILLER_48_1224 ();
 sg13g2_decap_4 FILLER_48_1244 ();
 sg13g2_fill_2 FILLER_48_1248 ();
 sg13g2_decap_8 FILLER_48_1260 ();
 sg13g2_decap_8 FILLER_48_1267 ();
 sg13g2_fill_1 FILLER_48_1294 ();
 sg13g2_fill_2 FILLER_48_1325 ();
 sg13g2_fill_1 FILLER_48_1327 ();
 sg13g2_decap_8 FILLER_48_1338 ();
 sg13g2_decap_8 FILLER_48_1345 ();
 sg13g2_fill_2 FILLER_48_1352 ();
 sg13g2_fill_2 FILLER_48_1379 ();
 sg13g2_fill_1 FILLER_48_1381 ();
 sg13g2_decap_8 FILLER_48_1390 ();
 sg13g2_fill_2 FILLER_48_1397 ();
 sg13g2_fill_2 FILLER_48_1412 ();
 sg13g2_fill_1 FILLER_48_1424 ();
 sg13g2_decap_8 FILLER_48_1430 ();
 sg13g2_decap_8 FILLER_48_1437 ();
 sg13g2_decap_8 FILLER_48_1444 ();
 sg13g2_decap_8 FILLER_48_1451 ();
 sg13g2_decap_8 FILLER_48_1458 ();
 sg13g2_fill_1 FILLER_48_1477 ();
 sg13g2_fill_1 FILLER_48_1486 ();
 sg13g2_fill_2 FILLER_48_1495 ();
 sg13g2_fill_1 FILLER_48_1512 ();
 sg13g2_decap_4 FILLER_48_1534 ();
 sg13g2_decap_8 FILLER_48_1558 ();
 sg13g2_decap_8 FILLER_48_1565 ();
 sg13g2_fill_2 FILLER_48_1572 ();
 sg13g2_fill_1 FILLER_48_1574 ();
 sg13g2_decap_8 FILLER_48_1594 ();
 sg13g2_decap_4 FILLER_48_1617 ();
 sg13g2_fill_2 FILLER_48_1639 ();
 sg13g2_fill_2 FILLER_48_1645 ();
 sg13g2_fill_1 FILLER_48_1647 ();
 sg13g2_fill_1 FILLER_48_1652 ();
 sg13g2_decap_8 FILLER_48_1668 ();
 sg13g2_decap_4 FILLER_48_1675 ();
 sg13g2_fill_2 FILLER_48_1679 ();
 sg13g2_fill_2 FILLER_48_1703 ();
 sg13g2_fill_1 FILLER_48_1705 ();
 sg13g2_fill_1 FILLER_48_1721 ();
 sg13g2_fill_2 FILLER_48_1730 ();
 sg13g2_fill_1 FILLER_48_1748 ();
 sg13g2_fill_2 FILLER_48_1765 ();
 sg13g2_fill_1 FILLER_48_1767 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_51 ();
 sg13g2_fill_1 FILLER_49_97 ();
 sg13g2_fill_1 FILLER_49_177 ();
 sg13g2_fill_1 FILLER_49_268 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_295 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_330 ();
 sg13g2_fill_1 FILLER_49_332 ();
 sg13g2_decap_4 FILLER_49_365 ();
 sg13g2_fill_2 FILLER_49_409 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_decap_4 FILLER_49_422 ();
 sg13g2_fill_1 FILLER_49_426 ();
 sg13g2_fill_2 FILLER_49_441 ();
 sg13g2_fill_1 FILLER_49_466 ();
 sg13g2_decap_4 FILLER_49_475 ();
 sg13g2_fill_1 FILLER_49_489 ();
 sg13g2_fill_1 FILLER_49_494 ();
 sg13g2_fill_1 FILLER_49_521 ();
 sg13g2_decap_8 FILLER_49_550 ();
 sg13g2_decap_4 FILLER_49_557 ();
 sg13g2_fill_2 FILLER_49_561 ();
 sg13g2_fill_2 FILLER_49_589 ();
 sg13g2_fill_2 FILLER_49_604 ();
 sg13g2_decap_8 FILLER_49_638 ();
 sg13g2_decap_8 FILLER_49_645 ();
 sg13g2_fill_1 FILLER_49_652 ();
 sg13g2_fill_2 FILLER_49_657 ();
 sg13g2_fill_1 FILLER_49_676 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_fill_2 FILLER_49_749 ();
 sg13g2_fill_2 FILLER_49_764 ();
 sg13g2_fill_1 FILLER_49_766 ();
 sg13g2_fill_1 FILLER_49_772 ();
 sg13g2_fill_1 FILLER_49_795 ();
 sg13g2_decap_8 FILLER_49_912 ();
 sg13g2_fill_1 FILLER_49_919 ();
 sg13g2_fill_2 FILLER_49_928 ();
 sg13g2_fill_1 FILLER_49_930 ();
 sg13g2_fill_2 FILLER_49_974 ();
 sg13g2_fill_1 FILLER_49_1009 ();
 sg13g2_fill_2 FILLER_49_1023 ();
 sg13g2_fill_1 FILLER_49_1025 ();
 sg13g2_fill_2 FILLER_49_1049 ();
 sg13g2_fill_2 FILLER_49_1060 ();
 sg13g2_fill_1 FILLER_49_1062 ();
 sg13g2_fill_2 FILLER_49_1076 ();
 sg13g2_fill_1 FILLER_49_1078 ();
 sg13g2_fill_2 FILLER_49_1089 ();
 sg13g2_fill_2 FILLER_49_1106 ();
 sg13g2_fill_1 FILLER_49_1108 ();
 sg13g2_fill_1 FILLER_49_1150 ();
 sg13g2_decap_8 FILLER_49_1194 ();
 sg13g2_decap_4 FILLER_49_1201 ();
 sg13g2_fill_1 FILLER_49_1205 ();
 sg13g2_fill_2 FILLER_49_1295 ();
 sg13g2_decap_4 FILLER_49_1315 ();
 sg13g2_decap_4 FILLER_49_1323 ();
 sg13g2_fill_1 FILLER_49_1327 ();
 sg13g2_decap_8 FILLER_49_1338 ();
 sg13g2_decap_8 FILLER_49_1345 ();
 sg13g2_fill_2 FILLER_49_1379 ();
 sg13g2_fill_1 FILLER_49_1381 ();
 sg13g2_decap_8 FILLER_49_1404 ();
 sg13g2_fill_2 FILLER_49_1411 ();
 sg13g2_fill_1 FILLER_49_1413 ();
 sg13g2_fill_2 FILLER_49_1433 ();
 sg13g2_fill_1 FILLER_49_1435 ();
 sg13g2_decap_8 FILLER_49_1442 ();
 sg13g2_decap_8 FILLER_49_1464 ();
 sg13g2_decap_4 FILLER_49_1471 ();
 sg13g2_decap_4 FILLER_49_1493 ();
 sg13g2_fill_1 FILLER_49_1497 ();
 sg13g2_decap_8 FILLER_49_1516 ();
 sg13g2_fill_1 FILLER_49_1523 ();
 sg13g2_decap_8 FILLER_49_1563 ();
 sg13g2_decap_8 FILLER_49_1570 ();
 sg13g2_fill_1 FILLER_49_1577 ();
 sg13g2_fill_2 FILLER_49_1595 ();
 sg13g2_fill_1 FILLER_49_1597 ();
 sg13g2_decap_4 FILLER_49_1607 ();
 sg13g2_fill_1 FILLER_49_1611 ();
 sg13g2_decap_8 FILLER_49_1622 ();
 sg13g2_decap_8 FILLER_49_1629 ();
 sg13g2_fill_1 FILLER_49_1636 ();
 sg13g2_decap_8 FILLER_49_1657 ();
 sg13g2_fill_2 FILLER_49_1664 ();
 sg13g2_decap_4 FILLER_49_1670 ();
 sg13g2_fill_1 FILLER_49_1674 ();
 sg13g2_fill_1 FILLER_49_1688 ();
 sg13g2_decap_8 FILLER_49_1703 ();
 sg13g2_decap_8 FILLER_49_1715 ();
 sg13g2_decap_8 FILLER_49_1722 ();
 sg13g2_decap_4 FILLER_49_1729 ();
 sg13g2_fill_2 FILLER_49_1733 ();
 sg13g2_fill_1 FILLER_49_1749 ();
 sg13g2_decap_4 FILLER_49_1763 ();
 sg13g2_fill_1 FILLER_49_1767 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_7 ();
 sg13g2_fill_1 FILLER_50_9 ();
 sg13g2_fill_1 FILLER_50_67 ();
 sg13g2_decap_4 FILLER_50_104 ();
 sg13g2_fill_2 FILLER_50_123 ();
 sg13g2_fill_2 FILLER_50_145 ();
 sg13g2_fill_2 FILLER_50_156 ();
 sg13g2_fill_1 FILLER_50_194 ();
 sg13g2_fill_1 FILLER_50_211 ();
 sg13g2_fill_2 FILLER_50_221 ();
 sg13g2_decap_8 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_254 ();
 sg13g2_fill_1 FILLER_50_256 ();
 sg13g2_fill_2 FILLER_50_301 ();
 sg13g2_fill_2 FILLER_50_317 ();
 sg13g2_decap_4 FILLER_50_343 ();
 sg13g2_decap_4 FILLER_50_400 ();
 sg13g2_fill_2 FILLER_50_431 ();
 sg13g2_fill_2 FILLER_50_454 ();
 sg13g2_fill_1 FILLER_50_456 ();
 sg13g2_fill_2 FILLER_50_462 ();
 sg13g2_fill_1 FILLER_50_464 ();
 sg13g2_decap_8 FILLER_50_480 ();
 sg13g2_decap_4 FILLER_50_487 ();
 sg13g2_fill_1 FILLER_50_491 ();
 sg13g2_decap_4 FILLER_50_502 ();
 sg13g2_fill_2 FILLER_50_546 ();
 sg13g2_decap_4 FILLER_50_570 ();
 sg13g2_decap_4 FILLER_50_579 ();
 sg13g2_fill_2 FILLER_50_583 ();
 sg13g2_decap_4 FILLER_50_595 ();
 sg13g2_fill_2 FILLER_50_599 ();
 sg13g2_fill_2 FILLER_50_611 ();
 sg13g2_fill_1 FILLER_50_613 ();
 sg13g2_decap_4 FILLER_50_643 ();
 sg13g2_fill_2 FILLER_50_662 ();
 sg13g2_fill_1 FILLER_50_664 ();
 sg13g2_fill_2 FILLER_50_675 ();
 sg13g2_fill_1 FILLER_50_677 ();
 sg13g2_fill_2 FILLER_50_700 ();
 sg13g2_decap_4 FILLER_50_711 ();
 sg13g2_fill_1 FILLER_50_715 ();
 sg13g2_decap_8 FILLER_50_725 ();
 sg13g2_fill_2 FILLER_50_732 ();
 sg13g2_fill_1 FILLER_50_734 ();
 sg13g2_fill_1 FILLER_50_771 ();
 sg13g2_fill_1 FILLER_50_805 ();
 sg13g2_decap_4 FILLER_50_810 ();
 sg13g2_fill_2 FILLER_50_814 ();
 sg13g2_decap_8 FILLER_50_824 ();
 sg13g2_decap_4 FILLER_50_856 ();
 sg13g2_fill_1 FILLER_50_860 ();
 sg13g2_fill_1 FILLER_50_877 ();
 sg13g2_fill_1 FILLER_50_918 ();
 sg13g2_fill_2 FILLER_50_946 ();
 sg13g2_fill_2 FILLER_50_979 ();
 sg13g2_fill_1 FILLER_50_994 ();
 sg13g2_fill_2 FILLER_50_1008 ();
 sg13g2_fill_1 FILLER_50_1010 ();
 sg13g2_fill_2 FILLER_50_1048 ();
 sg13g2_fill_1 FILLER_50_1078 ();
 sg13g2_fill_2 FILLER_50_1089 ();
 sg13g2_fill_1 FILLER_50_1091 ();
 sg13g2_decap_8 FILLER_50_1102 ();
 sg13g2_decap_4 FILLER_50_1109 ();
 sg13g2_fill_1 FILLER_50_1113 ();
 sg13g2_decap_8 FILLER_50_1141 ();
 sg13g2_fill_2 FILLER_50_1148 ();
 sg13g2_fill_1 FILLER_50_1150 ();
 sg13g2_decap_4 FILLER_50_1173 ();
 sg13g2_fill_2 FILLER_50_1177 ();
 sg13g2_decap_8 FILLER_50_1191 ();
 sg13g2_decap_8 FILLER_50_1198 ();
 sg13g2_decap_4 FILLER_50_1205 ();
 sg13g2_fill_1 FILLER_50_1218 ();
 sg13g2_decap_8 FILLER_50_1252 ();
 sg13g2_decap_8 FILLER_50_1262 ();
 sg13g2_decap_8 FILLER_50_1269 ();
 sg13g2_decap_8 FILLER_50_1276 ();
 sg13g2_decap_4 FILLER_50_1283 ();
 sg13g2_fill_2 FILLER_50_1305 ();
 sg13g2_fill_2 FILLER_50_1322 ();
 sg13g2_fill_1 FILLER_50_1324 ();
 sg13g2_decap_8 FILLER_50_1339 ();
 sg13g2_decap_4 FILLER_50_1346 ();
 sg13g2_fill_2 FILLER_50_1365 ();
 sg13g2_fill_1 FILLER_50_1367 ();
 sg13g2_decap_4 FILLER_50_1386 ();
 sg13g2_fill_1 FILLER_50_1390 ();
 sg13g2_decap_4 FILLER_50_1405 ();
 sg13g2_fill_2 FILLER_50_1427 ();
 sg13g2_fill_2 FILLER_50_1439 ();
 sg13g2_fill_1 FILLER_50_1441 ();
 sg13g2_decap_8 FILLER_50_1468 ();
 sg13g2_decap_4 FILLER_50_1475 ();
 sg13g2_fill_2 FILLER_50_1479 ();
 sg13g2_decap_8 FILLER_50_1485 ();
 sg13g2_decap_4 FILLER_50_1492 ();
 sg13g2_fill_2 FILLER_50_1496 ();
 sg13g2_fill_2 FILLER_50_1511 ();
 sg13g2_fill_1 FILLER_50_1513 ();
 sg13g2_decap_8 FILLER_50_1522 ();
 sg13g2_decap_8 FILLER_50_1529 ();
 sg13g2_decap_4 FILLER_50_1536 ();
 sg13g2_fill_2 FILLER_50_1540 ();
 sg13g2_decap_8 FILLER_50_1560 ();
 sg13g2_fill_1 FILLER_50_1567 ();
 sg13g2_decap_8 FILLER_50_1593 ();
 sg13g2_decap_8 FILLER_50_1600 ();
 sg13g2_fill_2 FILLER_50_1607 ();
 sg13g2_fill_1 FILLER_50_1609 ();
 sg13g2_decap_8 FILLER_50_1638 ();
 sg13g2_decap_4 FILLER_50_1645 ();
 sg13g2_fill_2 FILLER_50_1663 ();
 sg13g2_fill_1 FILLER_50_1665 ();
 sg13g2_decap_4 FILLER_50_1680 ();
 sg13g2_fill_2 FILLER_50_1689 ();
 sg13g2_fill_2 FILLER_50_1709 ();
 sg13g2_fill_2 FILLER_50_1729 ();
 sg13g2_fill_1 FILLER_50_1731 ();
 sg13g2_fill_1 FILLER_50_1742 ();
 sg13g2_fill_1 FILLER_50_1752 ();
 sg13g2_decap_8 FILLER_50_1761 ();
 sg13g2_decap_4 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_4 ();
 sg13g2_fill_2 FILLER_51_33 ();
 sg13g2_fill_2 FILLER_51_62 ();
 sg13g2_decap_8 FILLER_51_73 ();
 sg13g2_fill_2 FILLER_51_157 ();
 sg13g2_fill_1 FILLER_51_172 ();
 sg13g2_fill_2 FILLER_51_192 ();
 sg13g2_fill_1 FILLER_51_202 ();
 sg13g2_fill_1 FILLER_51_261 ();
 sg13g2_fill_2 FILLER_51_326 ();
 sg13g2_fill_2 FILLER_51_350 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_fill_2 FILLER_51_382 ();
 sg13g2_fill_1 FILLER_51_388 ();
 sg13g2_fill_2 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_51_413 ();
 sg13g2_decap_8 FILLER_51_420 ();
 sg13g2_fill_2 FILLER_51_427 ();
 sg13g2_fill_1 FILLER_51_437 ();
 sg13g2_fill_2 FILLER_51_461 ();
 sg13g2_fill_1 FILLER_51_468 ();
 sg13g2_decap_8 FILLER_51_474 ();
 sg13g2_fill_2 FILLER_51_481 ();
 sg13g2_fill_1 FILLER_51_523 ();
 sg13g2_fill_1 FILLER_51_578 ();
 sg13g2_fill_2 FILLER_51_604 ();
 sg13g2_fill_2 FILLER_51_609 ();
 sg13g2_fill_1 FILLER_51_611 ();
 sg13g2_decap_8 FILLER_51_641 ();
 sg13g2_fill_2 FILLER_51_648 ();
 sg13g2_fill_1 FILLER_51_660 ();
 sg13g2_fill_1 FILLER_51_697 ();
 sg13g2_decap_4 FILLER_51_704 ();
 sg13g2_fill_1 FILLER_51_708 ();
 sg13g2_decap_4 FILLER_51_746 ();
 sg13g2_fill_1 FILLER_51_750 ();
 sg13g2_fill_2 FILLER_51_756 ();
 sg13g2_fill_1 FILLER_51_762 ();
 sg13g2_fill_1 FILLER_51_781 ();
 sg13g2_fill_2 FILLER_51_828 ();
 sg13g2_fill_1 FILLER_51_830 ();
 sg13g2_fill_2 FILLER_51_868 ();
 sg13g2_fill_1 FILLER_51_876 ();
 sg13g2_decap_8 FILLER_51_881 ();
 sg13g2_fill_2 FILLER_51_888 ();
 sg13g2_decap_4 FILLER_51_924 ();
 sg13g2_fill_2 FILLER_51_928 ();
 sg13g2_fill_1 FILLER_51_934 ();
 sg13g2_fill_2 FILLER_51_952 ();
 sg13g2_fill_1 FILLER_51_954 ();
 sg13g2_fill_2 FILLER_51_1013 ();
 sg13g2_fill_1 FILLER_51_1015 ();
 sg13g2_fill_2 FILLER_51_1042 ();
 sg13g2_fill_2 FILLER_51_1085 ();
 sg13g2_fill_1 FILLER_51_1087 ();
 sg13g2_fill_1 FILLER_51_1121 ();
 sg13g2_fill_2 FILLER_51_1155 ();
 sg13g2_fill_2 FILLER_51_1172 ();
 sg13g2_fill_1 FILLER_51_1174 ();
 sg13g2_decap_4 FILLER_51_1248 ();
 sg13g2_fill_1 FILLER_51_1252 ();
 sg13g2_decap_8 FILLER_51_1280 ();
 sg13g2_decap_8 FILLER_51_1287 ();
 sg13g2_decap_4 FILLER_51_1294 ();
 sg13g2_fill_1 FILLER_51_1298 ();
 sg13g2_fill_2 FILLER_51_1308 ();
 sg13g2_fill_1 FILLER_51_1310 ();
 sg13g2_decap_8 FILLER_51_1321 ();
 sg13g2_fill_1 FILLER_51_1328 ();
 sg13g2_decap_8 FILLER_51_1349 ();
 sg13g2_fill_2 FILLER_51_1356 ();
 sg13g2_fill_1 FILLER_51_1363 ();
 sg13g2_decap_4 FILLER_51_1374 ();
 sg13g2_fill_2 FILLER_51_1378 ();
 sg13g2_fill_2 FILLER_51_1412 ();
 sg13g2_fill_1 FILLER_51_1414 ();
 sg13g2_fill_2 FILLER_51_1429 ();
 sg13g2_decap_4 FILLER_51_1446 ();
 sg13g2_fill_2 FILLER_51_1450 ();
 sg13g2_decap_4 FILLER_51_1461 ();
 sg13g2_fill_1 FILLER_51_1465 ();
 sg13g2_fill_1 FILLER_51_1477 ();
 sg13g2_decap_8 FILLER_51_1495 ();
 sg13g2_decap_8 FILLER_51_1531 ();
 sg13g2_fill_2 FILLER_51_1548 ();
 sg13g2_fill_1 FILLER_51_1550 ();
 sg13g2_decap_8 FILLER_51_1559 ();
 sg13g2_decap_4 FILLER_51_1566 ();
 sg13g2_fill_2 FILLER_51_1570 ();
 sg13g2_fill_2 FILLER_51_1583 ();
 sg13g2_fill_1 FILLER_51_1612 ();
 sg13g2_fill_1 FILLER_51_1622 ();
 sg13g2_decap_8 FILLER_51_1628 ();
 sg13g2_decap_8 FILLER_51_1635 ();
 sg13g2_fill_1 FILLER_51_1642 ();
 sg13g2_fill_2 FILLER_51_1661 ();
 sg13g2_fill_2 FILLER_51_1672 ();
 sg13g2_decap_8 FILLER_51_1679 ();
 sg13g2_fill_2 FILLER_51_1686 ();
 sg13g2_fill_1 FILLER_51_1688 ();
 sg13g2_decap_8 FILLER_51_1693 ();
 sg13g2_fill_2 FILLER_51_1700 ();
 sg13g2_fill_1 FILLER_51_1705 ();
 sg13g2_fill_2 FILLER_51_1712 ();
 sg13g2_fill_1 FILLER_51_1723 ();
 sg13g2_decap_4 FILLER_51_1730 ();
 sg13g2_fill_2 FILLER_51_1734 ();
 sg13g2_fill_2 FILLER_51_1745 ();
 sg13g2_fill_1 FILLER_51_1747 ();
 sg13g2_decap_8 FILLER_51_1756 ();
 sg13g2_decap_4 FILLER_51_1763 ();
 sg13g2_fill_1 FILLER_51_1767 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_107 ();
 sg13g2_fill_2 FILLER_52_143 ();
 sg13g2_fill_1 FILLER_52_145 ();
 sg13g2_fill_1 FILLER_52_190 ();
 sg13g2_decap_4 FILLER_52_196 ();
 sg13g2_decap_8 FILLER_52_204 ();
 sg13g2_fill_2 FILLER_52_211 ();
 sg13g2_fill_1 FILLER_52_213 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_fill_2 FILLER_52_242 ();
 sg13g2_fill_2 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_323 ();
 sg13g2_decap_4 FILLER_52_337 ();
 sg13g2_decap_4 FILLER_52_359 ();
 sg13g2_fill_2 FILLER_52_363 ();
 sg13g2_decap_4 FILLER_52_392 ();
 sg13g2_decap_4 FILLER_52_399 ();
 sg13g2_fill_1 FILLER_52_403 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_fill_1 FILLER_52_415 ();
 sg13g2_fill_1 FILLER_52_435 ();
 sg13g2_fill_2 FILLER_52_445 ();
 sg13g2_fill_2 FILLER_52_459 ();
 sg13g2_fill_2 FILLER_52_466 ();
 sg13g2_fill_1 FILLER_52_468 ();
 sg13g2_decap_8 FILLER_52_540 ();
 sg13g2_fill_2 FILLER_52_547 ();
 sg13g2_fill_1 FILLER_52_549 ();
 sg13g2_fill_1 FILLER_52_558 ();
 sg13g2_fill_2 FILLER_52_580 ();
 sg13g2_fill_1 FILLER_52_582 ();
 sg13g2_fill_1 FILLER_52_601 ();
 sg13g2_decap_8 FILLER_52_606 ();
 sg13g2_decap_8 FILLER_52_637 ();
 sg13g2_fill_1 FILLER_52_644 ();
 sg13g2_decap_8 FILLER_52_650 ();
 sg13g2_decap_8 FILLER_52_657 ();
 sg13g2_decap_8 FILLER_52_664 ();
 sg13g2_fill_1 FILLER_52_671 ();
 sg13g2_decap_4 FILLER_52_693 ();
 sg13g2_fill_2 FILLER_52_697 ();
 sg13g2_fill_2 FILLER_52_712 ();
 sg13g2_fill_1 FILLER_52_714 ();
 sg13g2_fill_1 FILLER_52_728 ();
 sg13g2_fill_1 FILLER_52_742 ();
 sg13g2_fill_1 FILLER_52_793 ();
 sg13g2_fill_2 FILLER_52_808 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_fill_1 FILLER_52_841 ();
 sg13g2_fill_2 FILLER_52_856 ();
 sg13g2_fill_1 FILLER_52_858 ();
 sg13g2_decap_8 FILLER_52_906 ();
 sg13g2_fill_2 FILLER_52_913 ();
 sg13g2_fill_1 FILLER_52_915 ();
 sg13g2_fill_1 FILLER_52_979 ();
 sg13g2_fill_2 FILLER_52_1008 ();
 sg13g2_fill_1 FILLER_52_1087 ();
 sg13g2_decap_4 FILLER_52_1110 ();
 sg13g2_decap_8 FILLER_52_1158 ();
 sg13g2_decap_8 FILLER_52_1165 ();
 sg13g2_fill_1 FILLER_52_1172 ();
 sg13g2_fill_2 FILLER_52_1206 ();
 sg13g2_fill_1 FILLER_52_1208 ();
 sg13g2_fill_1 FILLER_52_1267 ();
 sg13g2_decap_8 FILLER_52_1287 ();
 sg13g2_decap_8 FILLER_52_1294 ();
 sg13g2_decap_4 FILLER_52_1301 ();
 sg13g2_decap_4 FILLER_52_1326 ();
 sg13g2_fill_2 FILLER_52_1330 ();
 sg13g2_decap_8 FILLER_52_1352 ();
 sg13g2_fill_2 FILLER_52_1359 ();
 sg13g2_fill_1 FILLER_52_1391 ();
 sg13g2_decap_8 FILLER_52_1407 ();
 sg13g2_fill_2 FILLER_52_1414 ();
 sg13g2_fill_1 FILLER_52_1416 ();
 sg13g2_fill_2 FILLER_52_1421 ();
 sg13g2_fill_1 FILLER_52_1433 ();
 sg13g2_decap_8 FILLER_52_1438 ();
 sg13g2_fill_1 FILLER_52_1445 ();
 sg13g2_decap_8 FILLER_52_1459 ();
 sg13g2_decap_4 FILLER_52_1466 ();
 sg13g2_fill_2 FILLER_52_1470 ();
 sg13g2_decap_4 FILLER_52_1482 ();
 sg13g2_fill_2 FILLER_52_1486 ();
 sg13g2_decap_8 FILLER_52_1491 ();
 sg13g2_fill_2 FILLER_52_1498 ();
 sg13g2_fill_1 FILLER_52_1510 ();
 sg13g2_decap_8 FILLER_52_1518 ();
 sg13g2_fill_2 FILLER_52_1525 ();
 sg13g2_fill_1 FILLER_52_1540 ();
 sg13g2_fill_2 FILLER_52_1562 ();
 sg13g2_fill_1 FILLER_52_1564 ();
 sg13g2_fill_1 FILLER_52_1591 ();
 sg13g2_decap_8 FILLER_52_1596 ();
 sg13g2_decap_4 FILLER_52_1603 ();
 sg13g2_fill_2 FILLER_52_1607 ();
 sg13g2_fill_1 FILLER_52_1621 ();
 sg13g2_fill_2 FILLER_52_1626 ();
 sg13g2_fill_1 FILLER_52_1628 ();
 sg13g2_fill_1 FILLER_52_1637 ();
 sg13g2_decap_4 FILLER_52_1647 ();
 sg13g2_fill_1 FILLER_52_1655 ();
 sg13g2_decap_8 FILLER_52_1661 ();
 sg13g2_fill_2 FILLER_52_1668 ();
 sg13g2_fill_1 FILLER_52_1670 ();
 sg13g2_fill_1 FILLER_52_1676 ();
 sg13g2_fill_2 FILLER_52_1704 ();
 sg13g2_fill_1 FILLER_52_1706 ();
 sg13g2_decap_4 FILLER_52_1762 ();
 sg13g2_fill_2 FILLER_52_1766 ();
 sg13g2_fill_1 FILLER_53_27 ();
 sg13g2_fill_2 FILLER_53_37 ();
 sg13g2_fill_2 FILLER_53_63 ();
 sg13g2_fill_1 FILLER_53_65 ();
 sg13g2_decap_8 FILLER_53_78 ();
 sg13g2_fill_1 FILLER_53_85 ();
 sg13g2_fill_2 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_1 FILLER_53_179 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_2 FILLER_53_249 ();
 sg13g2_fill_1 FILLER_53_251 ();
 sg13g2_fill_1 FILLER_53_261 ();
 sg13g2_fill_1 FILLER_53_271 ();
 sg13g2_decap_4 FILLER_53_280 ();
 sg13g2_fill_2 FILLER_53_284 ();
 sg13g2_decap_4 FILLER_53_323 ();
 sg13g2_decap_8 FILLER_53_337 ();
 sg13g2_fill_2 FILLER_53_361 ();
 sg13g2_fill_2 FILLER_53_370 ();
 sg13g2_fill_1 FILLER_53_372 ();
 sg13g2_decap_8 FILLER_53_391 ();
 sg13g2_fill_1 FILLER_53_398 ();
 sg13g2_decap_8 FILLER_53_435 ();
 sg13g2_fill_1 FILLER_53_442 ();
 sg13g2_fill_2 FILLER_53_454 ();
 sg13g2_fill_1 FILLER_53_476 ();
 sg13g2_fill_2 FILLER_53_488 ();
 sg13g2_fill_2 FILLER_53_541 ();
 sg13g2_fill_1 FILLER_53_543 ();
 sg13g2_fill_1 FILLER_53_553 ();
 sg13g2_decap_8 FILLER_53_566 ();
 sg13g2_decap_4 FILLER_53_627 ();
 sg13g2_fill_1 FILLER_53_631 ();
 sg13g2_decap_4 FILLER_53_642 ();
 sg13g2_fill_2 FILLER_53_656 ();
 sg13g2_fill_1 FILLER_53_663 ();
 sg13g2_fill_2 FILLER_53_686 ();
 sg13g2_fill_2 FILLER_53_708 ();
 sg13g2_fill_1 FILLER_53_752 ();
 sg13g2_fill_2 FILLER_53_794 ();
 sg13g2_decap_8 FILLER_53_829 ();
 sg13g2_fill_2 FILLER_53_836 ();
 sg13g2_decap_4 FILLER_53_851 ();
 sg13g2_fill_1 FILLER_53_855 ();
 sg13g2_fill_1 FILLER_53_888 ();
 sg13g2_decap_4 FILLER_53_902 ();
 sg13g2_fill_2 FILLER_53_906 ();
 sg13g2_fill_2 FILLER_53_918 ();
 sg13g2_fill_2 FILLER_53_935 ();
 sg13g2_fill_1 FILLER_53_937 ();
 sg13g2_fill_2 FILLER_53_966 ();
 sg13g2_fill_1 FILLER_53_987 ();
 sg13g2_fill_1 FILLER_53_1029 ();
 sg13g2_fill_2 FILLER_53_1039 ();
 sg13g2_fill_1 FILLER_53_1091 ();
 sg13g2_fill_2 FILLER_53_1141 ();
 sg13g2_fill_1 FILLER_53_1143 ();
 sg13g2_fill_2 FILLER_53_1185 ();
 sg13g2_fill_2 FILLER_53_1206 ();
 sg13g2_fill_1 FILLER_53_1214 ();
 sg13g2_fill_1 FILLER_53_1223 ();
 sg13g2_fill_1 FILLER_53_1298 ();
 sg13g2_decap_8 FILLER_53_1373 ();
 sg13g2_decap_8 FILLER_53_1380 ();
 sg13g2_fill_1 FILLER_53_1387 ();
 sg13g2_fill_1 FILLER_53_1398 ();
 sg13g2_fill_2 FILLER_53_1412 ();
 sg13g2_fill_1 FILLER_53_1414 ();
 sg13g2_decap_8 FILLER_53_1461 ();
 sg13g2_fill_1 FILLER_53_1468 ();
 sg13g2_decap_4 FILLER_53_1494 ();
 sg13g2_decap_8 FILLER_53_1518 ();
 sg13g2_fill_2 FILLER_53_1525 ();
 sg13g2_decap_4 FILLER_53_1540 ();
 sg13g2_fill_2 FILLER_53_1557 ();
 sg13g2_fill_1 FILLER_53_1559 ();
 sg13g2_fill_2 FILLER_53_1568 ();
 sg13g2_decap_8 FILLER_53_1588 ();
 sg13g2_decap_8 FILLER_53_1595 ();
 sg13g2_decap_8 FILLER_53_1625 ();
 sg13g2_fill_2 FILLER_53_1632 ();
 sg13g2_fill_1 FILLER_53_1634 ();
 sg13g2_decap_4 FILLER_53_1643 ();
 sg13g2_fill_2 FILLER_53_1661 ();
 sg13g2_decap_8 FILLER_53_1681 ();
 sg13g2_fill_2 FILLER_53_1688 ();
 sg13g2_fill_1 FILLER_53_1690 ();
 sg13g2_decap_4 FILLER_53_1713 ();
 sg13g2_fill_2 FILLER_53_1717 ();
 sg13g2_decap_8 FILLER_53_1728 ();
 sg13g2_decap_8 FILLER_53_1754 ();
 sg13g2_decap_8 FILLER_53_1761 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_4 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_46 ();
 sg13g2_fill_2 FILLER_54_57 ();
 sg13g2_decap_8 FILLER_54_84 ();
 sg13g2_fill_2 FILLER_54_91 ();
 sg13g2_fill_2 FILLER_54_120 ();
 sg13g2_fill_1 FILLER_54_122 ();
 sg13g2_decap_4 FILLER_54_140 ();
 sg13g2_fill_2 FILLER_54_149 ();
 sg13g2_fill_1 FILLER_54_192 ();
 sg13g2_decap_8 FILLER_54_199 ();
 sg13g2_decap_8 FILLER_54_206 ();
 sg13g2_decap_8 FILLER_54_213 ();
 sg13g2_decap_4 FILLER_54_220 ();
 sg13g2_fill_1 FILLER_54_224 ();
 sg13g2_fill_1 FILLER_54_237 ();
 sg13g2_decap_8 FILLER_54_282 ();
 sg13g2_decap_4 FILLER_54_289 ();
 sg13g2_fill_2 FILLER_54_293 ();
 sg13g2_fill_2 FILLER_54_299 ();
 sg13g2_fill_2 FILLER_54_305 ();
 sg13g2_fill_1 FILLER_54_307 ();
 sg13g2_fill_2 FILLER_54_312 ();
 sg13g2_decap_8 FILLER_54_322 ();
 sg13g2_fill_1 FILLER_54_329 ();
 sg13g2_fill_2 FILLER_54_358 ();
 sg13g2_fill_1 FILLER_54_364 ();
 sg13g2_fill_2 FILLER_54_427 ();
 sg13g2_fill_2 FILLER_54_462 ();
 sg13g2_fill_1 FILLER_54_464 ();
 sg13g2_decap_4 FILLER_54_497 ();
 sg13g2_decap_8 FILLER_54_524 ();
 sg13g2_fill_1 FILLER_54_531 ();
 sg13g2_decap_8 FILLER_54_544 ();
 sg13g2_fill_1 FILLER_54_551 ();
 sg13g2_fill_2 FILLER_54_574 ();
 sg13g2_fill_1 FILLER_54_589 ();
 sg13g2_decap_4 FILLER_54_604 ();
 sg13g2_fill_1 FILLER_54_608 ();
 sg13g2_decap_4 FILLER_54_639 ();
 sg13g2_decap_4 FILLER_54_658 ();
 sg13g2_fill_1 FILLER_54_693 ();
 sg13g2_fill_1 FILLER_54_705 ();
 sg13g2_fill_1 FILLER_54_711 ();
 sg13g2_fill_1 FILLER_54_778 ();
 sg13g2_fill_2 FILLER_54_784 ();
 sg13g2_fill_1 FILLER_54_822 ();
 sg13g2_decap_4 FILLER_54_855 ();
 sg13g2_fill_2 FILLER_54_859 ();
 sg13g2_decap_8 FILLER_54_865 ();
 sg13g2_decap_4 FILLER_54_872 ();
 sg13g2_fill_1 FILLER_54_876 ();
 sg13g2_decap_8 FILLER_54_883 ();
 sg13g2_decap_8 FILLER_54_890 ();
 sg13g2_decap_4 FILLER_54_897 ();
 sg13g2_fill_2 FILLER_54_901 ();
 sg13g2_fill_2 FILLER_54_1021 ();
 sg13g2_fill_2 FILLER_54_1051 ();
 sg13g2_fill_1 FILLER_54_1053 ();
 sg13g2_fill_1 FILLER_54_1072 ();
 sg13g2_fill_1 FILLER_54_1095 ();
 sg13g2_decap_4 FILLER_54_1142 ();
 sg13g2_decap_8 FILLER_54_1155 ();
 sg13g2_decap_8 FILLER_54_1162 ();
 sg13g2_fill_2 FILLER_54_1169 ();
 sg13g2_fill_1 FILLER_54_1171 ();
 sg13g2_fill_2 FILLER_54_1189 ();
 sg13g2_fill_1 FILLER_54_1191 ();
 sg13g2_fill_2 FILLER_54_1207 ();
 sg13g2_fill_1 FILLER_54_1209 ();
 sg13g2_fill_2 FILLER_54_1219 ();
 sg13g2_fill_2 FILLER_54_1239 ();
 sg13g2_fill_1 FILLER_54_1241 ();
 sg13g2_decap_8 FILLER_54_1291 ();
 sg13g2_decap_8 FILLER_54_1298 ();
 sg13g2_fill_1 FILLER_54_1305 ();
 sg13g2_fill_2 FILLER_54_1324 ();
 sg13g2_fill_1 FILLER_54_1326 ();
 sg13g2_fill_1 FILLER_54_1331 ();
 sg13g2_decap_8 FILLER_54_1336 ();
 sg13g2_fill_2 FILLER_54_1343 ();
 sg13g2_decap_8 FILLER_54_1355 ();
 sg13g2_decap_8 FILLER_54_1376 ();
 sg13g2_decap_4 FILLER_54_1383 ();
 sg13g2_decap_8 FILLER_54_1409 ();
 sg13g2_decap_4 FILLER_54_1416 ();
 sg13g2_fill_1 FILLER_54_1420 ();
 sg13g2_decap_4 FILLER_54_1439 ();
 sg13g2_decap_8 FILLER_54_1456 ();
 sg13g2_fill_2 FILLER_54_1463 ();
 sg13g2_decap_4 FILLER_54_1485 ();
 sg13g2_decap_4 FILLER_54_1493 ();
 sg13g2_decap_4 FILLER_54_1513 ();
 sg13g2_fill_2 FILLER_54_1517 ();
 sg13g2_decap_4 FILLER_54_1553 ();
 sg13g2_fill_1 FILLER_54_1557 ();
 sg13g2_decap_4 FILLER_54_1562 ();
 sg13g2_fill_2 FILLER_54_1566 ();
 sg13g2_decap_4 FILLER_54_1573 ();
 sg13g2_decap_4 FILLER_54_1580 ();
 sg13g2_fill_2 FILLER_54_1584 ();
 sg13g2_fill_2 FILLER_54_1606 ();
 sg13g2_fill_1 FILLER_54_1608 ();
 sg13g2_decap_8 FILLER_54_1616 ();
 sg13g2_decap_4 FILLER_54_1623 ();
 sg13g2_fill_1 FILLER_54_1627 ();
 sg13g2_decap_4 FILLER_54_1647 ();
 sg13g2_fill_1 FILLER_54_1651 ();
 sg13g2_decap_4 FILLER_54_1660 ();
 sg13g2_fill_1 FILLER_54_1664 ();
 sg13g2_fill_2 FILLER_54_1678 ();
 sg13g2_decap_8 FILLER_54_1710 ();
 sg13g2_fill_2 FILLER_54_1717 ();
 sg13g2_fill_1 FILLER_54_1719 ();
 sg13g2_fill_1 FILLER_54_1725 ();
 sg13g2_fill_1 FILLER_54_1739 ();
 sg13g2_fill_1 FILLER_54_1745 ();
 sg13g2_decap_8 FILLER_54_1759 ();
 sg13g2_fill_2 FILLER_54_1766 ();
 sg13g2_decap_4 FILLER_55_0 ();
 sg13g2_fill_1 FILLER_55_4 ();
 sg13g2_decap_8 FILLER_55_9 ();
 sg13g2_decap_8 FILLER_55_16 ();
 sg13g2_fill_2 FILLER_55_37 ();
 sg13g2_fill_2 FILLER_55_102 ();
 sg13g2_decap_8 FILLER_55_108 ();
 sg13g2_decap_4 FILLER_55_115 ();
 sg13g2_fill_2 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_153 ();
 sg13g2_fill_1 FILLER_55_155 ();
 sg13g2_fill_1 FILLER_55_179 ();
 sg13g2_fill_2 FILLER_55_189 ();
 sg13g2_fill_1 FILLER_55_191 ();
 sg13g2_decap_8 FILLER_55_225 ();
 sg13g2_decap_4 FILLER_55_232 ();
 sg13g2_fill_1 FILLER_55_236 ();
 sg13g2_fill_2 FILLER_55_242 ();
 sg13g2_decap_8 FILLER_55_257 ();
 sg13g2_fill_1 FILLER_55_264 ();
 sg13g2_fill_1 FILLER_55_346 ();
 sg13g2_fill_2 FILLER_55_358 ();
 sg13g2_fill_2 FILLER_55_378 ();
 sg13g2_fill_1 FILLER_55_380 ();
 sg13g2_fill_1 FILLER_55_412 ();
 sg13g2_decap_4 FILLER_55_459 ();
 sg13g2_fill_1 FILLER_55_491 ();
 sg13g2_fill_2 FILLER_55_522 ();
 sg13g2_fill_2 FILLER_55_541 ();
 sg13g2_decap_4 FILLER_55_572 ();
 sg13g2_decap_4 FILLER_55_616 ();
 sg13g2_fill_1 FILLER_55_620 ();
 sg13g2_decap_4 FILLER_55_630 ();
 sg13g2_fill_2 FILLER_55_634 ();
 sg13g2_fill_1 FILLER_55_660 ();
 sg13g2_fill_2 FILLER_55_684 ();
 sg13g2_fill_2 FILLER_55_702 ();
 sg13g2_fill_1 FILLER_55_704 ();
 sg13g2_decap_4 FILLER_55_724 ();
 sg13g2_fill_1 FILLER_55_767 ();
 sg13g2_fill_1 FILLER_55_813 ();
 sg13g2_fill_1 FILLER_55_878 ();
 sg13g2_decap_8 FILLER_55_911 ();
 sg13g2_decap_4 FILLER_55_918 ();
 sg13g2_fill_2 FILLER_55_985 ();
 sg13g2_fill_2 FILLER_55_1006 ();
 sg13g2_fill_2 FILLER_55_1017 ();
 sg13g2_fill_1 FILLER_55_1019 ();
 sg13g2_fill_1 FILLER_55_1057 ();
 sg13g2_fill_1 FILLER_55_1099 ();
 sg13g2_fill_1 FILLER_55_1122 ();
 sg13g2_fill_2 FILLER_55_1127 ();
 sg13g2_fill_1 FILLER_55_1129 ();
 sg13g2_decap_4 FILLER_55_1154 ();
 sg13g2_fill_2 FILLER_55_1158 ();
 sg13g2_decap_8 FILLER_55_1173 ();
 sg13g2_fill_2 FILLER_55_1180 ();
 sg13g2_fill_2 FILLER_55_1188 ();
 sg13g2_fill_1 FILLER_55_1242 ();
 sg13g2_fill_1 FILLER_55_1254 ();
 sg13g2_decap_8 FILLER_55_1301 ();
 sg13g2_decap_8 FILLER_55_1308 ();
 sg13g2_fill_1 FILLER_55_1315 ();
 sg13g2_fill_1 FILLER_55_1324 ();
 sg13g2_fill_2 FILLER_55_1362 ();
 sg13g2_fill_1 FILLER_55_1364 ();
 sg13g2_fill_2 FILLER_55_1378 ();
 sg13g2_fill_1 FILLER_55_1380 ();
 sg13g2_decap_8 FILLER_55_1408 ();
 sg13g2_fill_2 FILLER_55_1415 ();
 sg13g2_fill_2 FILLER_55_1427 ();
 sg13g2_fill_2 FILLER_55_1433 ();
 sg13g2_fill_1 FILLER_55_1435 ();
 sg13g2_decap_4 FILLER_55_1453 ();
 sg13g2_decap_4 FILLER_55_1460 ();
 sg13g2_fill_1 FILLER_55_1464 ();
 sg13g2_decap_4 FILLER_55_1483 ();
 sg13g2_fill_1 FILLER_55_1487 ();
 sg13g2_decap_4 FILLER_55_1495 ();
 sg13g2_decap_8 FILLER_55_1512 ();
 sg13g2_fill_1 FILLER_55_1519 ();
 sg13g2_decap_4 FILLER_55_1541 ();
 sg13g2_fill_1 FILLER_55_1550 ();
 sg13g2_decap_8 FILLER_55_1555 ();
 sg13g2_fill_2 FILLER_55_1562 ();
 sg13g2_fill_1 FILLER_55_1564 ();
 sg13g2_decap_8 FILLER_55_1573 ();
 sg13g2_decap_4 FILLER_55_1580 ();
 sg13g2_fill_1 FILLER_55_1584 ();
 sg13g2_decap_4 FILLER_55_1607 ();
 sg13g2_fill_1 FILLER_55_1611 ();
 sg13g2_decap_8 FILLER_55_1633 ();
 sg13g2_fill_1 FILLER_55_1657 ();
 sg13g2_fill_2 FILLER_55_1663 ();
 sg13g2_fill_1 FILLER_55_1682 ();
 sg13g2_decap_8 FILLER_55_1688 ();
 sg13g2_fill_1 FILLER_55_1695 ();
 sg13g2_fill_2 FILLER_55_1706 ();
 sg13g2_fill_1 FILLER_55_1708 ();
 sg13g2_fill_2 FILLER_55_1714 ();
 sg13g2_decap_4 FILLER_55_1739 ();
 sg13g2_decap_8 FILLER_55_1760 ();
 sg13g2_fill_1 FILLER_55_1767 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_15 ();
 sg13g2_fill_2 FILLER_56_22 ();
 sg13g2_fill_1 FILLER_56_24 ();
 sg13g2_fill_2 FILLER_56_61 ();
 sg13g2_fill_1 FILLER_56_63 ();
 sg13g2_decap_8 FILLER_56_85 ();
 sg13g2_decap_8 FILLER_56_92 ();
 sg13g2_fill_2 FILLER_56_99 ();
 sg13g2_fill_1 FILLER_56_101 ();
 sg13g2_decap_8 FILLER_56_130 ();
 sg13g2_fill_1 FILLER_56_159 ();
 sg13g2_fill_2 FILLER_56_166 ();
 sg13g2_fill_1 FILLER_56_168 ();
 sg13g2_decap_8 FILLER_56_181 ();
 sg13g2_fill_1 FILLER_56_192 ();
 sg13g2_fill_2 FILLER_56_203 ();
 sg13g2_fill_1 FILLER_56_222 ();
 sg13g2_decap_8 FILLER_56_257 ();
 sg13g2_fill_2 FILLER_56_280 ();
 sg13g2_fill_1 FILLER_56_282 ();
 sg13g2_fill_2 FILLER_56_289 ();
 sg13g2_decap_8 FILLER_56_309 ();
 sg13g2_decap_4 FILLER_56_329 ();
 sg13g2_fill_2 FILLER_56_349 ();
 sg13g2_fill_1 FILLER_56_351 ();
 sg13g2_fill_2 FILLER_56_389 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_decap_8 FILLER_56_515 ();
 sg13g2_decap_8 FILLER_56_535 ();
 sg13g2_decap_4 FILLER_56_542 ();
 sg13g2_fill_1 FILLER_56_546 ();
 sg13g2_fill_2 FILLER_56_568 ();
 sg13g2_decap_4 FILLER_56_574 ();
 sg13g2_fill_1 FILLER_56_578 ();
 sg13g2_fill_2 FILLER_56_584 ();
 sg13g2_fill_1 FILLER_56_586 ();
 sg13g2_fill_2 FILLER_56_626 ();
 sg13g2_fill_1 FILLER_56_628 ();
 sg13g2_fill_2 FILLER_56_647 ();
 sg13g2_fill_2 FILLER_56_654 ();
 sg13g2_fill_2 FILLER_56_671 ();
 sg13g2_fill_1 FILLER_56_673 ();
 sg13g2_fill_1 FILLER_56_679 ();
 sg13g2_decap_4 FILLER_56_693 ();
 sg13g2_fill_2 FILLER_56_697 ();
 sg13g2_fill_2 FILLER_56_723 ();
 sg13g2_fill_1 FILLER_56_725 ();
 sg13g2_fill_2 FILLER_56_782 ();
 sg13g2_fill_1 FILLER_56_784 ();
 sg13g2_fill_1 FILLER_56_794 ();
 sg13g2_fill_2 FILLER_56_808 ();
 sg13g2_fill_1 FILLER_56_810 ();
 sg13g2_fill_2 FILLER_56_842 ();
 sg13g2_decap_4 FILLER_56_870 ();
 sg13g2_fill_1 FILLER_56_874 ();
 sg13g2_fill_1 FILLER_56_899 ();
 sg13g2_fill_2 FILLER_56_936 ();
 sg13g2_fill_2 FILLER_56_972 ();
 sg13g2_fill_1 FILLER_56_974 ();
 sg13g2_fill_2 FILLER_56_993 ();
 sg13g2_fill_2 FILLER_56_1067 ();
 sg13g2_fill_2 FILLER_56_1078 ();
 sg13g2_fill_1 FILLER_56_1089 ();
 sg13g2_fill_1 FILLER_56_1110 ();
 sg13g2_decap_4 FILLER_56_1151 ();
 sg13g2_fill_2 FILLER_56_1187 ();
 sg13g2_fill_1 FILLER_56_1189 ();
 sg13g2_decap_8 FILLER_56_1194 ();
 sg13g2_decap_8 FILLER_56_1201 ();
 sg13g2_fill_1 FILLER_56_1208 ();
 sg13g2_fill_2 FILLER_56_1227 ();
 sg13g2_fill_1 FILLER_56_1276 ();
 sg13g2_fill_2 FILLER_56_1308 ();
 sg13g2_decap_4 FILLER_56_1336 ();
 sg13g2_fill_1 FILLER_56_1340 ();
 sg13g2_decap_8 FILLER_56_1350 ();
 sg13g2_decap_4 FILLER_56_1357 ();
 sg13g2_fill_2 FILLER_56_1361 ();
 sg13g2_fill_1 FILLER_56_1373 ();
 sg13g2_decap_8 FILLER_56_1379 ();
 sg13g2_decap_4 FILLER_56_1386 ();
 sg13g2_fill_1 FILLER_56_1390 ();
 sg13g2_fill_1 FILLER_56_1394 ();
 sg13g2_fill_2 FILLER_56_1399 ();
 sg13g2_fill_1 FILLER_56_1401 ();
 sg13g2_decap_8 FILLER_56_1429 ();
 sg13g2_fill_2 FILLER_56_1436 ();
 sg13g2_fill_1 FILLER_56_1438 ();
 sg13g2_fill_1 FILLER_56_1473 ();
 sg13g2_decap_8 FILLER_56_1478 ();
 sg13g2_fill_2 FILLER_56_1485 ();
 sg13g2_fill_1 FILLER_56_1487 ();
 sg13g2_fill_1 FILLER_56_1493 ();
 sg13g2_decap_8 FILLER_56_1511 ();
 sg13g2_fill_2 FILLER_56_1518 ();
 sg13g2_fill_1 FILLER_56_1520 ();
 sg13g2_fill_2 FILLER_56_1532 ();
 sg13g2_fill_2 FILLER_56_1551 ();
 sg13g2_fill_1 FILLER_56_1553 ();
 sg13g2_decap_4 FILLER_56_1571 ();
 sg13g2_fill_1 FILLER_56_1575 ();
 sg13g2_decap_4 FILLER_56_1589 ();
 sg13g2_fill_2 FILLER_56_1593 ();
 sg13g2_fill_1 FILLER_56_1608 ();
 sg13g2_fill_1 FILLER_56_1640 ();
 sg13g2_fill_1 FILLER_56_1646 ();
 sg13g2_fill_2 FILLER_56_1660 ();
 sg13g2_decap_4 FILLER_56_1680 ();
 sg13g2_fill_2 FILLER_56_1684 ();
 sg13g2_fill_2 FILLER_56_1698 ();
 sg13g2_decap_8 FILLER_56_1709 ();
 sg13g2_fill_1 FILLER_56_1716 ();
 sg13g2_decap_8 FILLER_56_1733 ();
 sg13g2_decap_4 FILLER_56_1762 ();
 sg13g2_fill_2 FILLER_56_1766 ();
 sg13g2_decap_4 FILLER_57_59 ();
 sg13g2_decap_4 FILLER_57_103 ();
 sg13g2_decap_8 FILLER_57_111 ();
 sg13g2_fill_2 FILLER_57_118 ();
 sg13g2_fill_2 FILLER_57_152 ();
 sg13g2_fill_1 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_178 ();
 sg13g2_fill_1 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_218 ();
 sg13g2_decap_8 FILLER_57_225 ();
 sg13g2_decap_4 FILLER_57_232 ();
 sg13g2_fill_2 FILLER_57_236 ();
 sg13g2_fill_2 FILLER_57_243 ();
 sg13g2_decap_8 FILLER_57_250 ();
 sg13g2_fill_1 FILLER_57_271 ();
 sg13g2_fill_1 FILLER_57_290 ();
 sg13g2_fill_2 FILLER_57_329 ();
 sg13g2_fill_1 FILLER_57_375 ();
 sg13g2_fill_1 FILLER_57_427 ();
 sg13g2_fill_1 FILLER_57_464 ();
 sg13g2_decap_8 FILLER_57_496 ();
 sg13g2_fill_2 FILLER_57_503 ();
 sg13g2_fill_2 FILLER_57_510 ();
 sg13g2_fill_2 FILLER_57_561 ();
 sg13g2_decap_4 FILLER_57_585 ();
 sg13g2_fill_2 FILLER_57_589 ();
 sg13g2_decap_8 FILLER_57_601 ();
 sg13g2_fill_2 FILLER_57_613 ();
 sg13g2_fill_1 FILLER_57_615 ();
 sg13g2_fill_2 FILLER_57_626 ();
 sg13g2_fill_2 FILLER_57_641 ();
 sg13g2_fill_1 FILLER_57_643 ();
 sg13g2_fill_1 FILLER_57_659 ();
 sg13g2_decap_8 FILLER_57_677 ();
 sg13g2_decap_8 FILLER_57_697 ();
 sg13g2_fill_2 FILLER_57_704 ();
 sg13g2_fill_2 FILLER_57_735 ();
 sg13g2_fill_2 FILLER_57_748 ();
 sg13g2_fill_1 FILLER_57_750 ();
 sg13g2_fill_2 FILLER_57_786 ();
 sg13g2_fill_1 FILLER_57_788 ();
 sg13g2_fill_2 FILLER_57_804 ();
 sg13g2_fill_1 FILLER_57_806 ();
 sg13g2_fill_2 FILLER_57_840 ();
 sg13g2_fill_2 FILLER_57_846 ();
 sg13g2_fill_2 FILLER_57_880 ();
 sg13g2_fill_2 FILLER_57_920 ();
 sg13g2_fill_1 FILLER_57_922 ();
 sg13g2_fill_2 FILLER_57_1004 ();
 sg13g2_fill_1 FILLER_57_1047 ();
 sg13g2_fill_1 FILLER_57_1067 ();
 sg13g2_fill_2 FILLER_57_1099 ();
 sg13g2_fill_2 FILLER_57_1142 ();
 sg13g2_fill_1 FILLER_57_1144 ();
 sg13g2_decap_4 FILLER_57_1163 ();
 sg13g2_fill_1 FILLER_57_1184 ();
 sg13g2_fill_1 FILLER_57_1204 ();
 sg13g2_fill_2 FILLER_57_1261 ();
 sg13g2_fill_1 FILLER_57_1276 ();
 sg13g2_fill_2 FILLER_57_1287 ();
 sg13g2_fill_1 FILLER_57_1289 ();
 sg13g2_fill_1 FILLER_57_1296 ();
 sg13g2_decap_8 FILLER_57_1305 ();
 sg13g2_fill_2 FILLER_57_1312 ();
 sg13g2_fill_1 FILLER_57_1314 ();
 sg13g2_decap_4 FILLER_57_1332 ();
 sg13g2_fill_2 FILLER_57_1341 ();
 sg13g2_fill_1 FILLER_57_1343 ();
 sg13g2_decap_8 FILLER_57_1349 ();
 sg13g2_fill_1 FILLER_57_1356 ();
 sg13g2_decap_8 FILLER_57_1385 ();
 sg13g2_fill_1 FILLER_57_1392 ();
 sg13g2_decap_8 FILLER_57_1411 ();
 sg13g2_fill_2 FILLER_57_1418 ();
 sg13g2_fill_1 FILLER_57_1420 ();
 sg13g2_decap_8 FILLER_57_1429 ();
 sg13g2_decap_4 FILLER_57_1436 ();
 sg13g2_fill_1 FILLER_57_1440 ();
 sg13g2_fill_1 FILLER_57_1445 ();
 sg13g2_decap_8 FILLER_57_1458 ();
 sg13g2_fill_1 FILLER_57_1465 ();
 sg13g2_decap_4 FILLER_57_1472 ();
 sg13g2_fill_2 FILLER_57_1484 ();
 sg13g2_fill_1 FILLER_57_1486 ();
 sg13g2_fill_2 FILLER_57_1492 ();
 sg13g2_fill_1 FILLER_57_1494 ();
 sg13g2_decap_4 FILLER_57_1500 ();
 sg13g2_fill_2 FILLER_57_1509 ();
 sg13g2_decap_8 FILLER_57_1516 ();
 sg13g2_decap_8 FILLER_57_1528 ();
 sg13g2_fill_2 FILLER_57_1535 ();
 sg13g2_decap_4 FILLER_57_1546 ();
 sg13g2_fill_1 FILLER_57_1550 ();
 sg13g2_fill_2 FILLER_57_1556 ();
 sg13g2_fill_2 FILLER_57_1572 ();
 sg13g2_fill_1 FILLER_57_1574 ();
 sg13g2_decap_4 FILLER_57_1578 ();
 sg13g2_fill_1 FILLER_57_1582 ();
 sg13g2_fill_1 FILLER_57_1587 ();
 sg13g2_decap_8 FILLER_57_1601 ();
 sg13g2_decap_4 FILLER_57_1608 ();
 sg13g2_fill_2 FILLER_57_1636 ();
 sg13g2_fill_1 FILLER_57_1638 ();
 sg13g2_fill_1 FILLER_57_1656 ();
 sg13g2_decap_8 FILLER_57_1680 ();
 sg13g2_fill_1 FILLER_57_1687 ();
 sg13g2_fill_2 FILLER_57_1710 ();
 sg13g2_fill_1 FILLER_57_1712 ();
 sg13g2_fill_2 FILLER_57_1718 ();
 sg13g2_decap_4 FILLER_57_1764 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_7 ();
 sg13g2_fill_2 FILLER_58_15 ();
 sg13g2_fill_1 FILLER_58_17 ();
 sg13g2_fill_2 FILLER_58_83 ();
 sg13g2_fill_2 FILLER_58_117 ();
 sg13g2_fill_1 FILLER_58_119 ();
 sg13g2_fill_2 FILLER_58_164 ();
 sg13g2_fill_1 FILLER_58_166 ();
 sg13g2_decap_4 FILLER_58_186 ();
 sg13g2_fill_1 FILLER_58_205 ();
 sg13g2_fill_1 FILLER_58_211 ();
 sg13g2_decap_8 FILLER_58_219 ();
 sg13g2_fill_1 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_271 ();
 sg13g2_decap_4 FILLER_58_285 ();
 sg13g2_fill_1 FILLER_58_310 ();
 sg13g2_decap_8 FILLER_58_362 ();
 sg13g2_fill_2 FILLER_58_369 ();
 sg13g2_fill_1 FILLER_58_388 ();
 sg13g2_fill_2 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_414 ();
 sg13g2_fill_2 FILLER_58_462 ();
 sg13g2_fill_2 FILLER_58_513 ();
 sg13g2_fill_1 FILLER_58_529 ();
 sg13g2_decap_4 FILLER_58_534 ();
 sg13g2_fill_2 FILLER_58_538 ();
 sg13g2_decap_4 FILLER_58_562 ();
 sg13g2_fill_1 FILLER_58_606 ();
 sg13g2_fill_2 FILLER_58_611 ();
 sg13g2_fill_1 FILLER_58_617 ();
 sg13g2_decap_4 FILLER_58_645 ();
 sg13g2_fill_2 FILLER_58_662 ();
 sg13g2_fill_1 FILLER_58_664 ();
 sg13g2_decap_4 FILLER_58_696 ();
 sg13g2_fill_1 FILLER_58_700 ();
 sg13g2_fill_1 FILLER_58_720 ();
 sg13g2_fill_2 FILLER_58_755 ();
 sg13g2_fill_2 FILLER_58_803 ();
 sg13g2_fill_1 FILLER_58_805 ();
 sg13g2_fill_2 FILLER_58_832 ();
 sg13g2_fill_2 FILLER_58_848 ();
 sg13g2_fill_2 FILLER_58_883 ();
 sg13g2_fill_1 FILLER_58_885 ();
 sg13g2_decap_4 FILLER_58_914 ();
 sg13g2_fill_1 FILLER_58_918 ();
 sg13g2_fill_1 FILLER_58_948 ();
 sg13g2_fill_2 FILLER_58_968 ();
 sg13g2_fill_2 FILLER_58_997 ();
 sg13g2_fill_1 FILLER_58_999 ();
 sg13g2_fill_2 FILLER_58_1086 ();
 sg13g2_fill_1 FILLER_58_1088 ();
 sg13g2_fill_1 FILLER_58_1098 ();
 sg13g2_decap_8 FILLER_58_1125 ();
 sg13g2_fill_1 FILLER_58_1132 ();
 sg13g2_fill_2 FILLER_58_1146 ();
 sg13g2_fill_1 FILLER_58_1148 ();
 sg13g2_fill_2 FILLER_58_1225 ();
 sg13g2_fill_2 FILLER_58_1245 ();
 sg13g2_fill_1 FILLER_58_1247 ();
 sg13g2_fill_1 FILLER_58_1276 ();
 sg13g2_decap_4 FILLER_58_1311 ();
 sg13g2_fill_1 FILLER_58_1315 ();
 sg13g2_decap_8 FILLER_58_1330 ();
 sg13g2_fill_1 FILLER_58_1337 ();
 sg13g2_decap_8 FILLER_58_1358 ();
 sg13g2_decap_4 FILLER_58_1365 ();
 sg13g2_decap_8 FILLER_58_1379 ();
 sg13g2_decap_4 FILLER_58_1386 ();
 sg13g2_fill_1 FILLER_58_1404 ();
 sg13g2_decap_4 FILLER_58_1413 ();
 sg13g2_decap_4 FILLER_58_1429 ();
 sg13g2_decap_4 FILLER_58_1454 ();
 sg13g2_fill_2 FILLER_58_1458 ();
 sg13g2_decap_4 FILLER_58_1471 ();
 sg13g2_decap_4 FILLER_58_1494 ();
 sg13g2_fill_2 FILLER_58_1522 ();
 sg13g2_decap_4 FILLER_58_1541 ();
 sg13g2_fill_2 FILLER_58_1545 ();
 sg13g2_fill_2 FILLER_58_1560 ();
 sg13g2_fill_1 FILLER_58_1577 ();
 sg13g2_decap_4 FILLER_58_1591 ();
 sg13g2_fill_2 FILLER_58_1595 ();
 sg13g2_fill_2 FILLER_58_1610 ();
 sg13g2_decap_8 FILLER_58_1628 ();
 sg13g2_decap_4 FILLER_58_1635 ();
 sg13g2_fill_1 FILLER_58_1639 ();
 sg13g2_decap_8 FILLER_58_1653 ();
 sg13g2_fill_2 FILLER_58_1660 ();
 sg13g2_fill_1 FILLER_58_1662 ();
 sg13g2_fill_1 FILLER_58_1668 ();
 sg13g2_fill_2 FILLER_58_1677 ();
 sg13g2_fill_1 FILLER_58_1679 ();
 sg13g2_fill_2 FILLER_58_1685 ();
 sg13g2_fill_2 FILLER_58_1692 ();
 sg13g2_fill_1 FILLER_58_1694 ();
 sg13g2_decap_8 FILLER_58_1730 ();
 sg13g2_fill_1 FILLER_58_1737 ();
 sg13g2_decap_8 FILLER_58_1756 ();
 sg13g2_decap_4 FILLER_58_1763 ();
 sg13g2_fill_1 FILLER_58_1767 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_4 ();
 sg13g2_fill_1 FILLER_59_33 ();
 sg13g2_fill_2 FILLER_59_53 ();
 sg13g2_fill_1 FILLER_59_55 ();
 sg13g2_fill_2 FILLER_59_61 ();
 sg13g2_fill_2 FILLER_59_91 ();
 sg13g2_fill_2 FILLER_59_123 ();
 sg13g2_fill_2 FILLER_59_129 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_2 FILLER_59_182 ();
 sg13g2_decap_4 FILLER_59_204 ();
 sg13g2_decap_8 FILLER_59_221 ();
 sg13g2_fill_2 FILLER_59_228 ();
 sg13g2_fill_1 FILLER_59_230 ();
 sg13g2_fill_1 FILLER_59_244 ();
 sg13g2_fill_2 FILLER_59_252 ();
 sg13g2_fill_2 FILLER_59_269 ();
 sg13g2_fill_2 FILLER_59_293 ();
 sg13g2_fill_2 FILLER_59_304 ();
 sg13g2_fill_1 FILLER_59_318 ();
 sg13g2_fill_1 FILLER_59_338 ();
 sg13g2_fill_2 FILLER_59_394 ();
 sg13g2_fill_1 FILLER_59_396 ();
 sg13g2_fill_1 FILLER_59_449 ();
 sg13g2_decap_4 FILLER_59_460 ();
 sg13g2_fill_2 FILLER_59_481 ();
 sg13g2_fill_1 FILLER_59_483 ();
 sg13g2_fill_2 FILLER_59_498 ();
 sg13g2_fill_1 FILLER_59_508 ();
 sg13g2_fill_2 FILLER_59_518 ();
 sg13g2_fill_1 FILLER_59_520 ();
 sg13g2_decap_8 FILLER_59_549 ();
 sg13g2_decap_8 FILLER_59_556 ();
 sg13g2_fill_2 FILLER_59_563 ();
 sg13g2_fill_1 FILLER_59_565 ();
 sg13g2_fill_2 FILLER_59_580 ();
 sg13g2_decap_4 FILLER_59_591 ();
 sg13g2_fill_2 FILLER_59_595 ();
 sg13g2_fill_2 FILLER_59_637 ();
 sg13g2_fill_1 FILLER_59_639 ();
 sg13g2_fill_1 FILLER_59_651 ();
 sg13g2_fill_1 FILLER_59_671 ();
 sg13g2_fill_2 FILLER_59_681 ();
 sg13g2_decap_8 FILLER_59_693 ();
 sg13g2_fill_2 FILLER_59_700 ();
 sg13g2_fill_2 FILLER_59_715 ();
 sg13g2_fill_1 FILLER_59_736 ();
 sg13g2_fill_1 FILLER_59_746 ();
 sg13g2_fill_2 FILLER_59_753 ();
 sg13g2_fill_1 FILLER_59_784 ();
 sg13g2_fill_2 FILLER_59_809 ();
 sg13g2_fill_2 FILLER_59_849 ();
 sg13g2_fill_1 FILLER_59_851 ();
 sg13g2_decap_8 FILLER_59_874 ();
 sg13g2_decap_4 FILLER_59_881 ();
 sg13g2_fill_1 FILLER_59_885 ();
 sg13g2_fill_1 FILLER_59_905 ();
 sg13g2_fill_2 FILLER_59_966 ();
 sg13g2_fill_2 FILLER_59_987 ();
 sg13g2_fill_2 FILLER_59_1054 ();
 sg13g2_fill_1 FILLER_59_1071 ();
 sg13g2_fill_2 FILLER_59_1119 ();
 sg13g2_fill_1 FILLER_59_1121 ();
 sg13g2_decap_8 FILLER_59_1150 ();
 sg13g2_fill_2 FILLER_59_1189 ();
 sg13g2_fill_1 FILLER_59_1191 ();
 sg13g2_fill_1 FILLER_59_1201 ();
 sg13g2_fill_2 FILLER_59_1279 ();
 sg13g2_fill_1 FILLER_59_1281 ();
 sg13g2_fill_2 FILLER_59_1295 ();
 sg13g2_decap_8 FILLER_59_1306 ();
 sg13g2_decap_4 FILLER_59_1313 ();
 sg13g2_fill_2 FILLER_59_1317 ();
 sg13g2_decap_4 FILLER_59_1338 ();
 sg13g2_fill_2 FILLER_59_1342 ();
 sg13g2_decap_8 FILLER_59_1354 ();
 sg13g2_fill_1 FILLER_59_1370 ();
 sg13g2_fill_2 FILLER_59_1412 ();
 sg13g2_decap_4 FILLER_59_1419 ();
 sg13g2_fill_1 FILLER_59_1423 ();
 sg13g2_decap_4 FILLER_59_1431 ();
 sg13g2_fill_1 FILLER_59_1435 ();
 sg13g2_fill_2 FILLER_59_1457 ();
 sg13g2_decap_8 FILLER_59_1481 ();
 sg13g2_decap_4 FILLER_59_1488 ();
 sg13g2_fill_1 FILLER_59_1492 ();
 sg13g2_decap_8 FILLER_59_1518 ();
 sg13g2_fill_2 FILLER_59_1529 ();
 sg13g2_fill_1 FILLER_59_1531 ();
 sg13g2_fill_2 FILLER_59_1561 ();
 sg13g2_fill_1 FILLER_59_1563 ();
 sg13g2_fill_2 FILLER_59_1568 ();
 sg13g2_decap_8 FILLER_59_1595 ();
 sg13g2_decap_4 FILLER_59_1602 ();
 sg13g2_decap_8 FILLER_59_1614 ();
 sg13g2_decap_8 FILLER_59_1621 ();
 sg13g2_decap_8 FILLER_59_1628 ();
 sg13g2_decap_4 FILLER_59_1635 ();
 sg13g2_fill_1 FILLER_59_1639 ();
 sg13g2_fill_2 FILLER_59_1643 ();
 sg13g2_decap_8 FILLER_59_1649 ();
 sg13g2_decap_4 FILLER_59_1656 ();
 sg13g2_fill_1 FILLER_59_1660 ();
 sg13g2_decap_8 FILLER_59_1680 ();
 sg13g2_decap_8 FILLER_59_1687 ();
 sg13g2_decap_4 FILLER_59_1694 ();
 sg13g2_fill_2 FILLER_59_1698 ();
 sg13g2_decap_8 FILLER_59_1708 ();
 sg13g2_fill_2 FILLER_59_1728 ();
 sg13g2_fill_1 FILLER_59_1767 ();
 sg13g2_fill_2 FILLER_60_0 ();
 sg13g2_fill_2 FILLER_60_34 ();
 sg13g2_fill_1 FILLER_60_36 ();
 sg13g2_fill_2 FILLER_60_55 ();
 sg13g2_fill_1 FILLER_60_57 ();
 sg13g2_fill_2 FILLER_60_78 ();
 sg13g2_fill_2 FILLER_60_104 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_1 FILLER_60_147 ();
 sg13g2_fill_2 FILLER_60_189 ();
 sg13g2_fill_1 FILLER_60_191 ();
 sg13g2_fill_2 FILLER_60_210 ();
 sg13g2_fill_2 FILLER_60_227 ();
 sg13g2_fill_1 FILLER_60_229 ();
 sg13g2_decap_4 FILLER_60_252 ();
 sg13g2_fill_1 FILLER_60_256 ();
 sg13g2_fill_2 FILLER_60_267 ();
 sg13g2_fill_1 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_288 ();
 sg13g2_decap_4 FILLER_60_351 ();
 sg13g2_fill_2 FILLER_60_355 ();
 sg13g2_fill_1 FILLER_60_363 ();
 sg13g2_decap_4 FILLER_60_381 ();
 sg13g2_fill_1 FILLER_60_434 ();
 sg13g2_decap_4 FILLER_60_462 ();
 sg13g2_fill_1 FILLER_60_494 ();
 sg13g2_fill_2 FILLER_60_523 ();
 sg13g2_decap_4 FILLER_60_538 ();
 sg13g2_fill_2 FILLER_60_542 ();
 sg13g2_fill_1 FILLER_60_576 ();
 sg13g2_decap_8 FILLER_60_587 ();
 sg13g2_decap_4 FILLER_60_594 ();
 sg13g2_fill_1 FILLER_60_601 ();
 sg13g2_decap_4 FILLER_60_606 ();
 sg13g2_fill_2 FILLER_60_614 ();
 sg13g2_fill_2 FILLER_60_646 ();
 sg13g2_fill_1 FILLER_60_648 ();
 sg13g2_decap_8 FILLER_60_676 ();
 sg13g2_fill_1 FILLER_60_683 ();
 sg13g2_fill_1 FILLER_60_716 ();
 sg13g2_fill_1 FILLER_60_796 ();
 sg13g2_fill_1 FILLER_60_825 ();
 sg13g2_fill_2 FILLER_60_830 ();
 sg13g2_fill_2 FILLER_60_841 ();
 sg13g2_fill_1 FILLER_60_843 ();
 sg13g2_fill_1 FILLER_60_858 ();
 sg13g2_fill_2 FILLER_60_893 ();
 sg13g2_decap_8 FILLER_60_899 ();
 sg13g2_decap_4 FILLER_60_906 ();
 sg13g2_fill_1 FILLER_60_910 ();
 sg13g2_fill_1 FILLER_60_915 ();
 sg13g2_fill_2 FILLER_60_947 ();
 sg13g2_fill_1 FILLER_60_954 ();
 sg13g2_fill_1 FILLER_60_964 ();
 sg13g2_fill_1 FILLER_60_1005 ();
 sg13g2_fill_1 FILLER_60_1069 ();
 sg13g2_fill_2 FILLER_60_1101 ();
 sg13g2_fill_1 FILLER_60_1103 ();
 sg13g2_fill_2 FILLER_60_1155 ();
 sg13g2_fill_2 FILLER_60_1277 ();
 sg13g2_decap_4 FILLER_60_1293 ();
 sg13g2_fill_2 FILLER_60_1297 ();
 sg13g2_decap_8 FILLER_60_1319 ();
 sg13g2_fill_1 FILLER_60_1326 ();
 sg13g2_decap_4 FILLER_60_1336 ();
 sg13g2_fill_1 FILLER_60_1340 ();
 sg13g2_decap_4 FILLER_60_1349 ();
 sg13g2_fill_1 FILLER_60_1358 ();
 sg13g2_fill_2 FILLER_60_1371 ();
 sg13g2_fill_1 FILLER_60_1373 ();
 sg13g2_decap_8 FILLER_60_1387 ();
 sg13g2_fill_1 FILLER_60_1394 ();
 sg13g2_decap_4 FILLER_60_1417 ();
 sg13g2_fill_1 FILLER_60_1437 ();
 sg13g2_fill_1 FILLER_60_1466 ();
 sg13g2_decap_8 FILLER_60_1471 ();
 sg13g2_fill_2 FILLER_60_1486 ();
 sg13g2_fill_1 FILLER_60_1488 ();
 sg13g2_decap_8 FILLER_60_1515 ();
 sg13g2_decap_4 FILLER_60_1522 ();
 sg13g2_decap_8 FILLER_60_1534 ();
 sg13g2_fill_1 FILLER_60_1541 ();
 sg13g2_fill_2 FILLER_60_1552 ();
 sg13g2_decap_8 FILLER_60_1558 ();
 sg13g2_decap_8 FILLER_60_1565 ();
 sg13g2_decap_8 FILLER_60_1595 ();
 sg13g2_decap_8 FILLER_60_1602 ();
 sg13g2_decap_4 FILLER_60_1609 ();
 sg13g2_decap_8 FILLER_60_1619 ();
 sg13g2_fill_1 FILLER_60_1626 ();
 sg13g2_decap_8 FILLER_60_1632 ();
 sg13g2_fill_2 FILLER_60_1639 ();
 sg13g2_fill_2 FILLER_60_1650 ();
 sg13g2_fill_2 FILLER_60_1662 ();
 sg13g2_decap_8 FILLER_60_1686 ();
 sg13g2_decap_8 FILLER_60_1693 ();
 sg13g2_decap_8 FILLER_60_1704 ();
 sg13g2_decap_8 FILLER_60_1711 ();
 sg13g2_decap_8 FILLER_60_1731 ();
 sg13g2_fill_2 FILLER_60_1738 ();
 sg13g2_fill_1 FILLER_60_1740 ();
 sg13g2_decap_8 FILLER_60_1757 ();
 sg13g2_decap_4 FILLER_60_1764 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_2 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_103 ();
 sg13g2_fill_1 FILLER_61_105 ();
 sg13g2_decap_8 FILLER_61_124 ();
 sg13g2_decap_4 FILLER_61_131 ();
 sg13g2_fill_2 FILLER_61_162 ();
 sg13g2_fill_1 FILLER_61_164 ();
 sg13g2_fill_1 FILLER_61_178 ();
 sg13g2_decap_4 FILLER_61_225 ();
 sg13g2_decap_8 FILLER_61_247 ();
 sg13g2_decap_8 FILLER_61_290 ();
 sg13g2_fill_1 FILLER_61_305 ();
 sg13g2_fill_1 FILLER_61_309 ();
 sg13g2_decap_8 FILLER_61_337 ();
 sg13g2_decap_8 FILLER_61_392 ();
 sg13g2_fill_2 FILLER_61_399 ();
 sg13g2_fill_1 FILLER_61_401 ();
 sg13g2_fill_1 FILLER_61_409 ();
 sg13g2_fill_1 FILLER_61_419 ();
 sg13g2_fill_1 FILLER_61_429 ();
 sg13g2_fill_1 FILLER_61_444 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_decap_8 FILLER_61_466 ();
 sg13g2_decap_4 FILLER_61_473 ();
 sg13g2_fill_2 FILLER_61_488 ();
 sg13g2_decap_8 FILLER_61_494 ();
 sg13g2_decap_8 FILLER_61_501 ();
 sg13g2_fill_1 FILLER_61_536 ();
 sg13g2_fill_1 FILLER_61_568 ();
 sg13g2_fill_2 FILLER_61_610 ();
 sg13g2_fill_1 FILLER_61_612 ();
 sg13g2_fill_2 FILLER_61_648 ();
 sg13g2_fill_1 FILLER_61_663 ();
 sg13g2_fill_2 FILLER_61_696 ();
 sg13g2_fill_1 FILLER_61_698 ();
 sg13g2_fill_1 FILLER_61_708 ();
 sg13g2_fill_1 FILLER_61_727 ();
 sg13g2_decap_4 FILLER_61_736 ();
 sg13g2_fill_2 FILLER_61_740 ();
 sg13g2_fill_2 FILLER_61_747 ();
 sg13g2_fill_1 FILLER_61_749 ();
 sg13g2_fill_2 FILLER_61_760 ();
 sg13g2_fill_2 FILLER_61_788 ();
 sg13g2_fill_1 FILLER_61_790 ();
 sg13g2_fill_2 FILLER_61_804 ();
 sg13g2_fill_2 FILLER_61_830 ();
 sg13g2_fill_1 FILLER_61_832 ();
 sg13g2_fill_1 FILLER_61_863 ();
 sg13g2_fill_2 FILLER_61_877 ();
 sg13g2_fill_1 FILLER_61_879 ();
 sg13g2_fill_2 FILLER_61_923 ();
 sg13g2_fill_1 FILLER_61_925 ();
 sg13g2_fill_2 FILLER_61_934 ();
 sg13g2_fill_2 FILLER_61_950 ();
 sg13g2_fill_2 FILLER_61_966 ();
 sg13g2_fill_1 FILLER_61_1007 ();
 sg13g2_fill_2 FILLER_61_1026 ();
 sg13g2_fill_1 FILLER_61_1028 ();
 sg13g2_fill_1 FILLER_61_1048 ();
 sg13g2_fill_1 FILLER_61_1058 ();
 sg13g2_fill_1 FILLER_61_1080 ();
 sg13g2_fill_2 FILLER_61_1085 ();
 sg13g2_fill_2 FILLER_61_1145 ();
 sg13g2_fill_2 FILLER_61_1206 ();
 sg13g2_fill_2 FILLER_61_1214 ();
 sg13g2_fill_2 FILLER_61_1225 ();
 sg13g2_fill_2 FILLER_61_1249 ();
 sg13g2_fill_1 FILLER_61_1251 ();
 sg13g2_fill_2 FILLER_61_1282 ();
 sg13g2_fill_1 FILLER_61_1284 ();
 sg13g2_fill_2 FILLER_61_1300 ();
 sg13g2_decap_8 FILLER_61_1310 ();
 sg13g2_decap_4 FILLER_61_1317 ();
 sg13g2_decap_4 FILLER_61_1351 ();
 sg13g2_fill_2 FILLER_61_1368 ();
 sg13g2_fill_1 FILLER_61_1370 ();
 sg13g2_decap_8 FILLER_61_1375 ();
 sg13g2_decap_4 FILLER_61_1382 ();
 sg13g2_fill_1 FILLER_61_1386 ();
 sg13g2_decap_4 FILLER_61_1391 ();
 sg13g2_decap_8 FILLER_61_1408 ();
 sg13g2_decap_4 FILLER_61_1415 ();
 sg13g2_fill_2 FILLER_61_1419 ();
 sg13g2_decap_8 FILLER_61_1434 ();
 sg13g2_decap_4 FILLER_61_1441 ();
 sg13g2_decap_8 FILLER_61_1461 ();
 sg13g2_decap_8 FILLER_61_1468 ();
 sg13g2_fill_1 FILLER_61_1475 ();
 sg13g2_fill_2 FILLER_61_1491 ();
 sg13g2_fill_1 FILLER_61_1493 ();
 sg13g2_fill_2 FILLER_61_1516 ();
 sg13g2_decap_8 FILLER_61_1539 ();
 sg13g2_fill_2 FILLER_61_1546 ();
 sg13g2_fill_1 FILLER_61_1548 ();
 sg13g2_fill_1 FILLER_61_1554 ();
 sg13g2_decap_8 FILLER_61_1560 ();
 sg13g2_decap_8 FILLER_61_1567 ();
 sg13g2_decap_4 FILLER_61_1574 ();
 sg13g2_decap_8 FILLER_61_1594 ();
 sg13g2_fill_2 FILLER_61_1607 ();
 sg13g2_fill_2 FILLER_61_1618 ();
 sg13g2_decap_4 FILLER_61_1641 ();
 sg13g2_fill_2 FILLER_61_1645 ();
 sg13g2_fill_2 FILLER_61_1654 ();
 sg13g2_fill_1 FILLER_61_1656 ();
 sg13g2_decap_8 FILLER_61_1686 ();
 sg13g2_fill_1 FILLER_61_1699 ();
 sg13g2_fill_2 FILLER_61_1715 ();
 sg13g2_decap_8 FILLER_61_1730 ();
 sg13g2_fill_2 FILLER_61_1737 ();
 sg13g2_decap_8 FILLER_61_1756 ();
 sg13g2_decap_4 FILLER_61_1763 ();
 sg13g2_fill_1 FILLER_61_1767 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_2 ();
 sg13g2_fill_2 FILLER_62_35 ();
 sg13g2_fill_1 FILLER_62_37 ();
 sg13g2_fill_2 FILLER_62_64 ();
 sg13g2_fill_1 FILLER_62_73 ();
 sg13g2_decap_8 FILLER_62_131 ();
 sg13g2_fill_1 FILLER_62_138 ();
 sg13g2_fill_2 FILLER_62_157 ();
 sg13g2_fill_1 FILLER_62_159 ();
 sg13g2_decap_8 FILLER_62_174 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_decap_8 FILLER_62_240 ();
 sg13g2_fill_2 FILLER_62_257 ();
 sg13g2_fill_1 FILLER_62_263 ();
 sg13g2_decap_4 FILLER_62_273 ();
 sg13g2_fill_1 FILLER_62_277 ();
 sg13g2_fill_2 FILLER_62_290 ();
 sg13g2_decap_8 FILLER_62_319 ();
 sg13g2_decap_4 FILLER_62_326 ();
 sg13g2_fill_2 FILLER_62_334 ();
 sg13g2_fill_1 FILLER_62_336 ();
 sg13g2_fill_2 FILLER_62_350 ();
 sg13g2_fill_1 FILLER_62_352 ();
 sg13g2_decap_4 FILLER_62_357 ();
 sg13g2_decap_4 FILLER_62_375 ();
 sg13g2_fill_1 FILLER_62_379 ();
 sg13g2_decap_8 FILLER_62_383 ();
 sg13g2_decap_4 FILLER_62_390 ();
 sg13g2_fill_1 FILLER_62_394 ();
 sg13g2_decap_8 FILLER_62_465 ();
 sg13g2_fill_2 FILLER_62_472 ();
 sg13g2_fill_1 FILLER_62_474 ();
 sg13g2_decap_8 FILLER_62_492 ();
 sg13g2_fill_2 FILLER_62_499 ();
 sg13g2_fill_1 FILLER_62_501 ();
 sg13g2_decap_4 FILLER_62_508 ();
 sg13g2_fill_1 FILLER_62_512 ();
 sg13g2_fill_1 FILLER_62_517 ();
 sg13g2_decap_8 FILLER_62_581 ();
 sg13g2_fill_2 FILLER_62_606 ();
 sg13g2_fill_1 FILLER_62_664 ();
 sg13g2_fill_2 FILLER_62_678 ();
 sg13g2_fill_1 FILLER_62_680 ();
 sg13g2_decap_8 FILLER_62_685 ();
 sg13g2_decap_8 FILLER_62_692 ();
 sg13g2_fill_1 FILLER_62_699 ();
 sg13g2_fill_2 FILLER_62_724 ();
 sg13g2_decap_8 FILLER_62_730 ();
 sg13g2_decap_4 FILLER_62_737 ();
 sg13g2_fill_1 FILLER_62_741 ();
 sg13g2_fill_2 FILLER_62_748 ();
 sg13g2_fill_1 FILLER_62_750 ();
 sg13g2_fill_2 FILLER_62_771 ();
 sg13g2_fill_2 FILLER_62_777 ();
 sg13g2_fill_1 FILLER_62_779 ();
 sg13g2_fill_2 FILLER_62_793 ();
 sg13g2_decap_8 FILLER_62_895 ();
 sg13g2_decap_4 FILLER_62_902 ();
 sg13g2_decap_4 FILLER_62_920 ();
 sg13g2_fill_1 FILLER_62_924 ();
 sg13g2_fill_1 FILLER_62_952 ();
 sg13g2_fill_1 FILLER_62_985 ();
 sg13g2_fill_1 FILLER_62_1022 ();
 sg13g2_fill_1 FILLER_62_1059 ();
 sg13g2_fill_1 FILLER_62_1083 ();
 sg13g2_decap_8 FILLER_62_1144 ();
 sg13g2_fill_2 FILLER_62_1151 ();
 sg13g2_decap_4 FILLER_62_1188 ();
 sg13g2_decap_4 FILLER_62_1318 ();
 sg13g2_fill_2 FILLER_62_1322 ();
 sg13g2_decap_8 FILLER_62_1329 ();
 sg13g2_fill_2 FILLER_62_1336 ();
 sg13g2_fill_1 FILLER_62_1338 ();
 sg13g2_decap_8 FILLER_62_1343 ();
 sg13g2_decap_4 FILLER_62_1378 ();
 sg13g2_decap_4 FILLER_62_1410 ();
 sg13g2_decap_8 FILLER_62_1446 ();
 sg13g2_decap_8 FILLER_62_1453 ();
 sg13g2_decap_8 FILLER_62_1460 ();
 sg13g2_fill_2 FILLER_62_1467 ();
 sg13g2_decap_8 FILLER_62_1473 ();
 sg13g2_decap_4 FILLER_62_1480 ();
 sg13g2_decap_4 FILLER_62_1487 ();
 sg13g2_decap_8 FILLER_62_1498 ();
 sg13g2_decap_8 FILLER_62_1505 ();
 sg13g2_decap_4 FILLER_62_1512 ();
 sg13g2_fill_1 FILLER_62_1516 ();
 sg13g2_decap_8 FILLER_62_1537 ();
 sg13g2_fill_2 FILLER_62_1544 ();
 sg13g2_decap_8 FILLER_62_1565 ();
 sg13g2_fill_1 FILLER_62_1572 ();
 sg13g2_decap_8 FILLER_62_1589 ();
 sg13g2_decap_4 FILLER_62_1596 ();
 sg13g2_fill_2 FILLER_62_1609 ();
 sg13g2_decap_8 FILLER_62_1643 ();
 sg13g2_fill_2 FILLER_62_1664 ();
 sg13g2_fill_1 FILLER_62_1666 ();
 sg13g2_decap_8 FILLER_62_1672 ();
 sg13g2_fill_2 FILLER_62_1679 ();
 sg13g2_fill_1 FILLER_62_1681 ();
 sg13g2_decap_8 FILLER_62_1717 ();
 sg13g2_fill_2 FILLER_62_1724 ();
 sg13g2_fill_1 FILLER_62_1726 ();
 sg13g2_decap_8 FILLER_62_1759 ();
 sg13g2_fill_2 FILLER_62_1766 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_40 ();
 sg13g2_fill_1 FILLER_63_42 ();
 sg13g2_fill_1 FILLER_63_70 ();
 sg13g2_fill_2 FILLER_63_100 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_fill_2 FILLER_63_203 ();
 sg13g2_fill_1 FILLER_63_205 ();
 sg13g2_fill_2 FILLER_63_215 ();
 sg13g2_fill_2 FILLER_63_234 ();
 sg13g2_fill_1 FILLER_63_249 ();
 sg13g2_decap_8 FILLER_63_278 ();
 sg13g2_fill_2 FILLER_63_285 ();
 sg13g2_fill_1 FILLER_63_287 ();
 sg13g2_fill_1 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_403 ();
 sg13g2_decap_4 FILLER_63_435 ();
 sg13g2_fill_1 FILLER_63_443 ();
 sg13g2_fill_2 FILLER_63_475 ();
 sg13g2_fill_1 FILLER_63_477 ();
 sg13g2_fill_1 FILLER_63_494 ();
 sg13g2_fill_1 FILLER_63_504 ();
 sg13g2_fill_1 FILLER_63_532 ();
 sg13g2_fill_2 FILLER_63_537 ();
 sg13g2_fill_1 FILLER_63_539 ();
 sg13g2_decap_4 FILLER_63_553 ();
 sg13g2_fill_1 FILLER_63_557 ();
 sg13g2_decap_4 FILLER_63_562 ();
 sg13g2_fill_2 FILLER_63_566 ();
 sg13g2_fill_2 FILLER_63_576 ();
 sg13g2_fill_1 FILLER_63_578 ();
 sg13g2_fill_2 FILLER_63_622 ();
 sg13g2_decap_8 FILLER_63_666 ();
 sg13g2_fill_1 FILLER_63_673 ();
 sg13g2_fill_2 FILLER_63_706 ();
 sg13g2_fill_1 FILLER_63_708 ();
 sg13g2_fill_2 FILLER_63_718 ();
 sg13g2_fill_1 FILLER_63_720 ();
 sg13g2_fill_2 FILLER_63_758 ();
 sg13g2_fill_2 FILLER_63_766 ();
 sg13g2_fill_1 FILLER_63_802 ();
 sg13g2_fill_2 FILLER_63_942 ();
 sg13g2_fill_1 FILLER_63_944 ();
 sg13g2_fill_1 FILLER_63_955 ();
 sg13g2_fill_2 FILLER_63_961 ();
 sg13g2_fill_1 FILLER_63_963 ();
 sg13g2_fill_1 FILLER_63_992 ();
 sg13g2_fill_2 FILLER_63_1030 ();
 sg13g2_fill_1 FILLER_63_1048 ();
 sg13g2_decap_8 FILLER_63_1059 ();
 sg13g2_decap_4 FILLER_63_1066 ();
 sg13g2_fill_1 FILLER_63_1070 ();
 sg13g2_fill_2 FILLER_63_1088 ();
 sg13g2_fill_1 FILLER_63_1090 ();
 sg13g2_decap_4 FILLER_63_1131 ();
 sg13g2_fill_1 FILLER_63_1135 ();
 sg13g2_decap_4 FILLER_63_1153 ();
 sg13g2_decap_8 FILLER_63_1189 ();
 sg13g2_fill_1 FILLER_63_1228 ();
 sg13g2_fill_1 FILLER_63_1274 ();
 sg13g2_fill_2 FILLER_63_1288 ();
 sg13g2_fill_1 FILLER_63_1290 ();
 sg13g2_fill_1 FILLER_63_1310 ();
 sg13g2_decap_8 FILLER_63_1321 ();
 sg13g2_decap_4 FILLER_63_1328 ();
 sg13g2_fill_2 FILLER_63_1332 ();
 sg13g2_decap_8 FILLER_63_1349 ();
 sg13g2_decap_4 FILLER_63_1356 ();
 sg13g2_fill_1 FILLER_63_1360 ();
 sg13g2_decap_8 FILLER_63_1371 ();
 sg13g2_decap_8 FILLER_63_1382 ();
 sg13g2_fill_2 FILLER_63_1404 ();
 sg13g2_fill_1 FILLER_63_1406 ();
 sg13g2_fill_2 FILLER_63_1425 ();
 sg13g2_fill_1 FILLER_63_1500 ();
 sg13g2_decap_8 FILLER_63_1506 ();
 sg13g2_decap_8 FILLER_63_1513 ();
 sg13g2_fill_1 FILLER_63_1520 ();
 sg13g2_decap_4 FILLER_63_1537 ();
 sg13g2_fill_2 FILLER_63_1541 ();
 sg13g2_fill_1 FILLER_63_1569 ();
 sg13g2_decap_8 FILLER_63_1582 ();
 sg13g2_decap_8 FILLER_63_1589 ();
 sg13g2_decap_8 FILLER_63_1614 ();
 sg13g2_fill_1 FILLER_63_1621 ();
 sg13g2_fill_1 FILLER_63_1633 ();
 sg13g2_fill_2 FILLER_63_1639 ();
 sg13g2_decap_4 FILLER_63_1651 ();
 sg13g2_decap_8 FILLER_63_1670 ();
 sg13g2_decap_4 FILLER_63_1677 ();
 sg13g2_fill_1 FILLER_63_1681 ();
 sg13g2_fill_2 FILLER_63_1698 ();
 sg13g2_fill_1 FILLER_63_1700 ();
 sg13g2_decap_8 FILLER_63_1710 ();
 sg13g2_decap_8 FILLER_63_1729 ();
 sg13g2_fill_2 FILLER_63_1736 ();
 sg13g2_fill_1 FILLER_63_1738 ();
 sg13g2_decap_8 FILLER_63_1758 ();
 sg13g2_fill_2 FILLER_63_1765 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_decap_4 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_4 ();
 sg13g2_fill_1 FILLER_64_32 ();
 sg13g2_fill_2 FILLER_64_47 ();
 sg13g2_fill_2 FILLER_64_63 ();
 sg13g2_fill_2 FILLER_64_74 ();
 sg13g2_decap_4 FILLER_64_119 ();
 sg13g2_fill_1 FILLER_64_123 ();
 sg13g2_decap_8 FILLER_64_128 ();
 sg13g2_decap_8 FILLER_64_135 ();
 sg13g2_decap_8 FILLER_64_142 ();
 sg13g2_fill_2 FILLER_64_157 ();
 sg13g2_decap_4 FILLER_64_162 ();
 sg13g2_fill_1 FILLER_64_166 ();
 sg13g2_decap_4 FILLER_64_184 ();
 sg13g2_fill_1 FILLER_64_208 ();
 sg13g2_fill_1 FILLER_64_254 ();
 sg13g2_decap_8 FILLER_64_259 ();
 sg13g2_decap_8 FILLER_64_283 ();
 sg13g2_fill_2 FILLER_64_290 ();
 sg13g2_fill_1 FILLER_64_292 ();
 sg13g2_fill_2 FILLER_64_297 ();
 sg13g2_fill_1 FILLER_64_299 ();
 sg13g2_fill_2 FILLER_64_313 ();
 sg13g2_fill_1 FILLER_64_315 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_decap_8 FILLER_64_336 ();
 sg13g2_decap_8 FILLER_64_343 ();
 sg13g2_fill_2 FILLER_64_350 ();
 sg13g2_decap_8 FILLER_64_364 ();
 sg13g2_decap_4 FILLER_64_371 ();
 sg13g2_decap_8 FILLER_64_394 ();
 sg13g2_fill_2 FILLER_64_401 ();
 sg13g2_fill_2 FILLER_64_441 ();
 sg13g2_fill_2 FILLER_64_467 ();
 sg13g2_fill_1 FILLER_64_469 ();
 sg13g2_fill_2 FILLER_64_479 ();
 sg13g2_fill_1 FILLER_64_481 ();
 sg13g2_fill_2 FILLER_64_509 ();
 sg13g2_fill_1 FILLER_64_511 ();
 sg13g2_fill_2 FILLER_64_571 ();
 sg13g2_fill_1 FILLER_64_573 ();
 sg13g2_fill_2 FILLER_64_604 ();
 sg13g2_fill_1 FILLER_64_606 ();
 sg13g2_fill_2 FILLER_64_655 ();
 sg13g2_decap_8 FILLER_64_670 ();
 sg13g2_decap_4 FILLER_64_677 ();
 sg13g2_fill_2 FILLER_64_681 ();
 sg13g2_decap_8 FILLER_64_687 ();
 sg13g2_decap_4 FILLER_64_694 ();
 sg13g2_fill_1 FILLER_64_698 ();
 sg13g2_fill_1 FILLER_64_721 ();
 sg13g2_fill_2 FILLER_64_735 ();
 sg13g2_decap_4 FILLER_64_772 ();
 sg13g2_fill_2 FILLER_64_793 ();
 sg13g2_fill_2 FILLER_64_855 ();
 sg13g2_fill_1 FILLER_64_857 ();
 sg13g2_decap_4 FILLER_64_886 ();
 sg13g2_decap_8 FILLER_64_894 ();
 sg13g2_fill_2 FILLER_64_901 ();
 sg13g2_fill_1 FILLER_64_903 ();
 sg13g2_fill_2 FILLER_64_917 ();
 sg13g2_fill_1 FILLER_64_932 ();
 sg13g2_fill_2 FILLER_64_1058 ();
 sg13g2_decap_8 FILLER_64_1104 ();
 sg13g2_fill_2 FILLER_64_1111 ();
 sg13g2_decap_8 FILLER_64_1136 ();
 sg13g2_fill_2 FILLER_64_1143 ();
 sg13g2_fill_2 FILLER_64_1155 ();
 sg13g2_fill_1 FILLER_64_1157 ();
 sg13g2_decap_8 FILLER_64_1185 ();
 sg13g2_fill_2 FILLER_64_1192 ();
 sg13g2_fill_2 FILLER_64_1207 ();
 sg13g2_fill_2 FILLER_64_1284 ();
 sg13g2_fill_1 FILLER_64_1286 ();
 sg13g2_decap_4 FILLER_64_1291 ();
 sg13g2_fill_2 FILLER_64_1295 ();
 sg13g2_fill_2 FILLER_64_1302 ();
 sg13g2_fill_1 FILLER_64_1304 ();
 sg13g2_decap_8 FILLER_64_1315 ();
 sg13g2_fill_2 FILLER_64_1322 ();
 sg13g2_decap_4 FILLER_64_1367 ();
 sg13g2_fill_2 FILLER_64_1371 ();
 sg13g2_fill_1 FILLER_64_1400 ();
 sg13g2_fill_2 FILLER_64_1429 ();
 sg13g2_decap_8 FILLER_64_1463 ();
 sg13g2_decap_8 FILLER_64_1470 ();
 sg13g2_decap_8 FILLER_64_1517 ();
 sg13g2_fill_2 FILLER_64_1524 ();
 sg13g2_decap_4 FILLER_64_1530 ();
 sg13g2_fill_1 FILLER_64_1534 ();
 sg13g2_decap_8 FILLER_64_1541 ();
 sg13g2_fill_1 FILLER_64_1548 ();
 sg13g2_fill_1 FILLER_64_1573 ();
 sg13g2_decap_8 FILLER_64_1584 ();
 sg13g2_decap_4 FILLER_64_1591 ();
 sg13g2_fill_1 FILLER_64_1595 ();
 sg13g2_decap_8 FILLER_64_1611 ();
 sg13g2_decap_4 FILLER_64_1626 ();
 sg13g2_decap_8 FILLER_64_1635 ();
 sg13g2_fill_1 FILLER_64_1642 ();
 sg13g2_fill_1 FILLER_64_1656 ();
 sg13g2_fill_1 FILLER_64_1674 ();
 sg13g2_fill_1 FILLER_64_1684 ();
 sg13g2_decap_4 FILLER_64_1710 ();
 sg13g2_fill_1 FILLER_64_1714 ();
 sg13g2_fill_2 FILLER_64_1724 ();
 sg13g2_decap_4 FILLER_64_1731 ();
 sg13g2_fill_2 FILLER_64_1735 ();
 sg13g2_fill_2 FILLER_64_1766 ();
 sg13g2_decap_4 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_4 ();
 sg13g2_fill_1 FILLER_65_43 ();
 sg13g2_decap_4 FILLER_65_113 ();
 sg13g2_fill_1 FILLER_65_117 ();
 sg13g2_decap_4 FILLER_65_172 ();
 sg13g2_fill_1 FILLER_65_176 ();
 sg13g2_fill_1 FILLER_65_187 ();
 sg13g2_decap_8 FILLER_65_198 ();
 sg13g2_fill_2 FILLER_65_205 ();
 sg13g2_fill_1 FILLER_65_207 ();
 sg13g2_fill_1 FILLER_65_216 ();
 sg13g2_decap_8 FILLER_65_222 ();
 sg13g2_decap_8 FILLER_65_229 ();
 sg13g2_decap_4 FILLER_65_241 ();
 sg13g2_decap_4 FILLER_65_253 ();
 sg13g2_fill_1 FILLER_65_257 ();
 sg13g2_decap_4 FILLER_65_299 ();
 sg13g2_fill_1 FILLER_65_303 ();
 sg13g2_fill_1 FILLER_65_317 ();
 sg13g2_fill_2 FILLER_65_354 ();
 sg13g2_fill_1 FILLER_65_384 ();
 sg13g2_decap_8 FILLER_65_389 ();
 sg13g2_fill_1 FILLER_65_396 ();
 sg13g2_fill_1 FILLER_65_410 ();
 sg13g2_decap_8 FILLER_65_417 ();
 sg13g2_fill_2 FILLER_65_435 ();
 sg13g2_fill_1 FILLER_65_437 ();
 sg13g2_fill_2 FILLER_65_441 ();
 sg13g2_fill_2 FILLER_65_481 ();
 sg13g2_decap_4 FILLER_65_501 ();
 sg13g2_fill_1 FILLER_65_584 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_4 FILLER_65_658 ();
 sg13g2_fill_2 FILLER_65_731 ();
 sg13g2_fill_2 FILLER_65_773 ();
 sg13g2_fill_2 FILLER_65_807 ();
 sg13g2_fill_1 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_841 ();
 sg13g2_decap_4 FILLER_65_858 ();
 sg13g2_fill_1 FILLER_65_862 ();
 sg13g2_fill_1 FILLER_65_876 ();
 sg13g2_fill_1 FILLER_65_894 ();
 sg13g2_decap_4 FILLER_65_931 ();
 sg13g2_fill_1 FILLER_65_943 ();
 sg13g2_fill_1 FILLER_65_949 ();
 sg13g2_fill_2 FILLER_65_955 ();
 sg13g2_decap_4 FILLER_65_970 ();
 sg13g2_fill_2 FILLER_65_978 ();
 sg13g2_fill_1 FILLER_65_980 ();
 sg13g2_fill_2 FILLER_65_1012 ();
 sg13g2_fill_1 FILLER_65_1014 ();
 sg13g2_fill_2 FILLER_65_1038 ();
 sg13g2_decap_8 FILLER_65_1050 ();
 sg13g2_decap_4 FILLER_65_1057 ();
 sg13g2_fill_1 FILLER_65_1061 ();
 sg13g2_fill_1 FILLER_65_1080 ();
 sg13g2_decap_4 FILLER_65_1090 ();
 sg13g2_decap_4 FILLER_65_1114 ();
 sg13g2_decap_4 FILLER_65_1132 ();
 sg13g2_fill_1 FILLER_65_1136 ();
 sg13g2_decap_8 FILLER_65_1157 ();
 sg13g2_decap_8 FILLER_65_1164 ();
 sg13g2_decap_4 FILLER_65_1184 ();
 sg13g2_fill_1 FILLER_65_1188 ();
 sg13g2_decap_8 FILLER_65_1199 ();
 sg13g2_decap_8 FILLER_65_1219 ();
 sg13g2_fill_2 FILLER_65_1226 ();
 sg13g2_fill_2 FILLER_65_1245 ();
 sg13g2_fill_1 FILLER_65_1247 ();
 sg13g2_decap_4 FILLER_65_1275 ();
 sg13g2_fill_2 FILLER_65_1279 ();
 sg13g2_decap_8 FILLER_65_1291 ();
 sg13g2_fill_2 FILLER_65_1298 ();
 sg13g2_decap_4 FILLER_65_1350 ();
 sg13g2_fill_2 FILLER_65_1354 ();
 sg13g2_decap_8 FILLER_65_1376 ();
 sg13g2_fill_2 FILLER_65_1383 ();
 sg13g2_fill_1 FILLER_65_1385 ();
 sg13g2_fill_2 FILLER_65_1395 ();
 sg13g2_fill_2 FILLER_65_1415 ();
 sg13g2_fill_2 FILLER_65_1478 ();
 sg13g2_fill_1 FILLER_65_1480 ();
 sg13g2_fill_1 FILLER_65_1535 ();
 sg13g2_fill_2 FILLER_65_1549 ();
 sg13g2_fill_1 FILLER_65_1567 ();
 sg13g2_decap_8 FILLER_65_1573 ();
 sg13g2_decap_4 FILLER_65_1588 ();
 sg13g2_fill_2 FILLER_65_1592 ();
 sg13g2_decap_8 FILLER_65_1602 ();
 sg13g2_fill_2 FILLER_65_1609 ();
 sg13g2_fill_2 FILLER_65_1627 ();
 sg13g2_fill_1 FILLER_65_1629 ();
 sg13g2_fill_1 FILLER_65_1635 ();
 sg13g2_decap_8 FILLER_65_1643 ();
 sg13g2_decap_8 FILLER_65_1650 ();
 sg13g2_decap_8 FILLER_65_1657 ();
 sg13g2_decap_4 FILLER_65_1664 ();
 sg13g2_decap_8 FILLER_65_1687 ();
 sg13g2_fill_1 FILLER_65_1694 ();
 sg13g2_decap_8 FILLER_65_1700 ();
 sg13g2_fill_2 FILLER_65_1707 ();
 sg13g2_fill_1 FILLER_65_1709 ();
 sg13g2_fill_2 FILLER_65_1716 ();
 sg13g2_fill_2 FILLER_65_1743 ();
 sg13g2_fill_1 FILLER_65_1745 ();
 sg13g2_fill_2 FILLER_65_1766 ();
 sg13g2_fill_2 FILLER_66_44 ();
 sg13g2_fill_2 FILLER_66_100 ();
 sg13g2_decap_4 FILLER_66_106 ();
 sg13g2_fill_1 FILLER_66_110 ();
 sg13g2_fill_1 FILLER_66_154 ();
 sg13g2_decap_8 FILLER_66_175 ();
 sg13g2_fill_2 FILLER_66_182 ();
 sg13g2_fill_2 FILLER_66_238 ();
 sg13g2_fill_1 FILLER_66_240 ();
 sg13g2_fill_2 FILLER_66_257 ();
 sg13g2_decap_4 FILLER_66_263 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_1 FILLER_66_281 ();
 sg13g2_fill_2 FILLER_66_292 ();
 sg13g2_fill_1 FILLER_66_294 ();
 sg13g2_fill_2 FILLER_66_304 ();
 sg13g2_fill_2 FILLER_66_327 ();
 sg13g2_fill_1 FILLER_66_329 ();
 sg13g2_fill_2 FILLER_66_347 ();
 sg13g2_decap_4 FILLER_66_368 ();
 sg13g2_fill_1 FILLER_66_372 ();
 sg13g2_decap_4 FILLER_66_427 ();
 sg13g2_fill_1 FILLER_66_431 ();
 sg13g2_fill_2 FILLER_66_465 ();
 sg13g2_fill_1 FILLER_66_467 ();
 sg13g2_fill_1 FILLER_66_501 ();
 sg13g2_fill_2 FILLER_66_530 ();
 sg13g2_fill_1 FILLER_66_532 ();
 sg13g2_fill_2 FILLER_66_568 ();
 sg13g2_fill_1 FILLER_66_578 ();
 sg13g2_fill_2 FILLER_66_588 ();
 sg13g2_fill_1 FILLER_66_638 ();
 sg13g2_decap_4 FILLER_66_647 ();
 sg13g2_decap_4 FILLER_66_661 ();
 sg13g2_fill_2 FILLER_66_665 ();
 sg13g2_fill_1 FILLER_66_685 ();
 sg13g2_decap_8 FILLER_66_712 ();
 sg13g2_fill_1 FILLER_66_719 ();
 sg13g2_fill_2 FILLER_66_729 ();
 sg13g2_fill_1 FILLER_66_737 ();
 sg13g2_decap_8 FILLER_66_742 ();
 sg13g2_decap_4 FILLER_66_749 ();
 sg13g2_fill_1 FILLER_66_753 ();
 sg13g2_fill_2 FILLER_66_781 ();
 sg13g2_decap_4 FILLER_66_792 ();
 sg13g2_fill_1 FILLER_66_796 ();
 sg13g2_decap_8 FILLER_66_829 ();
 sg13g2_decap_4 FILLER_66_836 ();
 sg13g2_fill_2 FILLER_66_840 ();
 sg13g2_decap_8 FILLER_66_868 ();
 sg13g2_fill_2 FILLER_66_875 ();
 sg13g2_fill_2 FILLER_66_931 ();
 sg13g2_fill_2 FILLER_66_975 ();
 sg13g2_fill_1 FILLER_66_977 ();
 sg13g2_fill_2 FILLER_66_983 ();
 sg13g2_decap_4 FILLER_66_990 ();
 sg13g2_fill_1 FILLER_66_994 ();
 sg13g2_fill_2 FILLER_66_1018 ();
 sg13g2_decap_8 FILLER_66_1047 ();
 sg13g2_decap_4 FILLER_66_1054 ();
 sg13g2_fill_2 FILLER_66_1080 ();
 sg13g2_fill_1 FILLER_66_1082 ();
 sg13g2_decap_4 FILLER_66_1093 ();
 sg13g2_fill_1 FILLER_66_1097 ();
 sg13g2_fill_2 FILLER_66_1112 ();
 sg13g2_fill_1 FILLER_66_1114 ();
 sg13g2_fill_2 FILLER_66_1135 ();
 sg13g2_decap_8 FILLER_66_1147 ();
 sg13g2_decap_8 FILLER_66_1154 ();
 sg13g2_decap_4 FILLER_66_1161 ();
 sg13g2_fill_1 FILLER_66_1165 ();
 sg13g2_decap_4 FILLER_66_1186 ();
 sg13g2_fill_1 FILLER_66_1190 ();
 sg13g2_fill_2 FILLER_66_1211 ();
 sg13g2_fill_1 FILLER_66_1213 ();
 sg13g2_decap_8 FILLER_66_1224 ();
 sg13g2_fill_2 FILLER_66_1231 ();
 sg13g2_decap_4 FILLER_66_1277 ();
 sg13g2_fill_1 FILLER_66_1281 ();
 sg13g2_fill_2 FILLER_66_1302 ();
 sg13g2_fill_1 FILLER_66_1304 ();
 sg13g2_decap_4 FILLER_66_1315 ();
 sg13g2_fill_1 FILLER_66_1319 ();
 sg13g2_decap_8 FILLER_66_1330 ();
 sg13g2_fill_1 FILLER_66_1337 ();
 sg13g2_fill_2 FILLER_66_1348 ();
 sg13g2_decap_8 FILLER_66_1378 ();
 sg13g2_decap_4 FILLER_66_1385 ();
 sg13g2_fill_1 FILLER_66_1397 ();
 sg13g2_decap_4 FILLER_66_1416 ();
 sg13g2_fill_1 FILLER_66_1448 ();
 sg13g2_decap_4 FILLER_66_1472 ();
 sg13g2_fill_2 FILLER_66_1504 ();
 sg13g2_fill_2 FILLER_66_1534 ();
 sg13g2_fill_2 FILLER_66_1554 ();
 sg13g2_decap_8 FILLER_66_1574 ();
 sg13g2_fill_2 FILLER_66_1581 ();
 sg13g2_fill_1 FILLER_66_1583 ();
 sg13g2_fill_2 FILLER_66_1589 ();
 sg13g2_fill_1 FILLER_66_1591 ();
 sg13g2_decap_4 FILLER_66_1604 ();
 sg13g2_fill_1 FILLER_66_1608 ();
 sg13g2_fill_2 FILLER_66_1656 ();
 sg13g2_fill_2 FILLER_66_1688 ();
 sg13g2_fill_1 FILLER_66_1707 ();
 sg13g2_decap_4 FILLER_66_1712 ();
 sg13g2_fill_1 FILLER_66_1716 ();
 sg13g2_decap_4 FILLER_66_1727 ();
 sg13g2_decap_8 FILLER_66_1736 ();
 sg13g2_decap_8 FILLER_66_1754 ();
 sg13g2_decap_8 FILLER_66_1761 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_fill_2 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_61 ();
 sg13g2_fill_2 FILLER_67_95 ();
 sg13g2_fill_2 FILLER_67_172 ();
 sg13g2_fill_1 FILLER_67_174 ();
 sg13g2_decap_8 FILLER_67_193 ();
 sg13g2_fill_2 FILLER_67_200 ();
 sg13g2_fill_1 FILLER_67_202 ();
 sg13g2_fill_1 FILLER_67_264 ();
 sg13g2_decap_8 FILLER_67_379 ();
 sg13g2_decap_8 FILLER_67_386 ();
 sg13g2_fill_2 FILLER_67_393 ();
 sg13g2_fill_1 FILLER_67_395 ();
 sg13g2_fill_1 FILLER_67_422 ();
 sg13g2_decap_4 FILLER_67_460 ();
 sg13g2_fill_2 FILLER_67_464 ();
 sg13g2_decap_8 FILLER_67_505 ();
 sg13g2_decap_4 FILLER_67_512 ();
 sg13g2_fill_1 FILLER_67_562 ();
 sg13g2_fill_1 FILLER_67_590 ();
 sg13g2_fill_2 FILLER_67_595 ();
 sg13g2_fill_1 FILLER_67_597 ();
 sg13g2_fill_1 FILLER_67_625 ();
 sg13g2_fill_2 FILLER_67_630 ();
 sg13g2_fill_1 FILLER_67_632 ();
 sg13g2_fill_2 FILLER_67_665 ();
 sg13g2_fill_1 FILLER_67_667 ();
 sg13g2_decap_8 FILLER_67_704 ();
 sg13g2_fill_1 FILLER_67_711 ();
 sg13g2_decap_8 FILLER_67_716 ();
 sg13g2_decap_4 FILLER_67_723 ();
 sg13g2_fill_1 FILLER_67_727 ();
 sg13g2_fill_1 FILLER_67_754 ();
 sg13g2_fill_1 FILLER_67_759 ();
 sg13g2_fill_1 FILLER_67_801 ();
 sg13g2_decap_4 FILLER_67_824 ();
 sg13g2_fill_2 FILLER_67_828 ();
 sg13g2_fill_2 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_863 ();
 sg13g2_decap_8 FILLER_67_883 ();
 sg13g2_decap_4 FILLER_67_890 ();
 sg13g2_fill_2 FILLER_67_894 ();
 sg13g2_fill_1 FILLER_67_913 ();
 sg13g2_fill_2 FILLER_67_928 ();
 sg13g2_fill_1 FILLER_67_930 ();
 sg13g2_decap_8 FILLER_67_944 ();
 sg13g2_decap_8 FILLER_67_951 ();
 sg13g2_fill_2 FILLER_67_958 ();
 sg13g2_fill_1 FILLER_67_992 ();
 sg13g2_fill_2 FILLER_67_1011 ();
 sg13g2_decap_4 FILLER_67_1038 ();
 sg13g2_fill_2 FILLER_67_1042 ();
 sg13g2_fill_2 FILLER_67_1050 ();
 sg13g2_fill_1 FILLER_67_1052 ();
 sg13g2_fill_1 FILLER_67_1058 ();
 sg13g2_fill_1 FILLER_67_1094 ();
 sg13g2_fill_2 FILLER_67_1123 ();
 sg13g2_fill_1 FILLER_67_1125 ();
 sg13g2_fill_2 FILLER_67_1135 ();
 sg13g2_fill_2 FILLER_67_1165 ();
 sg13g2_decap_4 FILLER_67_1177 ();
 sg13g2_fill_1 FILLER_67_1207 ();
 sg13g2_fill_1 FILLER_67_1218 ();
 sg13g2_fill_1 FILLER_67_1253 ();
 sg13g2_fill_2 FILLER_67_1263 ();
 sg13g2_decap_8 FILLER_67_1275 ();
 sg13g2_decap_4 FILLER_67_1282 ();
 sg13g2_fill_1 FILLER_67_1296 ();
 sg13g2_decap_8 FILLER_67_1325 ();
 sg13g2_decap_4 FILLER_67_1332 ();
 sg13g2_fill_2 FILLER_67_1336 ();
 sg13g2_fill_2 FILLER_67_1417 ();
 sg13g2_fill_1 FILLER_67_1419 ();
 sg13g2_fill_1 FILLER_67_1461 ();
 sg13g2_fill_2 FILLER_67_1478 ();
 sg13g2_fill_1 FILLER_67_1480 ();
 sg13g2_fill_1 FILLER_67_1485 ();
 sg13g2_decap_4 FILLER_67_1504 ();
 sg13g2_fill_2 FILLER_67_1543 ();
 sg13g2_decap_4 FILLER_67_1573 ();
 sg13g2_fill_2 FILLER_67_1577 ();
 sg13g2_decap_8 FILLER_67_1603 ();
 sg13g2_fill_2 FILLER_67_1610 ();
 sg13g2_fill_1 FILLER_67_1612 ();
 sg13g2_decap_8 FILLER_67_1626 ();
 sg13g2_decap_8 FILLER_67_1633 ();
 sg13g2_fill_2 FILLER_67_1640 ();
 sg13g2_fill_1 FILLER_67_1642 ();
 sg13g2_fill_2 FILLER_67_1689 ();
 sg13g2_fill_1 FILLER_67_1691 ();
 sg13g2_decap_4 FILLER_67_1705 ();
 sg13g2_fill_1 FILLER_67_1709 ();
 sg13g2_fill_2 FILLER_67_1719 ();
 sg13g2_fill_2 FILLER_67_1734 ();
 sg13g2_fill_1 FILLER_67_1736 ();
 sg13g2_decap_8 FILLER_67_1750 ();
 sg13g2_decap_8 FILLER_67_1757 ();
 sg13g2_decap_4 FILLER_67_1764 ();
 sg13g2_fill_2 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_54 ();
 sg13g2_fill_2 FILLER_68_94 ();
 sg13g2_fill_1 FILLER_68_110 ();
 sg13g2_decap_8 FILLER_68_117 ();
 sg13g2_decap_4 FILLER_68_124 ();
 sg13g2_fill_1 FILLER_68_128 ();
 sg13g2_fill_1 FILLER_68_155 ();
 sg13g2_fill_2 FILLER_68_165 ();
 sg13g2_fill_2 FILLER_68_180 ();
 sg13g2_fill_1 FILLER_68_182 ();
 sg13g2_fill_1 FILLER_68_193 ();
 sg13g2_fill_1 FILLER_68_253 ();
 sg13g2_decap_8 FILLER_68_332 ();
 sg13g2_fill_2 FILLER_68_339 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_fill_2 FILLER_68_364 ();
 sg13g2_decap_8 FILLER_68_378 ();
 sg13g2_decap_8 FILLER_68_457 ();
 sg13g2_decap_4 FILLER_68_464 ();
 sg13g2_fill_2 FILLER_68_468 ();
 sg13g2_fill_1 FILLER_68_506 ();
 sg13g2_fill_2 FILLER_68_525 ();
 sg13g2_decap_4 FILLER_68_578 ();
 sg13g2_fill_2 FILLER_68_582 ();
 sg13g2_decap_4 FILLER_68_588 ();
 sg13g2_fill_1 FILLER_68_627 ();
 sg13g2_fill_2 FILLER_68_674 ();
 sg13g2_fill_2 FILLER_68_704 ();
 sg13g2_fill_1 FILLER_68_706 ();
 sg13g2_decap_8 FILLER_68_735 ();
 sg13g2_decap_8 FILLER_68_742 ();
 sg13g2_fill_1 FILLER_68_749 ();
 sg13g2_fill_1 FILLER_68_801 ();
 sg13g2_fill_2 FILLER_68_838 ();
 sg13g2_fill_1 FILLER_68_864 ();
 sg13g2_fill_2 FILLER_68_910 ();
 sg13g2_fill_1 FILLER_68_957 ();
 sg13g2_fill_2 FILLER_68_976 ();
 sg13g2_decap_8 FILLER_68_1006 ();
 sg13g2_decap_8 FILLER_68_1013 ();
 sg13g2_decap_8 FILLER_68_1025 ();
 sg13g2_fill_1 FILLER_68_1032 ();
 sg13g2_fill_1 FILLER_68_1057 ();
 sg13g2_fill_1 FILLER_68_1075 ();
 sg13g2_fill_2 FILLER_68_1091 ();
 sg13g2_fill_1 FILLER_68_1093 ();
 sg13g2_fill_1 FILLER_68_1103 ();
 sg13g2_fill_1 FILLER_68_1113 ();
 sg13g2_fill_2 FILLER_68_1119 ();
 sg13g2_fill_1 FILLER_68_1121 ();
 sg13g2_fill_1 FILLER_68_1145 ();
 sg13g2_fill_2 FILLER_68_1163 ();
 sg13g2_fill_2 FILLER_68_1201 ();
 sg13g2_fill_1 FILLER_68_1203 ();
 sg13g2_fill_1 FILLER_68_1227 ();
 sg13g2_decap_8 FILLER_68_1238 ();
 sg13g2_fill_1 FILLER_68_1245 ();
 sg13g2_fill_1 FILLER_68_1273 ();
 sg13g2_decap_4 FILLER_68_1278 ();
 sg13g2_fill_1 FILLER_68_1282 ();
 sg13g2_fill_1 FILLER_68_1306 ();
 sg13g2_decap_8 FILLER_68_1324 ();
 sg13g2_fill_1 FILLER_68_1331 ();
 sg13g2_fill_1 FILLER_68_1358 ();
 sg13g2_fill_1 FILLER_68_1368 ();
 sg13g2_decap_8 FILLER_68_1386 ();
 sg13g2_fill_2 FILLER_68_1393 ();
 sg13g2_fill_2 FILLER_68_1417 ();
 sg13g2_fill_1 FILLER_68_1487 ();
 sg13g2_fill_1 FILLER_68_1501 ();
 sg13g2_fill_1 FILLER_68_1535 ();
 sg13g2_decap_8 FILLER_68_1569 ();
 sg13g2_fill_1 FILLER_68_1576 ();
 sg13g2_decap_8 FILLER_68_1581 ();
 sg13g2_decap_8 FILLER_68_1600 ();
 sg13g2_fill_2 FILLER_68_1607 ();
 sg13g2_fill_1 FILLER_68_1609 ();
 sg13g2_fill_2 FILLER_68_1628 ();
 sg13g2_decap_8 FILLER_68_1639 ();
 sg13g2_fill_2 FILLER_68_1651 ();
 sg13g2_fill_2 FILLER_68_1658 ();
 sg13g2_fill_1 FILLER_68_1660 ();
 sg13g2_decap_4 FILLER_68_1679 ();
 sg13g2_decap_8 FILLER_68_1687 ();
 sg13g2_fill_1 FILLER_68_1694 ();
 sg13g2_decap_8 FILLER_68_1704 ();
 sg13g2_decap_8 FILLER_68_1711 ();
 sg13g2_fill_1 FILLER_68_1718 ();
 sg13g2_fill_1 FILLER_68_1732 ();
 sg13g2_decap_4 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_4 ();
 sg13g2_fill_2 FILLER_69_37 ();
 sg13g2_fill_1 FILLER_69_128 ();
 sg13g2_decap_4 FILLER_69_194 ();
 sg13g2_fill_2 FILLER_69_208 ();
 sg13g2_fill_1 FILLER_69_210 ();
 sg13g2_fill_1 FILLER_69_224 ();
 sg13g2_fill_1 FILLER_69_304 ();
 sg13g2_fill_2 FILLER_69_377 ();
 sg13g2_decap_4 FILLER_69_410 ();
 sg13g2_fill_1 FILLER_69_414 ();
 sg13g2_fill_1 FILLER_69_477 ();
 sg13g2_decap_4 FILLER_69_516 ();
 sg13g2_fill_2 FILLER_69_520 ();
 sg13g2_fill_2 FILLER_69_625 ();
 sg13g2_fill_1 FILLER_69_627 ();
 sg13g2_fill_1 FILLER_69_641 ();
 sg13g2_decap_4 FILLER_69_719 ();
 sg13g2_fill_2 FILLER_69_810 ();
 sg13g2_fill_2 FILLER_69_830 ();
 sg13g2_fill_2 FILLER_69_872 ();
 sg13g2_fill_2 FILLER_69_888 ();
 sg13g2_decap_4 FILLER_69_937 ();
 sg13g2_fill_1 FILLER_69_1018 ();
 sg13g2_fill_2 FILLER_69_1059 ();
 sg13g2_fill_2 FILLER_69_1102 ();
 sg13g2_fill_2 FILLER_69_1110 ();
 sg13g2_decap_4 FILLER_69_1177 ();
 sg13g2_fill_2 FILLER_69_1181 ();
 sg13g2_decap_4 FILLER_69_1188 ();
 sg13g2_fill_1 FILLER_69_1209 ();
 sg13g2_fill_1 FILLER_69_1238 ();
 sg13g2_fill_2 FILLER_69_1267 ();
 sg13g2_fill_1 FILLER_69_1282 ();
 sg13g2_decap_4 FILLER_69_1321 ();
 sg13g2_fill_2 FILLER_69_1336 ();
 sg13g2_decap_8 FILLER_69_1375 ();
 sg13g2_fill_2 FILLER_69_1382 ();
 sg13g2_decap_4 FILLER_69_1388 ();
 sg13g2_decap_4 FILLER_69_1425 ();
 sg13g2_fill_2 FILLER_69_1447 ();
 sg13g2_fill_1 FILLER_69_1462 ();
 sg13g2_decap_8 FILLER_69_1472 ();
 sg13g2_decap_4 FILLER_69_1479 ();
 sg13g2_fill_1 FILLER_69_1483 ();
 sg13g2_decap_8 FILLER_69_1502 ();
 sg13g2_fill_2 FILLER_69_1509 ();
 sg13g2_fill_1 FILLER_69_1511 ();
 sg13g2_decap_4 FILLER_69_1516 ();
 sg13g2_fill_1 FILLER_69_1520 ();
 sg13g2_fill_2 FILLER_69_1545 ();
 sg13g2_fill_2 FILLER_69_1551 ();
 sg13g2_fill_1 FILLER_69_1553 ();
 sg13g2_decap_8 FILLER_69_1563 ();
 sg13g2_fill_1 FILLER_69_1570 ();
 sg13g2_decap_8 FILLER_69_1604 ();
 sg13g2_decap_8 FILLER_69_1611 ();
 sg13g2_fill_2 FILLER_69_1618 ();
 sg13g2_fill_2 FILLER_69_1629 ();
 sg13g2_decap_8 FILLER_69_1641 ();
 sg13g2_decap_8 FILLER_69_1666 ();
 sg13g2_fill_1 FILLER_69_1673 ();
 sg13g2_decap_8 FILLER_69_1678 ();
 sg13g2_decap_8 FILLER_69_1685 ();
 sg13g2_decap_8 FILLER_69_1711 ();
 sg13g2_decap_4 FILLER_69_1718 ();
 sg13g2_fill_1 FILLER_69_1722 ();
 sg13g2_decap_4 FILLER_69_1728 ();
 sg13g2_fill_2 FILLER_69_1751 ();
 sg13g2_fill_1 FILLER_69_1753 ();
 sg13g2_fill_1 FILLER_69_1767 ();
 sg13g2_fill_2 FILLER_70_95 ();
 sg13g2_fill_1 FILLER_70_128 ();
 sg13g2_fill_1 FILLER_70_147 ();
 sg13g2_fill_1 FILLER_70_165 ();
 sg13g2_decap_4 FILLER_70_170 ();
 sg13g2_fill_2 FILLER_70_174 ();
 sg13g2_decap_8 FILLER_70_200 ();
 sg13g2_fill_2 FILLER_70_211 ();
 sg13g2_fill_1 FILLER_70_213 ();
 sg13g2_fill_2 FILLER_70_219 ();
 sg13g2_fill_2 FILLER_70_256 ();
 sg13g2_fill_2 FILLER_70_347 ();
 sg13g2_decap_4 FILLER_70_365 ();
 sg13g2_fill_1 FILLER_70_369 ();
 sg13g2_fill_2 FILLER_70_390 ();
 sg13g2_fill_1 FILLER_70_398 ();
 sg13g2_decap_8 FILLER_70_407 ();
 sg13g2_fill_2 FILLER_70_414 ();
 sg13g2_fill_1 FILLER_70_416 ();
 sg13g2_fill_2 FILLER_70_430 ();
 sg13g2_fill_1 FILLER_70_432 ();
 sg13g2_fill_2 FILLER_70_448 ();
 sg13g2_fill_1 FILLER_70_450 ();
 sg13g2_fill_2 FILLER_70_464 ();
 sg13g2_decap_4 FILLER_70_505 ();
 sg13g2_fill_1 FILLER_70_509 ();
 sg13g2_fill_2 FILLER_70_523 ();
 sg13g2_fill_1 FILLER_70_525 ();
 sg13g2_decap_4 FILLER_70_534 ();
 sg13g2_fill_1 FILLER_70_538 ();
 sg13g2_fill_1 FILLER_70_603 ();
 sg13g2_fill_1 FILLER_70_627 ();
 sg13g2_fill_2 FILLER_70_691 ();
 sg13g2_fill_1 FILLER_70_698 ();
 sg13g2_fill_1 FILLER_70_727 ();
 sg13g2_decap_4 FILLER_70_797 ();
 sg13g2_fill_1 FILLER_70_801 ();
 sg13g2_fill_2 FILLER_70_832 ();
 sg13g2_fill_1 FILLER_70_834 ();
 sg13g2_fill_2 FILLER_70_848 ();
 sg13g2_fill_2 FILLER_70_854 ();
 sg13g2_fill_2 FILLER_70_865 ();
 sg13g2_decap_4 FILLER_70_900 ();
 sg13g2_fill_2 FILLER_70_920 ();
 sg13g2_fill_2 FILLER_70_974 ();
 sg13g2_fill_2 FILLER_70_989 ();
 sg13g2_decap_8 FILLER_70_1030 ();
 sg13g2_decap_8 FILLER_70_1037 ();
 sg13g2_fill_2 FILLER_70_1044 ();
 sg13g2_fill_2 FILLER_70_1064 ();
 sg13g2_fill_1 FILLER_70_1116 ();
 sg13g2_fill_2 FILLER_70_1145 ();
 sg13g2_fill_2 FILLER_70_1165 ();
 sg13g2_fill_1 FILLER_70_1167 ();
 sg13g2_fill_2 FILLER_70_1182 ();
 sg13g2_fill_2 FILLER_70_1216 ();
 sg13g2_fill_1 FILLER_70_1218 ();
 sg13g2_fill_2 FILLER_70_1326 ();
 sg13g2_fill_1 FILLER_70_1328 ();
 sg13g2_fill_1 FILLER_70_1461 ();
 sg13g2_decap_4 FILLER_70_1479 ();
 sg13g2_fill_2 FILLER_70_1483 ();
 sg13g2_decap_8 FILLER_70_1502 ();
 sg13g2_fill_2 FILLER_70_1509 ();
 sg13g2_fill_1 FILLER_70_1511 ();
 sg13g2_fill_1 FILLER_70_1517 ();
 sg13g2_fill_1 FILLER_70_1531 ();
 sg13g2_fill_2 FILLER_70_1565 ();
 sg13g2_fill_1 FILLER_70_1567 ();
 sg13g2_decap_4 FILLER_70_1585 ();
 sg13g2_fill_2 FILLER_70_1589 ();
 sg13g2_decap_8 FILLER_70_1604 ();
 sg13g2_decap_8 FILLER_70_1611 ();
 sg13g2_fill_2 FILLER_70_1623 ();
 sg13g2_fill_1 FILLER_70_1625 ();
 sg13g2_fill_1 FILLER_70_1660 ();
 sg13g2_fill_2 FILLER_70_1686 ();
 sg13g2_decap_8 FILLER_70_1717 ();
 sg13g2_decap_4 FILLER_70_1724 ();
 sg13g2_decap_4 FILLER_70_1762 ();
 sg13g2_fill_2 FILLER_70_1766 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_9 ();
 sg13g2_decap_4 FILLER_71_14 ();
 sg13g2_fill_2 FILLER_71_18 ();
 sg13g2_fill_1 FILLER_71_130 ();
 sg13g2_fill_2 FILLER_71_144 ();
 sg13g2_decap_8 FILLER_71_167 ();
 sg13g2_fill_2 FILLER_71_200 ();
 sg13g2_fill_2 FILLER_71_222 ();
 sg13g2_fill_1 FILLER_71_224 ();
 sg13g2_fill_2 FILLER_71_243 ();
 sg13g2_fill_1 FILLER_71_258 ();
 sg13g2_fill_2 FILLER_71_291 ();
 sg13g2_fill_2 FILLER_71_337 ();
 sg13g2_decap_8 FILLER_71_367 ();
 sg13g2_decap_8 FILLER_71_374 ();
 sg13g2_fill_2 FILLER_71_381 ();
 sg13g2_fill_2 FILLER_71_499 ();
 sg13g2_fill_1 FILLER_71_501 ();
 sg13g2_fill_2 FILLER_71_508 ();
 sg13g2_fill_1 FILLER_71_510 ();
 sg13g2_fill_2 FILLER_71_539 ();
 sg13g2_fill_1 FILLER_71_541 ();
 sg13g2_fill_1 FILLER_71_574 ();
 sg13g2_fill_2 FILLER_71_617 ();
 sg13g2_fill_1 FILLER_71_619 ();
 sg13g2_fill_2 FILLER_71_645 ();
 sg13g2_fill_1 FILLER_71_647 ();
 sg13g2_fill_1 FILLER_71_672 ();
 sg13g2_decap_8 FILLER_71_705 ();
 sg13g2_decap_8 FILLER_71_712 ();
 sg13g2_decap_4 FILLER_71_719 ();
 sg13g2_fill_1 FILLER_71_723 ();
 sg13g2_fill_1 FILLER_71_729 ();
 sg13g2_decap_8 FILLER_71_786 ();
 sg13g2_decap_8 FILLER_71_793 ();
 sg13g2_fill_1 FILLER_71_800 ();
 sg13g2_decap_4 FILLER_71_843 ();
 sg13g2_decap_4 FILLER_71_852 ();
 sg13g2_fill_1 FILLER_71_856 ();
 sg13g2_fill_2 FILLER_71_877 ();
 sg13g2_decap_8 FILLER_71_910 ();
 sg13g2_fill_2 FILLER_71_917 ();
 sg13g2_fill_2 FILLER_71_928 ();
 sg13g2_fill_1 FILLER_71_943 ();
 sg13g2_fill_2 FILLER_71_949 ();
 sg13g2_fill_1 FILLER_71_951 ();
 sg13g2_fill_2 FILLER_71_965 ();
 sg13g2_fill_1 FILLER_71_967 ();
 sg13g2_fill_1 FILLER_71_973 ();
 sg13g2_fill_2 FILLER_71_987 ();
 sg13g2_fill_1 FILLER_71_989 ();
 sg13g2_fill_2 FILLER_71_999 ();
 sg13g2_decap_8 FILLER_71_1006 ();
 sg13g2_fill_2 FILLER_71_1013 ();
 sg13g2_fill_2 FILLER_71_1020 ();
 sg13g2_fill_1 FILLER_71_1022 ();
 sg13g2_fill_2 FILLER_71_1063 ();
 sg13g2_fill_1 FILLER_71_1065 ();
 sg13g2_fill_2 FILLER_71_1079 ();
 sg13g2_fill_2 FILLER_71_1109 ();
 sg13g2_fill_1 FILLER_71_1111 ();
 sg13g2_fill_1 FILLER_71_1142 ();
 sg13g2_fill_1 FILLER_71_1174 ();
 sg13g2_fill_2 FILLER_71_1203 ();
 sg13g2_fill_2 FILLER_71_1248 ();
 sg13g2_fill_1 FILLER_71_1250 ();
 sg13g2_fill_1 FILLER_71_1274 ();
 sg13g2_fill_2 FILLER_71_1311 ();
 sg13g2_fill_1 FILLER_71_1386 ();
 sg13g2_decap_8 FILLER_71_1444 ();
 sg13g2_fill_2 FILLER_71_1451 ();
 sg13g2_fill_1 FILLER_71_1453 ();
 sg13g2_fill_2 FILLER_71_1474 ();
 sg13g2_decap_4 FILLER_71_1485 ();
 sg13g2_fill_1 FILLER_71_1489 ();
 sg13g2_decap_4 FILLER_71_1500 ();
 sg13g2_fill_2 FILLER_71_1504 ();
 sg13g2_fill_2 FILLER_71_1512 ();
 sg13g2_fill_1 FILLER_71_1519 ();
 sg13g2_decap_8 FILLER_71_1525 ();
 sg13g2_decap_4 FILLER_71_1532 ();
 sg13g2_fill_2 FILLER_71_1549 ();
 sg13g2_fill_2 FILLER_71_1560 ();
 sg13g2_fill_2 FILLER_71_1568 ();
 sg13g2_decap_4 FILLER_71_1688 ();
 sg13g2_fill_2 FILLER_71_1692 ();
 sg13g2_fill_2 FILLER_71_1698 ();
 sg13g2_fill_1 FILLER_71_1700 ();
 sg13g2_fill_1 FILLER_71_1707 ();
 sg13g2_decap_4 FILLER_71_1712 ();
 sg13g2_decap_4 FILLER_71_1729 ();
 sg13g2_decap_4 FILLER_72_0 ();
 sg13g2_fill_1 FILLER_72_4 ();
 sg13g2_decap_8 FILLER_72_9 ();
 sg13g2_decap_8 FILLER_72_16 ();
 sg13g2_fill_1 FILLER_72_50 ();
 sg13g2_decap_4 FILLER_72_69 ();
 sg13g2_fill_1 FILLER_72_73 ();
 sg13g2_fill_1 FILLER_72_80 ();
 sg13g2_fill_1 FILLER_72_157 ();
 sg13g2_fill_2 FILLER_72_199 ();
 sg13g2_fill_1 FILLER_72_201 ();
 sg13g2_fill_2 FILLER_72_206 ();
 sg13g2_fill_2 FILLER_72_240 ();
 sg13g2_fill_1 FILLER_72_260 ();
 sg13g2_fill_1 FILLER_72_351 ();
 sg13g2_decap_4 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_372 ();
 sg13g2_fill_2 FILLER_72_379 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_72_434 ();
 sg13g2_fill_2 FILLER_72_441 ();
 sg13g2_fill_1 FILLER_72_456 ();
 sg13g2_fill_2 FILLER_72_466 ();
 sg13g2_decap_8 FILLER_72_484 ();
 sg13g2_decap_4 FILLER_72_491 ();
 sg13g2_fill_2 FILLER_72_495 ();
 sg13g2_fill_2 FILLER_72_519 ();
 sg13g2_fill_1 FILLER_72_521 ();
 sg13g2_decap_8 FILLER_72_531 ();
 sg13g2_decap_4 FILLER_72_547 ();
 sg13g2_fill_1 FILLER_72_576 ();
 sg13g2_fill_2 FILLER_72_591 ();
 sg13g2_fill_1 FILLER_72_593 ();
 sg13g2_fill_1 FILLER_72_604 ();
 sg13g2_fill_2 FILLER_72_609 ();
 sg13g2_fill_1 FILLER_72_611 ();
 sg13g2_fill_2 FILLER_72_661 ();
 sg13g2_fill_1 FILLER_72_668 ();
 sg13g2_fill_1 FILLER_72_719 ();
 sg13g2_decap_4 FILLER_72_761 ();
 sg13g2_fill_1 FILLER_72_765 ();
 sg13g2_fill_2 FILLER_72_807 ();
 sg13g2_fill_1 FILLER_72_809 ();
 sg13g2_fill_2 FILLER_72_827 ();
 sg13g2_fill_1 FILLER_72_829 ();
 sg13g2_fill_2 FILLER_72_981 ();
 sg13g2_decap_4 FILLER_72_1015 ();
 sg13g2_fill_1 FILLER_72_1019 ();
 sg13g2_decap_8 FILLER_72_1033 ();
 sg13g2_decap_4 FILLER_72_1040 ();
 sg13g2_fill_2 FILLER_72_1044 ();
 sg13g2_fill_1 FILLER_72_1059 ();
 sg13g2_fill_2 FILLER_72_1102 ();
 sg13g2_fill_2 FILLER_72_1145 ();
 sg13g2_fill_2 FILLER_72_1166 ();
 sg13g2_fill_1 FILLER_72_1168 ();
 sg13g2_fill_1 FILLER_72_1182 ();
 sg13g2_fill_1 FILLER_72_1214 ();
 sg13g2_fill_2 FILLER_72_1234 ();
 sg13g2_fill_1 FILLER_72_1255 ();
 sg13g2_fill_1 FILLER_72_1275 ();
 sg13g2_fill_2 FILLER_72_1297 ();
 sg13g2_fill_1 FILLER_72_1299 ();
 sg13g2_fill_1 FILLER_72_1316 ();
 sg13g2_fill_2 FILLER_72_1323 ();
 sg13g2_fill_1 FILLER_72_1368 ();
 sg13g2_fill_2 FILLER_72_1397 ();
 sg13g2_fill_1 FILLER_72_1399 ();
 sg13g2_decap_4 FILLER_72_1423 ();
 sg13g2_decap_4 FILLER_72_1468 ();
 sg13g2_fill_2 FILLER_72_1476 ();
 sg13g2_fill_2 FILLER_72_1482 ();
 sg13g2_fill_1 FILLER_72_1484 ();
 sg13g2_fill_2 FILLER_72_1503 ();
 sg13g2_fill_1 FILLER_72_1505 ();
 sg13g2_fill_1 FILLER_72_1514 ();
 sg13g2_decap_4 FILLER_72_1519 ();
 sg13g2_fill_1 FILLER_72_1523 ();
 sg13g2_decap_8 FILLER_72_1548 ();
 sg13g2_decap_4 FILLER_72_1555 ();
 sg13g2_decap_8 FILLER_72_1595 ();
 sg13g2_decap_4 FILLER_72_1602 ();
 sg13g2_fill_1 FILLER_72_1631 ();
 sg13g2_decap_4 FILLER_72_1642 ();
 sg13g2_fill_1 FILLER_72_1696 ();
 sg13g2_decap_4 FILLER_72_1764 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_9 ();
 sg13g2_decap_4 FILLER_73_37 ();
 sg13g2_fill_2 FILLER_73_54 ();
 sg13g2_fill_1 FILLER_73_56 ();
 sg13g2_fill_1 FILLER_73_105 ();
 sg13g2_fill_2 FILLER_73_111 ();
 sg13g2_fill_2 FILLER_73_122 ();
 sg13g2_decap_4 FILLER_73_175 ();
 sg13g2_fill_1 FILLER_73_179 ();
 sg13g2_fill_2 FILLER_73_196 ();
 sg13g2_fill_1 FILLER_73_198 ();
 sg13g2_fill_2 FILLER_73_252 ();
 sg13g2_fill_1 FILLER_73_267 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_315 ();
 sg13g2_decap_4 FILLER_73_355 ();
 sg13g2_fill_2 FILLER_73_399 ();
 sg13g2_fill_1 FILLER_73_401 ();
 sg13g2_fill_2 FILLER_73_415 ();
 sg13g2_fill_1 FILLER_73_417 ();
 sg13g2_decap_8 FILLER_73_433 ();
 sg13g2_fill_2 FILLER_73_440 ();
 sg13g2_fill_1 FILLER_73_442 ();
 sg13g2_fill_2 FILLER_73_483 ();
 sg13g2_fill_1 FILLER_73_485 ();
 sg13g2_decap_4 FILLER_73_496 ();
 sg13g2_decap_4 FILLER_73_561 ();
 sg13g2_fill_2 FILLER_73_565 ();
 sg13g2_fill_2 FILLER_73_594 ();
 sg13g2_fill_1 FILLER_73_627 ();
 sg13g2_fill_2 FILLER_73_660 ();
 sg13g2_fill_1 FILLER_73_662 ();
 sg13g2_fill_2 FILLER_73_702 ();
 sg13g2_fill_1 FILLER_73_704 ();
 sg13g2_fill_2 FILLER_73_732 ();
 sg13g2_decap_4 FILLER_73_747 ();
 sg13g2_fill_2 FILLER_73_751 ();
 sg13g2_fill_1 FILLER_73_771 ();
 sg13g2_fill_1 FILLER_73_797 ();
 sg13g2_fill_1 FILLER_73_807 ();
 sg13g2_fill_2 FILLER_73_840 ();
 sg13g2_fill_1 FILLER_73_861 ();
 sg13g2_decap_8 FILLER_73_907 ();
 sg13g2_fill_2 FILLER_73_914 ();
 sg13g2_fill_1 FILLER_73_916 ();
 sg13g2_fill_1 FILLER_73_935 ();
 sg13g2_fill_2 FILLER_73_972 ();
 sg13g2_decap_8 FILLER_73_1022 ();
 sg13g2_fill_1 FILLER_73_1029 ();
 sg13g2_fill_2 FILLER_73_1062 ();
 sg13g2_fill_1 FILLER_73_1073 ();
 sg13g2_fill_2 FILLER_73_1087 ();
 sg13g2_fill_2 FILLER_73_1107 ();
 sg13g2_fill_1 FILLER_73_1109 ();
 sg13g2_fill_1 FILLER_73_1131 ();
 sg13g2_fill_1 FILLER_73_1181 ();
 sg13g2_fill_1 FILLER_73_1197 ();
 sg13g2_fill_2 FILLER_73_1277 ();
 sg13g2_fill_2 FILLER_73_1309 ();
 sg13g2_fill_1 FILLER_73_1311 ();
 sg13g2_fill_2 FILLER_73_1321 ();
 sg13g2_fill_1 FILLER_73_1323 ();
 sg13g2_fill_2 FILLER_73_1329 ();
 sg13g2_fill_2 FILLER_73_1341 ();
 sg13g2_fill_2 FILLER_73_1383 ();
 sg13g2_fill_2 FILLER_73_1404 ();
 sg13g2_fill_1 FILLER_73_1406 ();
 sg13g2_fill_2 FILLER_73_1412 ();
 sg13g2_decap_4 FILLER_73_1450 ();
 sg13g2_fill_1 FILLER_73_1454 ();
 sg13g2_fill_1 FILLER_73_1460 ();
 sg13g2_decap_4 FILLER_73_1474 ();
 sg13g2_fill_2 FILLER_73_1478 ();
 sg13g2_fill_2 FILLER_73_1508 ();
 sg13g2_fill_2 FILLER_73_1528 ();
 sg13g2_decap_8 FILLER_73_1535 ();
 sg13g2_fill_2 FILLER_73_1542 ();
 sg13g2_decap_8 FILLER_73_1550 ();
 sg13g2_fill_2 FILLER_73_1557 ();
 sg13g2_fill_1 FILLER_73_1568 ();
 sg13g2_decap_4 FILLER_73_1577 ();
 sg13g2_fill_2 FILLER_73_1590 ();
 sg13g2_fill_2 FILLER_73_1619 ();
 sg13g2_fill_2 FILLER_73_1658 ();
 sg13g2_fill_1 FILLER_73_1660 ();
 sg13g2_fill_2 FILLER_73_1668 ();
 sg13g2_fill_1 FILLER_73_1679 ();
 sg13g2_fill_1 FILLER_73_1695 ();
 sg13g2_fill_1 FILLER_73_1702 ();
 sg13g2_fill_2 FILLER_73_1706 ();
 sg13g2_fill_2 FILLER_73_1712 ();
 sg13g2_decap_8 FILLER_73_1723 ();
 sg13g2_decap_8 FILLER_73_1730 ();
 sg13g2_fill_2 FILLER_73_1737 ();
 sg13g2_fill_1 FILLER_73_1739 ();
 sg13g2_decap_4 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_4 ();
 sg13g2_fill_1 FILLER_74_32 ();
 sg13g2_fill_2 FILLER_74_47 ();
 sg13g2_fill_1 FILLER_74_49 ();
 sg13g2_fill_1 FILLER_74_60 ();
 sg13g2_decap_4 FILLER_74_69 ();
 sg13g2_fill_1 FILLER_74_73 ();
 sg13g2_fill_2 FILLER_74_96 ();
 sg13g2_fill_1 FILLER_74_259 ();
 sg13g2_decap_4 FILLER_74_349 ();
 sg13g2_fill_1 FILLER_74_353 ();
 sg13g2_fill_1 FILLER_74_381 ();
 sg13g2_fill_2 FILLER_74_413 ();
 sg13g2_fill_1 FILLER_74_415 ();
 sg13g2_decap_8 FILLER_74_435 ();
 sg13g2_decap_4 FILLER_74_442 ();
 sg13g2_fill_1 FILLER_74_446 ();
 sg13g2_fill_2 FILLER_74_465 ();
 sg13g2_fill_1 FILLER_74_467 ();
 sg13g2_fill_2 FILLER_74_473 ();
 sg13g2_fill_2 FILLER_74_484 ();
 sg13g2_fill_1 FILLER_74_486 ();
 sg13g2_fill_2 FILLER_74_515 ();
 sg13g2_fill_2 FILLER_74_530 ();
 sg13g2_fill_1 FILLER_74_532 ();
 sg13g2_fill_1 FILLER_74_537 ();
 sg13g2_fill_2 FILLER_74_551 ();
 sg13g2_decap_8 FILLER_74_559 ();
 sg13g2_fill_2 FILLER_74_566 ();
 sg13g2_decap_8 FILLER_74_576 ();
 sg13g2_fill_2 FILLER_74_583 ();
 sg13g2_decap_4 FILLER_74_653 ();
 sg13g2_fill_2 FILLER_74_657 ();
 sg13g2_fill_2 FILLER_74_785 ();
 sg13g2_fill_2 FILLER_74_812 ();
 sg13g2_fill_2 FILLER_74_831 ();
 sg13g2_fill_1 FILLER_74_849 ();
 sg13g2_decap_4 FILLER_74_855 ();
 sg13g2_fill_2 FILLER_74_859 ();
 sg13g2_decap_4 FILLER_74_885 ();
 sg13g2_decap_4 FILLER_74_898 ();
 sg13g2_fill_1 FILLER_74_902 ();
 sg13g2_fill_2 FILLER_74_938 ();
 sg13g2_fill_2 FILLER_74_949 ();
 sg13g2_fill_1 FILLER_74_951 ();
 sg13g2_fill_2 FILLER_74_997 ();
 sg13g2_fill_2 FILLER_74_1088 ();
 sg13g2_fill_1 FILLER_74_1090 ();
 sg13g2_fill_1 FILLER_74_1133 ();
 sg13g2_fill_2 FILLER_74_1171 ();
 sg13g2_fill_1 FILLER_74_1173 ();
 sg13g2_fill_2 FILLER_74_1214 ();
 sg13g2_fill_1 FILLER_74_1216 ();
 sg13g2_fill_1 FILLER_74_1226 ();
 sg13g2_fill_2 FILLER_74_1246 ();
 sg13g2_fill_1 FILLER_74_1330 ();
 sg13g2_fill_1 FILLER_74_1403 ();
 sg13g2_fill_1 FILLER_74_1434 ();
 sg13g2_decap_4 FILLER_74_1451 ();
 sg13g2_decap_8 FILLER_74_1478 ();
 sg13g2_fill_2 FILLER_74_1490 ();
 sg13g2_fill_1 FILLER_74_1492 ();
 sg13g2_decap_8 FILLER_74_1503 ();
 sg13g2_decap_4 FILLER_74_1510 ();
 sg13g2_fill_2 FILLER_74_1514 ();
 sg13g2_fill_1 FILLER_74_1533 ();
 sg13g2_decap_4 FILLER_74_1539 ();
 sg13g2_decap_8 FILLER_74_1552 ();
 sg13g2_fill_1 FILLER_74_1559 ();
 sg13g2_fill_2 FILLER_74_1569 ();
 sg13g2_fill_1 FILLER_74_1571 ();
 sg13g2_decap_8 FILLER_74_1577 ();
 sg13g2_fill_2 FILLER_74_1601 ();
 sg13g2_decap_8 FILLER_74_1616 ();
 sg13g2_fill_1 FILLER_74_1623 ();
 sg13g2_decap_4 FILLER_74_1627 ();
 sg13g2_fill_2 FILLER_74_1631 ();
 sg13g2_decap_8 FILLER_74_1646 ();
 sg13g2_decap_8 FILLER_74_1653 ();
 sg13g2_fill_1 FILLER_74_1660 ();
 sg13g2_decap_4 FILLER_74_1689 ();
 sg13g2_fill_1 FILLER_74_1693 ();
 sg13g2_fill_2 FILLER_74_1701 ();
 sg13g2_decap_4 FILLER_74_1731 ();
 sg13g2_decap_4 FILLER_74_1742 ();
 sg13g2_decap_4 FILLER_74_1750 ();
 sg13g2_fill_2 FILLER_74_1754 ();
 sg13g2_fill_2 FILLER_74_1765 ();
 sg13g2_fill_1 FILLER_74_1767 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_fill_2 FILLER_75_51 ();
 sg13g2_fill_1 FILLER_75_66 ();
 sg13g2_fill_2 FILLER_75_156 ();
 sg13g2_fill_2 FILLER_75_162 ();
 sg13g2_fill_2 FILLER_75_173 ();
 sg13g2_fill_1 FILLER_75_185 ();
 sg13g2_fill_1 FILLER_75_241 ();
 sg13g2_fill_2 FILLER_75_296 ();
 sg13g2_fill_2 FILLER_75_378 ();
 sg13g2_fill_2 FILLER_75_421 ();
 sg13g2_fill_1 FILLER_75_423 ();
 sg13g2_fill_2 FILLER_75_461 ();
 sg13g2_fill_2 FILLER_75_470 ();
 sg13g2_fill_1 FILLER_75_472 ();
 sg13g2_decap_8 FILLER_75_480 ();
 sg13g2_fill_2 FILLER_75_487 ();
 sg13g2_fill_1 FILLER_75_489 ();
 sg13g2_fill_2 FILLER_75_502 ();
 sg13g2_fill_1 FILLER_75_504 ();
 sg13g2_decap_4 FILLER_75_522 ();
 sg13g2_fill_2 FILLER_75_526 ();
 sg13g2_fill_2 FILLER_75_565 ();
 sg13g2_fill_2 FILLER_75_598 ();
 sg13g2_fill_1 FILLER_75_600 ();
 sg13g2_decap_4 FILLER_75_669 ();
 sg13g2_fill_2 FILLER_75_673 ();
 sg13g2_fill_1 FILLER_75_688 ();
 sg13g2_fill_2 FILLER_75_710 ();
 sg13g2_fill_1 FILLER_75_712 ();
 sg13g2_fill_2 FILLER_75_721 ();
 sg13g2_decap_4 FILLER_75_746 ();
 sg13g2_fill_2 FILLER_75_750 ();
 sg13g2_decap_8 FILLER_75_756 ();
 sg13g2_fill_1 FILLER_75_763 ();
 sg13g2_fill_2 FILLER_75_803 ();
 sg13g2_fill_1 FILLER_75_818 ();
 sg13g2_fill_2 FILLER_75_825 ();
 sg13g2_fill_2 FILLER_75_850 ();
 sg13g2_fill_1 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_861 ();
 sg13g2_fill_1 FILLER_75_882 ();
 sg13g2_fill_1 FILLER_75_889 ();
 sg13g2_fill_2 FILLER_75_927 ();
 sg13g2_fill_1 FILLER_75_957 ();
 sg13g2_fill_2 FILLER_75_976 ();
 sg13g2_fill_1 FILLER_75_978 ();
 sg13g2_fill_2 FILLER_75_1038 ();
 sg13g2_fill_1 FILLER_75_1040 ();
 sg13g2_fill_1 FILLER_75_1050 ();
 sg13g2_fill_2 FILLER_75_1091 ();
 sg13g2_fill_1 FILLER_75_1093 ();
 sg13g2_fill_1 FILLER_75_1142 ();
 sg13g2_fill_1 FILLER_75_1179 ();
 sg13g2_fill_1 FILLER_75_1215 ();
 sg13g2_fill_2 FILLER_75_1242 ();
 sg13g2_fill_2 FILLER_75_1248 ();
 sg13g2_fill_2 FILLER_75_1290 ();
 sg13g2_fill_1 FILLER_75_1292 ();
 sg13g2_decap_4 FILLER_75_1331 ();
 sg13g2_decap_4 FILLER_75_1343 ();
 sg13g2_fill_1 FILLER_75_1347 ();
 sg13g2_decap_8 FILLER_75_1352 ();
 sg13g2_decap_4 FILLER_75_1359 ();
 sg13g2_fill_1 FILLER_75_1363 ();
 sg13g2_fill_1 FILLER_75_1373 ();
 sg13g2_fill_1 FILLER_75_1392 ();
 sg13g2_fill_2 FILLER_75_1417 ();
 sg13g2_fill_1 FILLER_75_1419 ();
 sg13g2_fill_2 FILLER_75_1430 ();
 sg13g2_fill_1 FILLER_75_1432 ();
 sg13g2_fill_1 FILLER_75_1439 ();
 sg13g2_decap_4 FILLER_75_1473 ();
 sg13g2_decap_4 FILLER_75_1487 ();
 sg13g2_fill_1 FILLER_75_1501 ();
 sg13g2_decap_4 FILLER_75_1507 ();
 sg13g2_fill_2 FILLER_75_1511 ();
 sg13g2_decap_8 FILLER_75_1528 ();
 sg13g2_fill_1 FILLER_75_1535 ();
 sg13g2_fill_1 FILLER_75_1546 ();
 sg13g2_decap_4 FILLER_75_1559 ();
 sg13g2_fill_2 FILLER_75_1588 ();
 sg13g2_decap_4 FILLER_75_1660 ();
 sg13g2_fill_2 FILLER_75_1664 ();
 sg13g2_decap_8 FILLER_75_1670 ();
 sg13g2_fill_2 FILLER_75_1677 ();
 sg13g2_fill_2 FILLER_75_1683 ();
 sg13g2_fill_2 FILLER_75_1690 ();
 sg13g2_decap_4 FILLER_75_1729 ();
 sg13g2_fill_1 FILLER_75_1738 ();
 sg13g2_fill_1 FILLER_75_1767 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_52 ();
 sg13g2_fill_2 FILLER_76_58 ();
 sg13g2_fill_1 FILLER_76_60 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_fill_1 FILLER_76_141 ();
 sg13g2_fill_1 FILLER_76_151 ();
 sg13g2_fill_2 FILLER_76_155 ();
 sg13g2_fill_1 FILLER_76_157 ();
 sg13g2_fill_1 FILLER_76_167 ();
 sg13g2_fill_1 FILLER_76_172 ();
 sg13g2_fill_1 FILLER_76_190 ();
 sg13g2_fill_1 FILLER_76_220 ();
 sg13g2_fill_1 FILLER_76_279 ();
 sg13g2_fill_1 FILLER_76_284 ();
 sg13g2_fill_1 FILLER_76_324 ();
 sg13g2_decap_8 FILLER_76_338 ();
 sg13g2_fill_2 FILLER_76_345 ();
 sg13g2_decap_8 FILLER_76_351 ();
 sg13g2_decap_8 FILLER_76_443 ();
 sg13g2_decap_4 FILLER_76_450 ();
 sg13g2_fill_1 FILLER_76_454 ();
 sg13g2_fill_1 FILLER_76_469 ();
 sg13g2_fill_2 FILLER_76_505 ();
 sg13g2_fill_1 FILLER_76_507 ();
 sg13g2_decap_4 FILLER_76_524 ();
 sg13g2_fill_1 FILLER_76_528 ();
 sg13g2_fill_2 FILLER_76_585 ();
 sg13g2_fill_2 FILLER_76_597 ();
 sg13g2_decap_4 FILLER_76_612 ();
 sg13g2_fill_2 FILLER_76_616 ();
 sg13g2_fill_1 FILLER_76_641 ();
 sg13g2_fill_1 FILLER_76_651 ();
 sg13g2_fill_1 FILLER_76_656 ();
 sg13g2_fill_1 FILLER_76_670 ();
 sg13g2_fill_2 FILLER_76_740 ();
 sg13g2_fill_1 FILLER_76_742 ();
 sg13g2_fill_1 FILLER_76_752 ();
 sg13g2_decap_8 FILLER_76_765 ();
 sg13g2_fill_1 FILLER_76_802 ();
 sg13g2_decap_4 FILLER_76_833 ();
 sg13g2_fill_2 FILLER_76_837 ();
 sg13g2_fill_2 FILLER_76_850 ();
 sg13g2_fill_2 FILLER_76_868 ();
 sg13g2_fill_1 FILLER_76_884 ();
 sg13g2_fill_1 FILLER_76_888 ();
 sg13g2_fill_1 FILLER_76_892 ();
 sg13g2_fill_2 FILLER_76_917 ();
 sg13g2_fill_2 FILLER_76_950 ();
 sg13g2_fill_2 FILLER_76_980 ();
 sg13g2_fill_1 FILLER_76_1017 ();
 sg13g2_fill_2 FILLER_76_1168 ();
 sg13g2_fill_1 FILLER_76_1170 ();
 sg13g2_fill_2 FILLER_76_1199 ();
 sg13g2_fill_2 FILLER_76_1218 ();
 sg13g2_fill_2 FILLER_76_1257 ();
 sg13g2_decap_8 FILLER_76_1341 ();
 sg13g2_decap_8 FILLER_76_1348 ();
 sg13g2_decap_4 FILLER_76_1355 ();
 sg13g2_fill_2 FILLER_76_1359 ();
 sg13g2_fill_2 FILLER_76_1388 ();
 sg13g2_decap_8 FILLER_76_1418 ();
 sg13g2_fill_2 FILLER_76_1425 ();
 sg13g2_fill_1 FILLER_76_1427 ();
 sg13g2_fill_2 FILLER_76_1434 ();
 sg13g2_fill_1 FILLER_76_1436 ();
 sg13g2_fill_2 FILLER_76_1445 ();
 sg13g2_decap_4 FILLER_76_1472 ();
 sg13g2_fill_2 FILLER_76_1476 ();
 sg13g2_decap_8 FILLER_76_1488 ();
 sg13g2_decap_4 FILLER_76_1495 ();
 sg13g2_fill_2 FILLER_76_1530 ();
 sg13g2_fill_1 FILLER_76_1532 ();
 sg13g2_fill_1 FILLER_76_1542 ();
 sg13g2_fill_2 FILLER_76_1553 ();
 sg13g2_fill_1 FILLER_76_1555 ();
 sg13g2_decap_4 FILLER_76_1566 ();
 sg13g2_fill_2 FILLER_76_1570 ();
 sg13g2_fill_2 FILLER_76_1580 ();
 sg13g2_fill_2 FILLER_76_1596 ();
 sg13g2_fill_1 FILLER_76_1607 ();
 sg13g2_fill_1 FILLER_76_1633 ();
 sg13g2_fill_2 FILLER_76_1647 ();
 sg13g2_fill_1 FILLER_76_1649 ();
 sg13g2_decap_4 FILLER_76_1706 ();
 sg13g2_fill_2 FILLER_76_1710 ();
 sg13g2_fill_2 FILLER_76_1741 ();
 sg13g2_fill_1 FILLER_76_1743 ();
 sg13g2_fill_2 FILLER_76_1748 ();
 sg13g2_decap_8 FILLER_76_1759 ();
 sg13g2_fill_2 FILLER_76_1766 ();
 sg13g2_decap_4 FILLER_77_0 ();
 sg13g2_fill_2 FILLER_77_4 ();
 sg13g2_fill_2 FILLER_77_33 ();
 sg13g2_fill_1 FILLER_77_35 ();
 sg13g2_fill_1 FILLER_77_91 ();
 sg13g2_fill_2 FILLER_77_134 ();
 sg13g2_fill_2 FILLER_77_199 ();
 sg13g2_fill_2 FILLER_77_210 ();
 sg13g2_fill_2 FILLER_77_226 ();
 sg13g2_decap_4 FILLER_77_294 ();
 sg13g2_fill_1 FILLER_77_298 ();
 sg13g2_fill_1 FILLER_77_330 ();
 sg13g2_fill_2 FILLER_77_336 ();
 sg13g2_fill_1 FILLER_77_347 ();
 sg13g2_fill_1 FILLER_77_356 ();
 sg13g2_fill_1 FILLER_77_361 ();
 sg13g2_fill_2 FILLER_77_371 ();
 sg13g2_fill_1 FILLER_77_373 ();
 sg13g2_fill_1 FILLER_77_428 ();
 sg13g2_fill_1 FILLER_77_457 ();
 sg13g2_fill_1 FILLER_77_472 ();
 sg13g2_decap_8 FILLER_77_487 ();
 sg13g2_fill_2 FILLER_77_494 ();
 sg13g2_fill_1 FILLER_77_496 ();
 sg13g2_fill_2 FILLER_77_503 ();
 sg13g2_fill_2 FILLER_77_513 ();
 sg13g2_fill_1 FILLER_77_538 ();
 sg13g2_decap_4 FILLER_77_579 ();
 sg13g2_fill_1 FILLER_77_583 ();
 sg13g2_fill_2 FILLER_77_621 ();
 sg13g2_fill_1 FILLER_77_623 ();
 sg13g2_fill_2 FILLER_77_738 ();
 sg13g2_decap_4 FILLER_77_750 ();
 sg13g2_fill_1 FILLER_77_754 ();
 sg13g2_fill_1 FILLER_77_818 ();
 sg13g2_fill_2 FILLER_77_844 ();
 sg13g2_fill_1 FILLER_77_846 ();
 sg13g2_fill_1 FILLER_77_856 ();
 sg13g2_decap_4 FILLER_77_865 ();
 sg13g2_fill_2 FILLER_77_869 ();
 sg13g2_decap_8 FILLER_77_894 ();
 sg13g2_decap_4 FILLER_77_951 ();
 sg13g2_fill_1 FILLER_77_955 ();
 sg13g2_fill_1 FILLER_77_993 ();
 sg13g2_fill_1 FILLER_77_1036 ();
 sg13g2_fill_2 FILLER_77_1069 ();
 sg13g2_fill_1 FILLER_77_1103 ();
 sg13g2_fill_2 FILLER_77_1118 ();
 sg13g2_fill_1 FILLER_77_1198 ();
 sg13g2_fill_1 FILLER_77_1227 ();
 sg13g2_fill_1 FILLER_77_1256 ();
 sg13g2_fill_2 FILLER_77_1280 ();
 sg13g2_fill_1 FILLER_77_1282 ();
 sg13g2_fill_1 FILLER_77_1296 ();
 sg13g2_fill_2 FILLER_77_1325 ();
 sg13g2_fill_1 FILLER_77_1327 ();
 sg13g2_fill_2 FILLER_77_1392 ();
 sg13g2_fill_1 FILLER_77_1394 ();
 sg13g2_fill_2 FILLER_77_1425 ();
 sg13g2_fill_1 FILLER_77_1427 ();
 sg13g2_fill_1 FILLER_77_1434 ();
 sg13g2_decap_8 FILLER_77_1449 ();
 sg13g2_decap_4 FILLER_77_1468 ();
 sg13g2_decap_8 FILLER_77_1487 ();
 sg13g2_decap_4 FILLER_77_1494 ();
 sg13g2_decap_4 FILLER_77_1502 ();
 sg13g2_fill_2 FILLER_77_1506 ();
 sg13g2_decap_8 FILLER_77_1513 ();
 sg13g2_decap_8 FILLER_77_1534 ();
 sg13g2_decap_8 FILLER_77_1545 ();
 sg13g2_fill_2 FILLER_77_1552 ();
 sg13g2_fill_2 FILLER_77_1563 ();
 sg13g2_fill_1 FILLER_77_1565 ();
 sg13g2_fill_2 FILLER_77_1576 ();
 sg13g2_decap_4 FILLER_77_1598 ();
 sg13g2_fill_1 FILLER_77_1602 ();
 sg13g2_decap_8 FILLER_77_1607 ();
 sg13g2_fill_2 FILLER_77_1614 ();
 sg13g2_fill_1 FILLER_77_1616 ();
 sg13g2_decap_8 FILLER_77_1645 ();
 sg13g2_fill_1 FILLER_77_1652 ();
 sg13g2_decap_8 FILLER_77_1666 ();
 sg13g2_decap_8 FILLER_77_1673 ();
 sg13g2_fill_2 FILLER_77_1680 ();
 sg13g2_decap_8 FILLER_77_1686 ();
 sg13g2_decap_8 FILLER_77_1758 ();
 sg13g2_fill_2 FILLER_77_1765 ();
 sg13g2_fill_1 FILLER_77_1767 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_2 ();
 sg13g2_fill_2 FILLER_78_31 ();
 sg13g2_fill_2 FILLER_78_52 ();
 sg13g2_fill_2 FILLER_78_64 ();
 sg13g2_decap_8 FILLER_78_154 ();
 sg13g2_decap_8 FILLER_78_169 ();
 sg13g2_decap_8 FILLER_78_176 ();
 sg13g2_decap_8 FILLER_78_183 ();
 sg13g2_fill_2 FILLER_78_217 ();
 sg13g2_fill_1 FILLER_78_234 ();
 sg13g2_fill_2 FILLER_78_271 ();
 sg13g2_fill_2 FILLER_78_298 ();
 sg13g2_fill_1 FILLER_78_351 ();
 sg13g2_fill_2 FILLER_78_386 ();
 sg13g2_fill_2 FILLER_78_393 ();
 sg13g2_fill_2 FILLER_78_443 ();
 sg13g2_fill_1 FILLER_78_445 ();
 sg13g2_fill_2 FILLER_78_469 ();
 sg13g2_decap_4 FILLER_78_510 ();
 sg13g2_fill_2 FILLER_78_514 ();
 sg13g2_fill_2 FILLER_78_587 ();
 sg13g2_fill_2 FILLER_78_620 ();
 sg13g2_fill_1 FILLER_78_622 ();
 sg13g2_fill_2 FILLER_78_654 ();
 sg13g2_fill_1 FILLER_78_656 ();
 sg13g2_fill_2 FILLER_78_679 ();
 sg13g2_fill_2 FILLER_78_726 ();
 sg13g2_fill_2 FILLER_78_777 ();
 sg13g2_fill_1 FILLER_78_779 ();
 sg13g2_fill_1 FILLER_78_799 ();
 sg13g2_fill_1 FILLER_78_809 ();
 sg13g2_fill_1 FILLER_78_837 ();
 sg13g2_decap_4 FILLER_78_852 ();
 sg13g2_decap_4 FILLER_78_865 ();
 sg13g2_fill_2 FILLER_78_873 ();
 sg13g2_fill_1 FILLER_78_875 ();
 sg13g2_decap_4 FILLER_78_889 ();
 sg13g2_fill_1 FILLER_78_893 ();
 sg13g2_fill_2 FILLER_78_912 ();
 sg13g2_fill_1 FILLER_78_914 ();
 sg13g2_fill_1 FILLER_78_924 ();
 sg13g2_decap_4 FILLER_78_948 ();
 sg13g2_fill_2 FILLER_78_974 ();
 sg13g2_fill_1 FILLER_78_976 ();
 sg13g2_fill_1 FILLER_78_994 ();
 sg13g2_fill_1 FILLER_78_1007 ();
 sg13g2_fill_2 FILLER_78_1041 ();
 sg13g2_fill_1 FILLER_78_1090 ();
 sg13g2_fill_1 FILLER_78_1172 ();
 sg13g2_fill_2 FILLER_78_1224 ();
 sg13g2_fill_2 FILLER_78_1240 ();
 sg13g2_fill_1 FILLER_78_1242 ();
 sg13g2_fill_2 FILLER_78_1373 ();
 sg13g2_fill_1 FILLER_78_1375 ();
 sg13g2_fill_2 FILLER_78_1385 ();
 sg13g2_fill_2 FILLER_78_1414 ();
 sg13g2_fill_1 FILLER_78_1416 ();
 sg13g2_decap_4 FILLER_78_1436 ();
 sg13g2_fill_2 FILLER_78_1446 ();
 sg13g2_fill_1 FILLER_78_1448 ();
 sg13g2_fill_2 FILLER_78_1460 ();
 sg13g2_fill_1 FILLER_78_1462 ();
 sg13g2_fill_2 FILLER_78_1494 ();
 sg13g2_fill_1 FILLER_78_1496 ();
 sg13g2_fill_2 FILLER_78_1537 ();
 sg13g2_fill_1 FILLER_78_1539 ();
 sg13g2_fill_2 FILLER_78_1560 ();
 sg13g2_fill_2 FILLER_78_1575 ();
 sg13g2_decap_8 FILLER_78_1595 ();
 sg13g2_decap_8 FILLER_78_1602 ();
 sg13g2_decap_4 FILLER_78_1616 ();
 sg13g2_fill_2 FILLER_78_1620 ();
 sg13g2_decap_8 FILLER_78_1626 ();
 sg13g2_decap_8 FILLER_78_1633 ();
 sg13g2_decap_8 FILLER_78_1640 ();
 sg13g2_fill_2 FILLER_78_1647 ();
 sg13g2_fill_1 FILLER_78_1705 ();
 sg13g2_fill_2 FILLER_78_1717 ();
 sg13g2_fill_1 FILLER_78_1719 ();
 sg13g2_decap_4 FILLER_78_1729 ();
 sg13g2_fill_1 FILLER_78_1733 ();
 sg13g2_decap_8 FILLER_78_1738 ();
 sg13g2_fill_2 FILLER_78_1745 ();
 sg13g2_fill_1 FILLER_78_1747 ();
 sg13g2_decap_8 FILLER_78_1757 ();
 sg13g2_decap_4 FILLER_78_1764 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_4 FILLER_79_7 ();
 sg13g2_fill_2 FILLER_79_43 ();
 sg13g2_fill_1 FILLER_79_45 ();
 sg13g2_fill_1 FILLER_79_150 ();
 sg13g2_fill_1 FILLER_79_168 ();
 sg13g2_fill_1 FILLER_79_209 ();
 sg13g2_fill_2 FILLER_79_294 ();
 sg13g2_fill_2 FILLER_79_366 ();
 sg13g2_decap_4 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_385 ();
 sg13g2_fill_2 FILLER_79_392 ();
 sg13g2_decap_8 FILLER_79_411 ();
 sg13g2_decap_4 FILLER_79_418 ();
 sg13g2_fill_1 FILLER_79_450 ();
 sg13g2_decap_8 FILLER_79_518 ();
 sg13g2_fill_2 FILLER_79_525 ();
 sg13g2_fill_1 FILLER_79_564 ();
 sg13g2_fill_2 FILLER_79_602 ();
 sg13g2_fill_1 FILLER_79_604 ();
 sg13g2_fill_2 FILLER_79_641 ();
 sg13g2_fill_2 FILLER_79_730 ();
 sg13g2_fill_2 FILLER_79_807 ();
 sg13g2_fill_2 FILLER_79_901 ();
 sg13g2_fill_1 FILLER_79_903 ();
 sg13g2_fill_2 FILLER_79_986 ();
 sg13g2_fill_1 FILLER_79_988 ();
 sg13g2_fill_2 FILLER_79_1017 ();
 sg13g2_fill_1 FILLER_79_1019 ();
 sg13g2_fill_1 FILLER_79_1043 ();
 sg13g2_fill_1 FILLER_79_1088 ();
 sg13g2_fill_1 FILLER_79_1098 ();
 sg13g2_fill_2 FILLER_79_1160 ();
 sg13g2_fill_1 FILLER_79_1175 ();
 sg13g2_fill_1 FILLER_79_1181 ();
 sg13g2_fill_2 FILLER_79_1261 ();
 sg13g2_fill_1 FILLER_79_1304 ();
 sg13g2_fill_1 FILLER_79_1354 ();
 sg13g2_fill_1 FILLER_79_1418 ();
 sg13g2_decap_8 FILLER_79_1452 ();
 sg13g2_fill_2 FILLER_79_1509 ();
 sg13g2_fill_1 FILLER_79_1511 ();
 sg13g2_fill_2 FILLER_79_1526 ();
 sg13g2_fill_1 FILLER_79_1532 ();
 sg13g2_fill_2 FILLER_79_1556 ();
 sg13g2_decap_8 FILLER_79_1576 ();
 sg13g2_fill_1 FILLER_79_1583 ();
 sg13g2_decap_8 FILLER_79_1588 ();
 sg13g2_decap_4 FILLER_79_1595 ();
 sg13g2_decap_8 FILLER_79_1632 ();
 sg13g2_decap_4 FILLER_79_1639 ();
 sg13g2_fill_1 FILLER_79_1643 ();
 sg13g2_fill_2 FILLER_79_1668 ();
 sg13g2_fill_1 FILLER_79_1670 ();
 sg13g2_decap_8 FILLER_79_1680 ();
 sg13g2_decap_8 FILLER_79_1687 ();
 sg13g2_decap_8 FILLER_79_1694 ();
 sg13g2_decap_8 FILLER_79_1701 ();
 sg13g2_decap_8 FILLER_79_1708 ();
 sg13g2_decap_8 FILLER_79_1715 ();
 sg13g2_decap_8 FILLER_79_1722 ();
 sg13g2_decap_8 FILLER_79_1729 ();
 sg13g2_decap_8 FILLER_79_1736 ();
 sg13g2_decap_8 FILLER_79_1743 ();
 sg13g2_decap_8 FILLER_79_1750 ();
 sg13g2_decap_8 FILLER_79_1757 ();
 sg13g2_decap_4 FILLER_79_1764 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_7 ();
 sg13g2_fill_1 FILLER_80_9 ();
 sg13g2_fill_2 FILLER_80_32 ();
 sg13g2_fill_2 FILLER_80_107 ();
 sg13g2_fill_1 FILLER_80_109 ();
 sg13g2_fill_2 FILLER_80_138 ();
 sg13g2_decap_8 FILLER_80_149 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_fill_1 FILLER_80_160 ();
 sg13g2_decap_4 FILLER_80_169 ();
 sg13g2_fill_1 FILLER_80_173 ();
 sg13g2_decap_4 FILLER_80_178 ();
 sg13g2_fill_1 FILLER_80_182 ();
 sg13g2_decap_8 FILLER_80_186 ();
 sg13g2_fill_2 FILLER_80_258 ();
 sg13g2_fill_2 FILLER_80_315 ();
 sg13g2_fill_1 FILLER_80_342 ();
 sg13g2_decap_4 FILLER_80_425 ();
 sg13g2_fill_1 FILLER_80_429 ();
 sg13g2_fill_2 FILLER_80_462 ();
 sg13g2_fill_1 FILLER_80_464 ();
 sg13g2_fill_2 FILLER_80_484 ();
 sg13g2_decap_8 FILLER_80_518 ();
 sg13g2_fill_1 FILLER_80_525 ();
 sg13g2_fill_2 FILLER_80_540 ();
 sg13g2_decap_4 FILLER_80_551 ();
 sg13g2_fill_2 FILLER_80_614 ();
 sg13g2_fill_2 FILLER_80_647 ();
 sg13g2_fill_1 FILLER_80_649 ();
 sg13g2_fill_2 FILLER_80_682 ();
 sg13g2_fill_1 FILLER_80_684 ();
 sg13g2_fill_2 FILLER_80_712 ();
 sg13g2_fill_2 FILLER_80_723 ();
 sg13g2_fill_1 FILLER_80_725 ();
 sg13g2_fill_2 FILLER_80_767 ();
 sg13g2_fill_1 FILLER_80_769 ();
 sg13g2_fill_2 FILLER_80_788 ();
 sg13g2_fill_1 FILLER_80_790 ();
 sg13g2_fill_1 FILLER_80_795 ();
 sg13g2_fill_1 FILLER_80_832 ();
 sg13g2_fill_1 FILLER_80_837 ();
 sg13g2_decap_8 FILLER_80_856 ();
 sg13g2_decap_8 FILLER_80_863 ();
 sg13g2_fill_2 FILLER_80_907 ();
 sg13g2_decap_4 FILLER_80_913 ();
 sg13g2_fill_1 FILLER_80_961 ();
 sg13g2_fill_1 FILLER_80_1012 ();
 sg13g2_fill_2 FILLER_80_1111 ();
 sg13g2_fill_2 FILLER_80_1138 ();
 sg13g2_fill_1 FILLER_80_1140 ();
 sg13g2_fill_2 FILLER_80_1201 ();
 sg13g2_fill_1 FILLER_80_1203 ();
 sg13g2_fill_2 FILLER_80_1232 ();
 sg13g2_fill_1 FILLER_80_1234 ();
 sg13g2_fill_2 FILLER_80_1267 ();
 sg13g2_fill_1 FILLER_80_1269 ();
 sg13g2_fill_2 FILLER_80_1298 ();
 sg13g2_fill_1 FILLER_80_1350 ();
 sg13g2_fill_2 FILLER_80_1359 ();
 sg13g2_decap_4 FILLER_80_1414 ();
 sg13g2_decap_8 FILLER_80_1450 ();
 sg13g2_decap_8 FILLER_80_1457 ();
 sg13g2_decap_8 FILLER_80_1464 ();
 sg13g2_decap_8 FILLER_80_1471 ();
 sg13g2_decap_8 FILLER_80_1478 ();
 sg13g2_decap_8 FILLER_80_1485 ();
 sg13g2_decap_4 FILLER_80_1492 ();
 sg13g2_fill_2 FILLER_80_1496 ();
 sg13g2_decap_4 FILLER_80_1511 ();
 sg13g2_decap_8 FILLER_80_1525 ();
 sg13g2_decap_8 FILLER_80_1532 ();
 sg13g2_decap_4 FILLER_80_1539 ();
 sg13g2_fill_2 FILLER_80_1563 ();
 sg13g2_fill_1 FILLER_80_1565 ();
 sg13g2_decap_8 FILLER_80_1615 ();
 sg13g2_decap_8 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1629 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_decap_8 FILLER_80_1657 ();
 sg13g2_decap_8 FILLER_80_1664 ();
 sg13g2_decap_8 FILLER_80_1671 ();
 sg13g2_decap_8 FILLER_80_1678 ();
 sg13g2_decap_8 FILLER_80_1685 ();
 sg13g2_decap_8 FILLER_80_1692 ();
 sg13g2_decap_8 FILLER_80_1699 ();
 sg13g2_decap_8 FILLER_80_1706 ();
 sg13g2_decap_8 FILLER_80_1713 ();
 sg13g2_decap_8 FILLER_80_1720 ();
 sg13g2_decap_8 FILLER_80_1727 ();
 sg13g2_decap_8 FILLER_80_1734 ();
 sg13g2_decap_8 FILLER_80_1741 ();
 sg13g2_decap_8 FILLER_80_1748 ();
 sg13g2_decap_8 FILLER_80_1755 ();
 sg13g2_decap_4 FILLER_80_1762 ();
 sg13g2_fill_2 FILLER_80_1766 ();
endmodule
