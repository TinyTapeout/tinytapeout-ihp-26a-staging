module tt_um_tomolt_rasterizer (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire clknet_0_clk;
 wire hsync;
 wire \raster.frame_counter[0] ;
 wire \raster.frame_counter[1] ;
 wire \raster.frame_counter[2] ;
 wire \raster.frame_counter[3] ;
 wire \raster.frame_counter[4] ;
 wire \raster.geometry[14] ;
 wire \raster.hpos[0] ;
 wire \raster.hpos[1] ;
 wire \raster.hpos[2] ;
 wire \raster.hpos[3] ;
 wire \raster.hpos[4] ;
 wire \raster.hpos[5] ;
 wire \raster.hpos[6] ;
 wire \raster.hpos[7] ;
 wire \raster.hpos[8] ;
 wire \raster.hpos[9] ;
 wire \raster.hvsync_gen.vpos[0] ;
 wire \raster.hvsync_gen.vpos[1] ;
 wire \raster.hvsync_gen.vpos[2] ;
 wire \raster.hvsync_gen.vpos[3] ;
 wire \raster.hvsync_gen.vpos[4] ;
 wire \raster.hvsync_gen.vpos[5] ;
 wire \raster.hvsync_gen.vpos[6] ;
 wire \raster.hvsync_gen.vpos[7] ;
 wire \raster.hvsync_gen.vpos[8] ;
 wire \raster.hvsync_gen.vpos[9] ;
 wire \raster.hvsync_gen.vsync ;
 wire \raster.tscan.left_err[0] ;
 wire \raster.tscan.left_err[1] ;
 wire \raster.tscan.left_err[2] ;
 wire \raster.tscan.left_err[3] ;
 wire \raster.tscan.left_err[4] ;
 wire \raster.tscan.left_err[5] ;
 wire \raster.tscan.left_err[6] ;
 wire \raster.tscan.left_err[7] ;
 wire \raster.tscan.left_err[8] ;
 wire \raster.tscan.left_err[9] ;
 wire \raster.tscan.left_x[0] ;
 wire \raster.tscan.left_x[1] ;
 wire \raster.tscan.left_x[2] ;
 wire \raster.tscan.left_x[3] ;
 wire \raster.tscan.left_x[4] ;
 wire \raster.tscan.left_x[5] ;
 wire \raster.tscan.left_x[6] ;
 wire \raster.tscan.left_x[7] ;
 wire \raster.tscan.left_x[8] ;
 wire \raster.tscan.left_x[9] ;
 wire \raster.tscan.right_err[0] ;
 wire \raster.tscan.right_err[1] ;
 wire \raster.tscan.right_err[2] ;
 wire \raster.tscan.right_err[3] ;
 wire \raster.tscan.right_err[4] ;
 wire \raster.tscan.right_err[5] ;
 wire \raster.tscan.right_err[6] ;
 wire \raster.tscan.right_err[7] ;
 wire \raster.tscan.right_err[8] ;
 wire \raster.tscan.right_err[9] ;
 wire \raster.tscan.right_x[0] ;
 wire \raster.tscan.right_x[1] ;
 wire \raster.tscan.right_x[2] ;
 wire \raster.tscan.right_x[3] ;
 wire \raster.tscan.right_x[4] ;
 wire \raster.tscan.right_x[5] ;
 wire \raster.tscan.right_x[6] ;
 wire \raster.tscan.right_x[7] ;
 wire \raster.tscan.right_x[8] ;
 wire \raster.tscan.right_x[9] ;
 wire \raster.tscan.state[1] ;
 wire \raster.tscan.state[2] ;
 wire \raster.tscan.state[3] ;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net1;
 wire net2;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;

 sg13g2_inv_2 _0754_ (.Y(\raster.geometry[14] ),
    .A(net155));
 sg13g2_inv_1 _0755_ (.Y(_0071_),
    .A(\raster.hpos[1] ));
 sg13g2_inv_1 _0756_ (.Y(_0072_),
    .A(\raster.hpos[0] ));
 sg13g2_inv_1 _0757_ (.Y(_0073_),
    .A(\raster.hpos[3] ));
 sg13g2_inv_1 _0758_ (.Y(_0074_),
    .A(\raster.hpos[2] ));
 sg13g2_inv_1 _0759_ (.Y(_0075_),
    .A(\raster.hpos[4] ));
 sg13g2_inv_2 _0760_ (.Y(_0076_),
    .A(net112));
 sg13g2_inv_2 _0761_ (.Y(_0077_),
    .A(\raster.hpos[7] ));
 sg13g2_inv_1 _0762_ (.Y(_0078_),
    .A(net166));
 sg13g2_inv_1 _0763_ (.Y(_0079_),
    .A(net164));
 sg13g2_inv_2 _0764_ (.Y(_0080_),
    .A(net95));
 sg13g2_inv_4 _0765_ (.A(net178),
    .Y(_0081_));
 sg13g2_inv_4 _0766_ (.A(net179),
    .Y(_0082_));
 sg13g2_inv_4 _0767_ (.A(net171),
    .Y(_0083_));
 sg13g2_inv_1 _0768_ (.Y(_0084_),
    .A(net205));
 sg13g2_inv_1 _0769_ (.Y(_0085_),
    .A(\raster.tscan.right_err[6] ));
 sg13g2_inv_1 _0770_ (.Y(_0086_),
    .A(net238));
 sg13g2_inv_1 _0771_ (.Y(_0087_),
    .A(net198));
 sg13g2_inv_1 _0772_ (.Y(_0088_),
    .A(net194));
 sg13g2_inv_1 _0773_ (.Y(_0089_),
    .A(net209));
 sg13g2_inv_1 _0774_ (.Y(_0090_),
    .A(\raster.tscan.right_x[4] ));
 sg13g2_inv_1 _0775_ (.Y(_0091_),
    .A(net183));
 sg13g2_inv_2 _0776_ (.Y(_0092_),
    .A(net186));
 sg13g2_inv_1 _0777_ (.Y(_0093_),
    .A(\raster.tscan.left_err[1] ));
 sg13g2_inv_2 _0778_ (.Y(_0094_),
    .A(net222));
 sg13g2_inv_1 _0779_ (.Y(_0095_),
    .A(\raster.tscan.left_err[4] ));
 sg13g2_inv_1 _0780_ (.Y(_0096_),
    .A(net197));
 sg13g2_inv_2 _0781_ (.Y(_0097_),
    .A(net202));
 sg13g2_inv_2 _0782_ (.Y(_0098_),
    .A(net229));
 sg13g2_inv_1 _0783_ (.Y(_0099_),
    .A(\raster.tscan.left_x[1] ));
 sg13g2_inv_1 _0784_ (.Y(_0100_),
    .A(net215));
 sg13g2_inv_2 _0785_ (.Y(_0101_),
    .A(net116));
 sg13g2_inv_1 _0786_ (.Y(_0102_),
    .A(net211));
 sg13g2_inv_1 _0787_ (.Y(_0103_),
    .A(net207));
 sg13g2_inv_1 _0788_ (.Y(_0104_),
    .A(net217));
 sg13g2_inv_1 _0789_ (.Y(_0105_),
    .A(\raster.tscan.right_x[9] ));
 sg13g2_inv_1 _0790_ (.Y(_0106_),
    .A(net90));
 sg13g2_nor3_1 _0791_ (.A(\raster.hpos[4] ),
    .B(\raster.hpos[5] ),
    .C(net167),
    .Y(_0107_));
 sg13g2_nand2_1 _0792_ (.Y(_0108_),
    .A(\raster.hpos[7] ),
    .B(\raster.hpos[9] ));
 sg13g2_nor2_1 _0793_ (.A(net166),
    .B(_0108_),
    .Y(_0109_));
 sg13g2_nor4_1 _0794_ (.A(\raster.hpos[1] ),
    .B(\raster.hpos[0] ),
    .C(\raster.hpos[3] ),
    .D(\raster.hpos[2] ),
    .Y(_0110_));
 sg13g2_and3_2 _0795_ (.X(_0111_),
    .A(_0107_),
    .B(_0109_),
    .C(_0110_));
 sg13g2_nand3_1 _0796_ (.B(_0109_),
    .C(_0110_),
    .A(_0107_),
    .Y(_0112_));
 sg13g2_nand2_1 _0797_ (.Y(_0113_),
    .A(net165),
    .B(net164));
 sg13g2_nand3_1 _0798_ (.B(net164),
    .C(\raster.hvsync_gen.vpos[2] ),
    .A(net165),
    .Y(_0114_));
 sg13g2_and4_1 _0799_ (.A(net165),
    .B(net164),
    .C(\raster.hvsync_gen.vpos[2] ),
    .D(\raster.hvsync_gen.vpos[3] ),
    .X(_0115_));
 sg13g2_nand2_1 _0800_ (.Y(_0116_),
    .A(net163),
    .B(_0115_));
 sg13g2_and2_1 _0801_ (.A(\raster.hvsync_gen.vpos[5] ),
    .B(\raster.hvsync_gen.vpos[6] ),
    .X(_0117_));
 sg13g2_nand3_1 _0802_ (.B(\raster.hvsync_gen.vpos[5] ),
    .C(_0115_),
    .A(net163),
    .Y(_0118_));
 sg13g2_nand3_1 _0803_ (.B(_0115_),
    .C(_0117_),
    .A(net163),
    .Y(_0119_));
 sg13g2_nand4_1 _0804_ (.B(\raster.hvsync_gen.vpos[7] ),
    .C(_0115_),
    .A(net163),
    .Y(_0120_),
    .D(_0117_));
 sg13g2_nor2b_1 _0805_ (.A(\raster.hvsync_gen.vpos[8] ),
    .B_N(_0120_),
    .Y(_0121_));
 sg13g2_nand3_1 _0806_ (.B(\raster.hvsync_gen.vpos[8] ),
    .C(_0117_),
    .A(\raster.hvsync_gen.vpos[7] ),
    .Y(_0122_));
 sg13g2_nor2_1 _0807_ (.A(_0116_),
    .B(_0122_),
    .Y(_0123_));
 sg13g2_xor2_1 _0808_ (.B(_0120_),
    .A(net104),
    .X(_0124_));
 sg13g2_o21ai_1 _0809_ (.B1(_0080_),
    .Y(_0125_),
    .A1(net147),
    .A2(_0121_));
 sg13g2_a21oi_2 _0810_ (.B1(_0125_),
    .Y(_0126_),
    .A2(_0124_),
    .A1(net147));
 sg13g2_xor2_1 _0811_ (.B(_0116_),
    .A(net193),
    .X(_0127_));
 sg13g2_xor2_1 _0812_ (.B(_0118_),
    .A(net182),
    .X(_0128_));
 sg13g2_nor3_1 _0813_ (.A(net151),
    .B(net149),
    .C(\raster.frame_counter[4] ),
    .Y(_0129_));
 sg13g2_or3_1 _0814_ (.A(net151),
    .B(net149),
    .C(\raster.frame_counter[4] ),
    .X(_0130_));
 sg13g2_nand2_2 _0815_ (.Y(_0131_),
    .A(net152),
    .B(_0130_));
 sg13g2_o21ai_1 _0816_ (.B1(_0127_),
    .Y(_0132_),
    .A1(_0128_),
    .A2(_0131_));
 sg13g2_xor2_1 _0817_ (.B(_0114_),
    .A(net188),
    .X(_0133_));
 sg13g2_xor2_1 _0818_ (.B(net150),
    .A(net151),
    .X(_0134_));
 sg13g2_nand2_1 _0819_ (.Y(_0135_),
    .A(net155),
    .B(_0134_));
 sg13g2_xnor2_1 _0820_ (.Y(_0136_),
    .A(_0133_),
    .B(_0135_));
 sg13g2_nand2b_1 _0821_ (.Y(_0137_),
    .B(_0113_),
    .A_N(\raster.hvsync_gen.vpos[2] ));
 sg13g2_xor2_1 _0822_ (.B(_0113_),
    .A(net99),
    .X(_0138_));
 sg13g2_nand2_2 _0823_ (.Y(_0139_),
    .A(net155),
    .B(net151));
 sg13g2_xnor2_1 _0824_ (.Y(_0140_),
    .A(_0138_),
    .B(_0139_));
 sg13g2_xnor2_1 _0825_ (.Y(_0141_),
    .A(net163),
    .B(_0115_));
 sg13g2_o21ai_1 _0826_ (.B1(\raster.frame_counter[4] ),
    .Y(_0142_),
    .A1(net151),
    .A2(net149));
 sg13g2_a21oi_2 _0827_ (.B1(net147),
    .Y(_0143_),
    .A2(_0142_),
    .A1(_0130_));
 sg13g2_nand2b_1 _0828_ (.Y(_0144_),
    .B(_0131_),
    .A_N(\raster.hvsync_gen.vpos[6] ));
 sg13g2_nand2b_1 _0829_ (.Y(_0145_),
    .B(_0144_),
    .A_N(_0127_));
 sg13g2_xor2_1 _0830_ (.B(_0119_),
    .A(net103),
    .X(_0146_));
 sg13g2_nor2_1 _0831_ (.A(net165),
    .B(net164),
    .Y(_0147_));
 sg13g2_xnor2_1 _0832_ (.Y(_0148_),
    .A(net165),
    .B(net164));
 sg13g2_nand2_2 _0833_ (.Y(_0149_),
    .A(net155),
    .B(\raster.frame_counter[1] ));
 sg13g2_xor2_1 _0834_ (.B(net165),
    .A(net156),
    .X(_0150_));
 sg13g2_xnor2_1 _0835_ (.Y(_0151_),
    .A(_0148_),
    .B(_0149_));
 sg13g2_nand2_1 _0836_ (.Y(_0152_),
    .A(_0150_),
    .B(_0151_));
 sg13g2_xnor2_1 _0837_ (.Y(_0153_),
    .A(_0141_),
    .B(_0143_));
 sg13g2_nor4_1 _0838_ (.A(_0136_),
    .B(_0140_),
    .C(_0152_),
    .D(_0153_),
    .Y(_0154_));
 sg13g2_and4_1 _0839_ (.A(_0132_),
    .B(_0145_),
    .C(_0146_),
    .D(_0154_),
    .X(_0155_));
 sg13g2_nand2_2 _0840_ (.Y(_0156_),
    .A(_0126_),
    .B(_0155_));
 sg13g2_and3_2 _0841_ (.X(_0157_),
    .A(net140),
    .B(_0126_),
    .C(_0155_));
 sg13g2_xnor2_1 _0842_ (.Y(_0158_),
    .A(net147),
    .B(_0146_));
 sg13g2_xnor2_1 _0843_ (.Y(_0159_),
    .A(net156),
    .B(_0146_));
 sg13g2_xnor2_1 _0844_ (.Y(_0160_),
    .A(net156),
    .B(_0128_));
 sg13g2_nand4_1 _0845_ (.B(\raster.hvsync_gen.vpos[5] ),
    .C(_0114_),
    .A(net156),
    .Y(_0161_),
    .D(_0137_));
 sg13g2_and2_1 _0846_ (.A(_0141_),
    .B(_0161_),
    .X(_0162_));
 sg13g2_nor2_1 _0847_ (.A(net156),
    .B(\raster.hvsync_gen.vpos[5] ),
    .Y(_0163_));
 sg13g2_a21o_1 _0848_ (.A2(_0163_),
    .A1(_0138_),
    .B1(_0141_),
    .X(_0164_));
 sg13g2_nand4_1 _0849_ (.B(net164),
    .C(_0133_),
    .A(net165),
    .Y(_0165_),
    .D(_0164_));
 sg13g2_nor4_1 _0850_ (.A(_0158_),
    .B(_0160_),
    .C(_0162_),
    .D(_0165_),
    .Y(_0166_));
 sg13g2_nand2_2 _0851_ (.Y(_0167_),
    .A(_0126_),
    .B(_0166_));
 sg13g2_nor2_1 _0852_ (.A(net135),
    .B(_0167_),
    .Y(_0168_));
 sg13g2_and4_1 _0853_ (.A(net178),
    .B(net140),
    .C(_0126_),
    .D(_0166_),
    .X(_0169_));
 sg13g2_a21o_2 _0854_ (.A2(_0157_),
    .A1(net171),
    .B1(_0169_),
    .X(_0170_));
 sg13g2_nor3_1 _0855_ (.A(\raster.hvsync_gen.vpos[3] ),
    .B(net163),
    .C(\raster.hvsync_gen.vpos[5] ),
    .Y(_0171_));
 sg13g2_nand4_1 _0856_ (.B(_0148_),
    .C(_0150_),
    .A(_0138_),
    .Y(_0172_),
    .D(_0171_));
 sg13g2_nor2b_1 _0857_ (.A(_0172_),
    .B_N(_0124_),
    .Y(_0173_));
 sg13g2_xnor2_1 _0858_ (.Y(_0174_),
    .A(net95),
    .B(_0123_));
 sg13g2_and4_1 _0859_ (.A(_0159_),
    .B(_0160_),
    .C(_0173_),
    .D(_0174_),
    .X(_0175_));
 sg13g2_nand2_1 _0860_ (.Y(_0176_),
    .A(net140),
    .B(_0175_));
 sg13g2_a21oi_1 _0861_ (.A1(_0106_),
    .A2(_0176_),
    .Y(_0010_),
    .B1(_0170_));
 sg13g2_nand2_1 _0862_ (.Y(_0177_),
    .A(net179),
    .B(_0167_));
 sg13g2_nand3_1 _0863_ (.B(_0157_),
    .C(_0167_),
    .A(net179),
    .Y(_0178_));
 sg13g2_nand2_1 _0864_ (.Y(_0179_),
    .A(net213),
    .B(net141));
 sg13g2_o21ai_1 _0865_ (.B1(_0178_),
    .Y(_0001_),
    .A1(_0081_),
    .A2(_0168_));
 sg13g2_nor2_1 _0866_ (.A(_0083_),
    .B(_0157_),
    .Y(_0180_));
 sg13g2_nor2_1 _0867_ (.A(_0167_),
    .B(_0179_),
    .Y(_0181_));
 sg13g2_nor2_2 _0868_ (.A(_0082_),
    .B(_0167_),
    .Y(_0182_));
 sg13g2_inv_2 _0869_ (.Y(_0183_),
    .A(_0182_));
 sg13g2_or2_1 _0870_ (.X(_0002_),
    .B(_0181_),
    .A(_0180_));
 sg13g2_or3_1 _0871_ (.A(_0082_),
    .B(_0157_),
    .C(_0168_),
    .X(_0184_));
 sg13g2_o21ai_1 _0872_ (.B1(_0184_),
    .Y(_0000_),
    .A1(net90),
    .A2(_0176_));
 sg13g2_and4_1 _0873_ (.A(\raster.hpos[4] ),
    .B(\raster.hpos[5] ),
    .C(\raster.hpos[7] ),
    .D(net167),
    .X(_0185_));
 sg13g2_nor4_1 _0874_ (.A(net87),
    .B(_0107_),
    .C(_0108_),
    .D(_0185_),
    .Y(_0003_));
 sg13g2_nand3b_1 _0875_ (.B(_0080_),
    .C(\raster.hvsync_gen.vpos[3] ),
    .Y(_0186_),
    .A_N(net163));
 sg13g2_nor4_1 _0876_ (.A(_0079_),
    .B(net99),
    .C(_0122_),
    .D(_0186_),
    .Y(_0004_));
 sg13g2_nand2b_1 _0877_ (.Y(_0187_),
    .B(\raster.tscan.left_x[6] ),
    .A_N(net167));
 sg13g2_a22oi_1 _0878_ (.Y(_0188_),
    .B1(\raster.tscan.left_x[1] ),
    .B2(_0071_),
    .A2(\raster.tscan.left_x[0] ),
    .A1(_0072_));
 sg13g2_a221oi_1 _0879_ (.B2(\raster.hpos[2] ),
    .C1(_0188_),
    .B1(_0101_),
    .A1(\raster.hpos[1] ),
    .Y(_0189_),
    .A2(_0099_));
 sg13g2_a221oi_1 _0880_ (.B2(_0074_),
    .C1(_0189_),
    .B1(\raster.tscan.left_x[2] ),
    .A1(_0073_),
    .Y(_0190_),
    .A2(\raster.tscan.left_x[3] ));
 sg13g2_a221oi_1 _0881_ (.B2(\raster.hpos[4] ),
    .C1(_0190_),
    .B1(_0102_),
    .A1(\raster.hpos[3] ),
    .Y(_0191_),
    .A2(_0100_));
 sg13g2_a221oi_1 _0882_ (.B2(_0076_),
    .C1(_0191_),
    .B1(\raster.tscan.left_x[5] ),
    .A1(_0075_),
    .Y(_0192_),
    .A2(\raster.tscan.left_x[4] ));
 sg13g2_nand2_1 _0883_ (.Y(_0193_),
    .A(\raster.hpos[6] ),
    .B(_0103_));
 sg13g2_o21ai_1 _0884_ (.B1(_0193_),
    .Y(_0194_),
    .A1(_0076_),
    .A2(\raster.tscan.left_x[5] ));
 sg13g2_o21ai_1 _0885_ (.B1(_0187_),
    .Y(_0195_),
    .A1(_0192_),
    .A2(_0194_));
 sg13g2_o21ai_1 _0886_ (.B1(_0195_),
    .Y(_0196_),
    .A1(_0077_),
    .A2(\raster.tscan.left_x[7] ));
 sg13g2_a22oi_1 _0887_ (.Y(_0197_),
    .B1(\raster.tscan.left_x[8] ),
    .B2(_0078_),
    .A2(\raster.tscan.left_x[7] ),
    .A1(_0077_));
 sg13g2_nor2b_1 _0888_ (.A(\raster.tscan.left_x[9] ),
    .B_N(\raster.hpos[9] ),
    .Y(_0198_));
 sg13g2_a221oi_1 _0889_ (.B2(_0197_),
    .C1(_0198_),
    .B1(_0196_),
    .A1(net166),
    .Y(_0199_),
    .A2(_0104_));
 sg13g2_nand2b_1 _0890_ (.Y(_0200_),
    .B(\raster.tscan.right_x[6] ),
    .A_N(net167));
 sg13g2_nand2b_1 _0891_ (.Y(_0201_),
    .B(\raster.tscan.right_x[1] ),
    .A_N(\raster.hpos[1] ));
 sg13g2_nand2b_1 _0892_ (.Y(_0202_),
    .B(\raster.tscan.right_x[0] ),
    .A_N(\raster.hpos[0] ));
 sg13g2_nor2b_1 _0893_ (.A(\raster.tscan.right_x[1] ),
    .B_N(\raster.hpos[1] ),
    .Y(_0203_));
 sg13g2_a221oi_1 _0894_ (.B2(_0202_),
    .C1(_0203_),
    .B1(_0201_),
    .A1(\raster.hpos[2] ),
    .Y(_0204_),
    .A2(_0088_));
 sg13g2_a221oi_1 _0895_ (.B2(_0073_),
    .C1(_0204_),
    .B1(\raster.tscan.right_x[3] ),
    .A1(_0074_),
    .Y(_0205_),
    .A2(\raster.tscan.right_x[2] ));
 sg13g2_a221oi_1 _0896_ (.B2(\raster.hpos[4] ),
    .C1(_0205_),
    .B1(_0090_),
    .A1(\raster.hpos[3] ),
    .Y(_0206_),
    .A2(_0089_));
 sg13g2_a221oi_1 _0897_ (.B2(_0076_),
    .C1(_0206_),
    .B1(\raster.tscan.right_x[5] ),
    .A1(_0075_),
    .Y(_0207_),
    .A2(\raster.tscan.right_x[4] ));
 sg13g2_nand2b_1 _0898_ (.Y(_0208_),
    .B(net167),
    .A_N(\raster.tscan.right_x[6] ));
 sg13g2_o21ai_1 _0899_ (.B1(_0208_),
    .Y(_0209_),
    .A1(_0076_),
    .A2(\raster.tscan.right_x[5] ));
 sg13g2_o21ai_1 _0900_ (.B1(_0200_),
    .Y(_0210_),
    .A1(_0207_),
    .A2(_0209_));
 sg13g2_o21ai_1 _0901_ (.B1(_0210_),
    .Y(_0211_),
    .A1(_0077_),
    .A2(\raster.tscan.right_x[7] ));
 sg13g2_a22oi_1 _0902_ (.Y(_0212_),
    .B1(\raster.tscan.right_x[8] ),
    .B2(_0078_),
    .A2(\raster.tscan.right_x[7] ),
    .A1(_0077_));
 sg13g2_a22oi_1 _0903_ (.Y(_0213_),
    .B1(_0211_),
    .B2(_0212_),
    .A2(_0092_),
    .A1(net166));
 sg13g2_xor2_1 _0904_ (.B(\raster.tscan.right_x[9] ),
    .A(\raster.hpos[9] ),
    .X(_0214_));
 sg13g2_nor2_1 _0905_ (.A(_0213_),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nand2b_1 _0906_ (.Y(_0216_),
    .B(\raster.tscan.left_x[9] ),
    .A_N(\raster.hpos[9] ));
 sg13g2_o21ai_1 _0907_ (.B1(\raster.hpos[9] ),
    .Y(_0217_),
    .A1(net166),
    .A2(_0105_));
 sg13g2_nor2_1 _0908_ (.A(net177),
    .B(net171),
    .Y(_0218_));
 sg13g2_nor2_2 _0909_ (.A(net177),
    .B(net179),
    .Y(_0219_));
 sg13g2_or2_1 _0910_ (.X(_0220_),
    .B(net179),
    .A(net177));
 sg13g2_nor2_1 _0911_ (.A(net171),
    .B(net161),
    .Y(_0221_));
 sg13g2_nand2_2 _0912_ (.Y(_0222_),
    .A(_0083_),
    .B(net162));
 sg13g2_nand2_1 _0913_ (.Y(_0223_),
    .A(_0080_),
    .B(_0108_));
 sg13g2_nand4_1 _0914_ (.B(_0216_),
    .C(_0217_),
    .A(_0122_),
    .Y(_0224_),
    .D(_0222_));
 sg13g2_nor4_2 _0915_ (.A(_0199_),
    .B(_0215_),
    .C(_0223_),
    .Y(uo_out[4]),
    .D(_0224_));
 sg13g2_xnor2_1 _0916_ (.Y(_0225_),
    .A(\raster.hpos[0] ),
    .B(net165));
 sg13g2_and3_2 _0917_ (.X(uo_out[5]),
    .A(net147),
    .B(uo_out[4]),
    .C(_0225_));
 sg13g2_xor2_1 _0918_ (.B(\raster.frame_counter[1] ),
    .A(net155),
    .X(_0005_));
 sg13g2_nand3_1 _0919_ (.B(\raster.frame_counter[1] ),
    .C(net151),
    .A(net152),
    .Y(_0226_));
 sg13g2_xnor2_1 _0920_ (.Y(_0006_),
    .A(\raster.frame_counter[2] ),
    .B(_0149_));
 sg13g2_nand4_1 _0921_ (.B(\raster.frame_counter[1] ),
    .C(net151),
    .A(net155),
    .Y(_0227_),
    .D(net149));
 sg13g2_xnor2_1 _0922_ (.Y(_0007_),
    .A(net149),
    .B(_0226_));
 sg13g2_xnor2_1 _0923_ (.Y(_0008_),
    .A(\raster.frame_counter[4] ),
    .B(_0227_));
 sg13g2_nor2_2 _0924_ (.A(net213),
    .B(net137),
    .Y(_0228_));
 sg13g2_nand2_1 _0925_ (.Y(_0229_),
    .A(_0009_),
    .B(_0228_));
 sg13g2_nand2_1 _0926_ (.Y(_0230_),
    .A(net180),
    .B(_0229_));
 sg13g2_nor3_2 _0927_ (.A(_0009_),
    .B(net138),
    .C(_0175_),
    .Y(_0231_));
 sg13g2_a21oi_1 _0928_ (.A1(\raster.tscan.left_err[9] ),
    .A2(net146),
    .Y(_0232_),
    .B1(net142));
 sg13g2_or2_1 _0929_ (.X(_0233_),
    .B(_0232_),
    .A(_0231_));
 sg13g2_nor2_1 _0930_ (.A(_0084_),
    .B(net142),
    .Y(_0234_));
 sg13g2_or2_1 _0931_ (.X(_0235_),
    .B(_0233_),
    .A(_0230_));
 sg13g2_nor2_2 _0932_ (.A(net135),
    .B(_0177_),
    .Y(_0236_));
 sg13g2_or2_1 _0933_ (.X(_0237_),
    .B(_0236_),
    .A(_0235_));
 sg13g2_nor2_2 _0934_ (.A(net141),
    .B(_0235_),
    .Y(_0238_));
 sg13g2_mux2_1 _0935_ (.A0(net128),
    .A1(_0238_),
    .S(_0098_),
    .X(_0011_));
 sg13g2_nor2_1 _0936_ (.A(net160),
    .B(net162),
    .Y(_0239_));
 sg13g2_nor3_1 _0937_ (.A(net160),
    .B(_0101_),
    .C(net162),
    .Y(_0240_));
 sg13g2_o21ai_1 _0938_ (.B1(_0101_),
    .Y(_0241_),
    .A1(net160),
    .A2(net162));
 sg13g2_nor2b_1 _0939_ (.A(_0240_),
    .B_N(_0241_),
    .Y(_0242_));
 sg13g2_nand3_1 _0940_ (.B(\raster.tscan.left_x[1] ),
    .C(net161),
    .A(net148),
    .Y(_0243_));
 sg13g2_a21oi_1 _0941_ (.A1(net148),
    .A2(_0220_),
    .Y(_0244_),
    .B1(\raster.tscan.left_x[1] ));
 sg13g2_xor2_1 _0942_ (.B(net144),
    .A(net121),
    .X(_0245_));
 sg13g2_o21ai_1 _0943_ (.B1(_0243_),
    .Y(_0246_),
    .A1(_0098_),
    .A2(_0244_));
 sg13g2_xnor2_1 _0944_ (.Y(_0247_),
    .A(_0242_),
    .B(_0246_));
 sg13g2_a22oi_1 _0945_ (.Y(_0012_),
    .B1(_0238_),
    .B2(_0247_),
    .A2(net128),
    .A1(_0101_));
 sg13g2_nand2_1 _0946_ (.Y(_0248_),
    .A(net106),
    .B(net128));
 sg13g2_nand2_1 _0947_ (.Y(_0249_),
    .A(\raster.tscan.left_x[8] ),
    .B(net143));
 sg13g2_xnor2_1 _0948_ (.Y(_0250_),
    .A(net217),
    .B(net143));
 sg13g2_xnor2_1 _0949_ (.Y(_0251_),
    .A(\raster.tscan.left_x[5] ),
    .B(net143));
 sg13g2_xnor2_1 _0950_ (.Y(_0252_),
    .A(net211),
    .B(net144));
 sg13g2_nor2_1 _0951_ (.A(\raster.tscan.left_x[3] ),
    .B(net144),
    .Y(_0253_));
 sg13g2_a21oi_1 _0952_ (.A1(_0241_),
    .A2(_0246_),
    .Y(_0254_),
    .B1(_0240_));
 sg13g2_a221oi_1 _0953_ (.B2(_0246_),
    .C1(_0240_),
    .B1(_0242_),
    .A1(\raster.tscan.left_x[3] ),
    .Y(_0255_),
    .A2(net144));
 sg13g2_nor3_1 _0954_ (.A(_0252_),
    .B(_0253_),
    .C(_0255_),
    .Y(_0256_));
 sg13g2_nor2b_2 _0955_ (.A(_0251_),
    .B_N(_0256_),
    .Y(_0257_));
 sg13g2_xor2_1 _0956_ (.B(net143),
    .A(net189),
    .X(_0258_));
 sg13g2_nand2_1 _0957_ (.Y(_0259_),
    .A(\raster.tscan.left_x[6] ),
    .B(net143));
 sg13g2_xnor2_1 _0958_ (.Y(_0260_),
    .A(_0103_),
    .B(net143));
 sg13g2_nand3_1 _0959_ (.B(_0258_),
    .C(_0260_),
    .A(_0257_),
    .Y(_0261_));
 sg13g2_o21ai_1 _0960_ (.B1(net143),
    .Y(_0262_),
    .A1(\raster.tscan.left_x[4] ),
    .A2(\raster.tscan.left_x[5] ));
 sg13g2_inv_1 _0961_ (.Y(_0263_),
    .A(_0262_));
 sg13g2_o21ai_1 _0962_ (.B1(net143),
    .Y(_0264_),
    .A1(\raster.tscan.left_x[6] ),
    .A2(\raster.tscan.left_x[7] ));
 sg13g2_and2_1 _0963_ (.A(_0262_),
    .B(_0264_),
    .X(_0265_));
 sg13g2_a21o_1 _0964_ (.A2(_0265_),
    .A1(_0261_),
    .B1(_0250_),
    .X(_0266_));
 sg13g2_xnor2_1 _0965_ (.Y(_0267_),
    .A(net106),
    .B(net144));
 sg13g2_nand3_1 _0966_ (.B(_0266_),
    .C(_0267_),
    .A(_0249_),
    .Y(_0268_));
 sg13g2_a21oi_1 _0967_ (.A1(_0249_),
    .A2(_0266_),
    .Y(_0269_),
    .B1(_0267_));
 sg13g2_nand2_1 _0968_ (.Y(_0270_),
    .A(_0238_),
    .B(_0268_));
 sg13g2_o21ai_1 _0969_ (.B1(_0248_),
    .Y(_0013_),
    .A1(_0269_),
    .A2(_0270_));
 sg13g2_nand3_1 _0970_ (.B(_0218_),
    .C(_0228_),
    .A(_0009_),
    .Y(_0271_));
 sg13g2_nand2_1 _0971_ (.Y(_0272_),
    .A(net180),
    .B(_0271_));
 sg13g2_nor3_1 _0972_ (.A(_0170_),
    .B(_0231_),
    .C(_0272_),
    .Y(_0273_));
 sg13g2_a21o_1 _0973_ (.A2(net146),
    .A1(\raster.tscan.right_err[9] ),
    .B1(net140),
    .X(_0274_));
 sg13g2_nor4_1 _0974_ (.A(_0170_),
    .B(_0181_),
    .C(_0231_),
    .D(_0272_),
    .Y(_0275_));
 sg13g2_and2_1 _0975_ (.A(_0274_),
    .B(_0275_),
    .X(_0276_));
 sg13g2_nor2_1 _0976_ (.A(_0149_),
    .B(net146),
    .Y(_0277_));
 sg13g2_nor2b_1 _0977_ (.A(_0218_),
    .B_N(\raster.tscan.right_err[0] ),
    .Y(_0278_));
 sg13g2_nor3_1 _0978_ (.A(net134),
    .B(_0277_),
    .C(_0278_),
    .Y(_0279_));
 sg13g2_nand2_1 _0979_ (.Y(_0280_),
    .A(_0156_),
    .B(_0279_));
 sg13g2_a21oi_1 _0980_ (.A1(net125),
    .A2(_0280_),
    .Y(_0281_),
    .B1(net97));
 sg13g2_nand2_1 _0981_ (.Y(_0282_),
    .A(net157),
    .B(net174));
 sg13g2_nor2_1 _0982_ (.A(net97),
    .B(_0282_),
    .Y(_0283_));
 sg13g2_a21oi_1 _0983_ (.A1(net97),
    .A2(_0282_),
    .Y(_0284_),
    .B1(net140));
 sg13g2_nand2b_1 _0984_ (.Y(_0285_),
    .B(_0284_),
    .A_N(_0283_));
 sg13g2_a21oi_1 _0985_ (.A1(_0126_),
    .A2(_0155_),
    .Y(_0286_),
    .B1(_0082_));
 sg13g2_o21ai_1 _0986_ (.B1(_0279_),
    .Y(_0287_),
    .A1(net164),
    .A2(_0082_));
 sg13g2_o21ai_1 _0987_ (.B1(_0285_),
    .Y(_0288_),
    .A1(_0286_),
    .A2(_0287_));
 sg13g2_a21oi_1 _0988_ (.A1(net125),
    .A2(_0288_),
    .Y(_0014_),
    .B1(net98));
 sg13g2_nand2_1 _0989_ (.Y(_0289_),
    .A(net139),
    .B(net145));
 sg13g2_nand2_1 _0990_ (.Y(_0290_),
    .A(\raster.tscan.right_err[1] ),
    .B(_0149_));
 sg13g2_xnor2_1 _0991_ (.Y(_0291_),
    .A(\raster.tscan.right_err[1] ),
    .B(_0149_));
 sg13g2_xor2_1 _0992_ (.B(_0291_),
    .A(_0283_),
    .X(_0292_));
 sg13g2_nor2_1 _0993_ (.A(net174),
    .B(\raster.tscan.right_err[1] ),
    .Y(_0293_));
 sg13g2_a21oi_1 _0994_ (.A1(_0083_),
    .A2(\raster.tscan.right_err[1] ),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_nor2_2 _0995_ (.A(_0082_),
    .B(_0156_),
    .Y(_0295_));
 sg13g2_nor2_1 _0996_ (.A(net218),
    .B(net124),
    .Y(_0296_));
 sg13g2_a21oi_1 _0997_ (.A1(net218),
    .A2(_0286_),
    .Y(_0297_),
    .B1(_0221_));
 sg13g2_a21oi_1 _0998_ (.A1(_0139_),
    .A2(_0295_),
    .Y(_0298_),
    .B1(_0294_));
 sg13g2_o21ai_1 _0999_ (.B1(net139),
    .Y(_0299_),
    .A1(_0139_),
    .A2(net145));
 sg13g2_a21oi_1 _1000_ (.A1(_0297_),
    .A2(_0298_),
    .Y(_0300_),
    .B1(_0299_));
 sg13g2_a21oi_1 _1001_ (.A1(net134),
    .A2(_0292_),
    .Y(_0301_),
    .B1(_0300_));
 sg13g2_a21oi_1 _1002_ (.A1(net124),
    .A2(_0301_),
    .Y(_0015_),
    .B1(_0296_));
 sg13g2_o21ai_1 _1003_ (.B1(_0290_),
    .Y(_0302_),
    .A1(_0283_),
    .A2(_0291_));
 sg13g2_nand2b_2 _1004_ (.Y(_0303_),
    .B(net153),
    .A_N(net151));
 sg13g2_nor2_1 _1005_ (.A(net174),
    .B(\raster.frame_counter[1] ),
    .Y(_0304_));
 sg13g2_nand2_1 _1006_ (.Y(_0305_),
    .A(net155),
    .B(_0081_));
 sg13g2_mux2_1 _1007_ (.A0(_0303_),
    .A1(_0139_),
    .S(_0304_),
    .X(_0306_));
 sg13g2_nor2b_1 _1008_ (.A(_0306_),
    .B_N(\raster.tscan.right_err[2] ),
    .Y(_0307_));
 sg13g2_xnor2_1 _1009_ (.Y(_0308_),
    .A(net170),
    .B(_0306_));
 sg13g2_o21ai_1 _1010_ (.B1(net133),
    .Y(_0309_),
    .A1(_0302_),
    .A2(_0308_));
 sg13g2_a21oi_1 _1011_ (.A1(_0302_),
    .A2(_0308_),
    .Y(_0310_),
    .B1(_0309_));
 sg13g2_or2_1 _1012_ (.X(_0311_),
    .B(_0286_),
    .A(net171));
 sg13g2_nand2b_1 _1013_ (.Y(_0312_),
    .B(_0311_),
    .A_N(net170));
 sg13g2_and2_1 _1014_ (.A(net154),
    .B(net150),
    .X(_0313_));
 sg13g2_nand2_1 _1015_ (.Y(_0314_),
    .A(net154),
    .B(net150));
 sg13g2_nor2_1 _1016_ (.A(\raster.tscan.right_err[1] ),
    .B(net170),
    .Y(_0315_));
 sg13g2_xnor2_1 _1017_ (.Y(_0316_),
    .A(\raster.tscan.right_err[1] ),
    .B(net170));
 sg13g2_a221oi_1 _1018_ (.B2(net174),
    .C1(_0221_),
    .B1(_0316_),
    .A1(_0295_),
    .Y(_0317_),
    .A2(_0313_));
 sg13g2_o21ai_1 _1019_ (.B1(net139),
    .Y(_0318_),
    .A1(net154),
    .A2(net145));
 sg13g2_a221oi_1 _1020_ (.B2(_0317_),
    .C1(_0318_),
    .B1(_0312_),
    .A1(_0134_),
    .Y(_0319_),
    .A2(_0289_));
 sg13g2_nor2_1 _1021_ (.A(_0310_),
    .B(_0319_),
    .Y(_0320_));
 sg13g2_nor2_1 _1022_ (.A(net170),
    .B(net124),
    .Y(_0321_));
 sg13g2_a21oi_1 _1023_ (.A1(net125),
    .A2(_0320_),
    .Y(_0016_),
    .B1(_0321_));
 sg13g2_nand3_1 _1024_ (.B(net174),
    .C(net150),
    .A(net155),
    .Y(_0322_));
 sg13g2_o21ai_1 _1025_ (.B1(_0322_),
    .Y(_0323_),
    .A1(_0007_),
    .A2(_0305_));
 sg13g2_nand2_1 _1026_ (.Y(_0324_),
    .A(net169),
    .B(_0323_));
 sg13g2_nor2_1 _1027_ (.A(net169),
    .B(_0323_),
    .Y(_0325_));
 sg13g2_xnor2_1 _1028_ (.Y(_0326_),
    .A(\raster.tscan.right_err[3] ),
    .B(_0323_));
 sg13g2_a21oi_1 _1029_ (.A1(_0302_),
    .A2(_0308_),
    .Y(_0327_),
    .B1(_0307_));
 sg13g2_xnor2_1 _1030_ (.Y(_0328_),
    .A(_0326_),
    .B(_0327_));
 sg13g2_xnor2_1 _1031_ (.Y(_0329_),
    .A(net170),
    .B(net169));
 sg13g2_o21ai_1 _1032_ (.B1(net153),
    .Y(_0330_),
    .A1(net149),
    .A2(\raster.frame_counter[4] ));
 sg13g2_a21oi_1 _1033_ (.A1(net149),
    .A2(\raster.frame_counter[4] ),
    .Y(_0331_),
    .B1(_0330_));
 sg13g2_a21o_2 _1034_ (.A2(\raster.frame_counter[4] ),
    .A1(net149),
    .B1(_0330_),
    .X(_0332_));
 sg13g2_nand2_1 _1035_ (.Y(_0333_),
    .A(net152),
    .B(net169));
 sg13g2_xnor2_1 _1036_ (.Y(_0334_),
    .A(net153),
    .B(net169));
 sg13g2_o21ai_1 _1037_ (.B1(net173),
    .Y(_0335_),
    .A1(_0315_),
    .A2(_0334_));
 sg13g2_a21oi_1 _1038_ (.A1(_0315_),
    .A2(_0334_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_a21oi_1 _1039_ (.A1(_0143_),
    .A2(_0221_),
    .Y(_0337_),
    .B1(net134));
 sg13g2_a221oi_1 _1040_ (.B2(_0295_),
    .C1(_0336_),
    .B1(_0331_),
    .A1(_0311_),
    .Y(_0338_),
    .A2(_0329_));
 sg13g2_a22oi_1 _1041_ (.Y(_0339_),
    .B1(_0337_),
    .B2(_0338_),
    .A2(_0328_),
    .A1(net133));
 sg13g2_mux2_1 _1042_ (.A0(net169),
    .A1(_0339_),
    .S(net124),
    .X(_0017_));
 sg13g2_or3_1 _1043_ (.A(\raster.frame_counter[1] ),
    .B(net150),
    .C(_0139_),
    .X(_0340_));
 sg13g2_or2_1 _1044_ (.X(_0341_),
    .B(_0340_),
    .A(_0143_));
 sg13g2_a21oi_1 _1045_ (.A1(_0143_),
    .A2(_0340_),
    .Y(_0342_),
    .B1(net173));
 sg13g2_a22oi_1 _1046_ (.Y(_0343_),
    .B1(_0341_),
    .B2(_0342_),
    .A2(_0332_),
    .A1(net173));
 sg13g2_and2_1 _1047_ (.A(\raster.tscan.right_err[4] ),
    .B(_0343_),
    .X(_0344_));
 sg13g2_or2_1 _1048_ (.X(_0345_),
    .B(_0343_),
    .A(\raster.tscan.right_err[4] ));
 sg13g2_nand2b_1 _1049_ (.Y(_0346_),
    .B(_0345_),
    .A_N(_0344_));
 sg13g2_o21ai_1 _1050_ (.B1(_0324_),
    .Y(_0347_),
    .A1(_0325_),
    .A2(_0327_));
 sg13g2_xnor2_1 _1051_ (.Y(_0348_),
    .A(_0346_),
    .B(_0347_));
 sg13g2_nor3_1 _1052_ (.A(net170),
    .B(net169),
    .C(\raster.tscan.right_err[4] ),
    .Y(_0349_));
 sg13g2_o21ai_1 _1053_ (.B1(\raster.tscan.right_err[4] ),
    .Y(_0350_),
    .A1(net170),
    .A2(net169));
 sg13g2_nand2b_1 _1054_ (.Y(_0351_),
    .B(_0350_),
    .A_N(_0349_));
 sg13g2_o21ai_1 _1055_ (.B1(_0333_),
    .Y(_0352_),
    .A1(_0315_),
    .A2(_0334_));
 sg13g2_and2_1 _1056_ (.A(\raster.tscan.right_err[4] ),
    .B(_0352_),
    .X(_0353_));
 sg13g2_o21ai_1 _1057_ (.B1(net173),
    .Y(_0354_),
    .A1(\raster.tscan.right_err[4] ),
    .A2(_0352_));
 sg13g2_o21ai_1 _1058_ (.B1(net145),
    .Y(_0355_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_a221oi_1 _1059_ (.B2(_0311_),
    .C1(_0355_),
    .B1(_0351_),
    .A1(_0295_),
    .Y(_0356_),
    .A2(_0330_));
 sg13g2_o21ai_1 _1060_ (.B1(net139),
    .Y(_0357_),
    .A1(_0131_),
    .A2(net145));
 sg13g2_nor2_1 _1061_ (.A(_0356_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_a21o_1 _1062_ (.A2(_0348_),
    .A1(net133),
    .B1(_0358_),
    .X(_0359_));
 sg13g2_mux2_1 _1063_ (.A0(net216),
    .A1(_0359_),
    .S(net124),
    .X(_0018_));
 sg13g2_a21oi_1 _1064_ (.A1(_0345_),
    .A2(_0347_),
    .Y(_0360_),
    .B1(_0344_));
 sg13g2_o21ai_1 _1065_ (.B1(_0330_),
    .Y(_0361_),
    .A1(net173),
    .A2(_0226_));
 sg13g2_inv_1 _1066_ (.Y(_0362_),
    .A(_0361_));
 sg13g2_nand2_1 _1067_ (.Y(_0363_),
    .A(\raster.tscan.right_err[5] ),
    .B(_0362_));
 sg13g2_xor2_1 _1068_ (.B(_0361_),
    .A(\raster.tscan.right_err[5] ),
    .X(_0364_));
 sg13g2_xor2_1 _1069_ (.B(_0364_),
    .A(_0360_),
    .X(_0365_));
 sg13g2_nor2b_1 _1070_ (.A(_0349_),
    .B_N(\raster.tscan.right_err[5] ),
    .Y(_0366_));
 sg13g2_xnor2_1 _1071_ (.Y(_0367_),
    .A(\raster.tscan.right_err[5] ),
    .B(_0349_));
 sg13g2_nor2_1 _1072_ (.A(\raster.tscan.right_err[5] ),
    .B(_0353_),
    .Y(_0368_));
 sg13g2_nand3_1 _1073_ (.B(\raster.tscan.right_err[5] ),
    .C(_0352_),
    .A(\raster.tscan.right_err[4] ),
    .Y(_0369_));
 sg13g2_nand2_1 _1074_ (.Y(_0370_),
    .A(net173),
    .B(_0369_));
 sg13g2_o21ai_1 _1075_ (.B1(net145),
    .Y(_0371_),
    .A1(_0368_),
    .A2(_0370_));
 sg13g2_a221oi_1 _1076_ (.B2(_0367_),
    .C1(_0371_),
    .B1(_0311_),
    .A1(net147),
    .Y(_0372_),
    .A2(_0295_));
 sg13g2_nor3_1 _1077_ (.A(net147),
    .B(_0130_),
    .C(net145),
    .Y(_0373_));
 sg13g2_nor3_1 _1078_ (.A(net133),
    .B(_0372_),
    .C(_0373_),
    .Y(_0374_));
 sg13g2_a21oi_1 _1079_ (.A1(net133),
    .A2(_0365_),
    .Y(_0375_),
    .B1(_0374_));
 sg13g2_nor2_1 _1080_ (.A(net204),
    .B(net124),
    .Y(_0376_));
 sg13g2_a21oi_1 _1081_ (.A1(net124),
    .A2(_0375_),
    .Y(_0019_),
    .B1(_0376_));
 sg13g2_o21ai_1 _1082_ (.B1(_0363_),
    .Y(_0377_),
    .A1(_0360_),
    .A2(_0364_));
 sg13g2_o21ai_1 _1083_ (.B1(net153),
    .Y(_0378_),
    .A1(net173),
    .A2(_0129_));
 sg13g2_o21ai_1 _1084_ (.B1(_0378_),
    .Y(_0379_),
    .A1(net173),
    .A2(_0341_));
 sg13g2_nor2_1 _1085_ (.A(_0085_),
    .B(_0379_),
    .Y(_0380_));
 sg13g2_nand2_1 _1086_ (.Y(_0381_),
    .A(_0085_),
    .B(_0379_));
 sg13g2_nor2b_1 _1087_ (.A(_0380_),
    .B_N(_0381_),
    .Y(_0382_));
 sg13g2_xnor2_1 _1088_ (.Y(_0383_),
    .A(_0377_),
    .B(_0382_));
 sg13g2_xor2_1 _1089_ (.B(\raster.tscan.right_err[6] ),
    .A(net152),
    .X(_0384_));
 sg13g2_nor2_2 _1090_ (.A(_0081_),
    .B(net133),
    .Y(_0385_));
 sg13g2_nor2b_1 _1091_ (.A(_0369_),
    .B_N(_0384_),
    .Y(_0386_));
 sg13g2_and2_1 _1092_ (.A(\raster.tscan.right_err[6] ),
    .B(_0366_),
    .X(_0387_));
 sg13g2_xnor2_1 _1093_ (.Y(_0388_),
    .A(_0085_),
    .B(_0366_));
 sg13g2_and2_1 _1094_ (.A(_0311_),
    .B(_0388_),
    .X(_0389_));
 sg13g2_xnor2_1 _1095_ (.Y(_0390_),
    .A(_0369_),
    .B(_0384_));
 sg13g2_a22oi_1 _1096_ (.Y(_0391_),
    .B1(_0390_),
    .B2(_0385_),
    .A2(_0389_),
    .A1(net139));
 sg13g2_o21ai_1 _1097_ (.B1(_0391_),
    .Y(_0392_),
    .A1(net139),
    .A2(_0383_));
 sg13g2_mux2_1 _1098_ (.A0(net196),
    .A1(_0392_),
    .S(net124),
    .X(_0020_));
 sg13g2_a21oi_1 _1099_ (.A1(_0377_),
    .A2(_0381_),
    .Y(_0393_),
    .B1(_0380_));
 sg13g2_o21ai_1 _1100_ (.B1(net133),
    .Y(_0394_),
    .A1(_0086_),
    .A2(_0393_));
 sg13g2_nand2_1 _1101_ (.Y(_0395_),
    .A(net125),
    .B(_0394_));
 sg13g2_a21oi_1 _1102_ (.A1(net125),
    .A2(_0394_),
    .Y(_0396_),
    .B1(_0086_));
 sg13g2_nor3_1 _1103_ (.A(net238),
    .B(net139),
    .C(_0393_),
    .Y(_0397_));
 sg13g2_xnor2_1 _1104_ (.Y(_0398_),
    .A(\raster.tscan.right_err[7] ),
    .B(_0387_));
 sg13g2_nand2_1 _1105_ (.Y(_0399_),
    .A(_0311_),
    .B(_0398_));
 sg13g2_a21oi_1 _1106_ (.A1(net152),
    .A2(\raster.tscan.right_err[6] ),
    .Y(_0400_),
    .B1(_0386_));
 sg13g2_nand2_1 _1107_ (.Y(_0401_),
    .A(net152),
    .B(\raster.tscan.right_err[7] ));
 sg13g2_nor2_1 _1108_ (.A(net152),
    .B(\raster.tscan.right_err[7] ),
    .Y(_0402_));
 sg13g2_xnor2_1 _1109_ (.Y(_0403_),
    .A(net152),
    .B(\raster.tscan.right_err[7] ));
 sg13g2_a21oi_1 _1110_ (.A1(_0400_),
    .A2(_0403_),
    .Y(_0404_),
    .B1(_0081_));
 sg13g2_o21ai_1 _1111_ (.B1(_0404_),
    .Y(_0405_),
    .A1(_0400_),
    .A2(_0403_));
 sg13g2_a21oi_1 _1112_ (.A1(_0399_),
    .A2(_0405_),
    .Y(_0406_),
    .B1(net133));
 sg13g2_o21ai_1 _1113_ (.B1(net125),
    .Y(_0407_),
    .A1(_0397_),
    .A2(_0406_));
 sg13g2_nand2b_1 _1114_ (.Y(_0021_),
    .B(_0407_),
    .A_N(_0396_));
 sg13g2_nor3_1 _1115_ (.A(_0086_),
    .B(_0087_),
    .C(_0393_),
    .Y(_0408_));
 sg13g2_or2_1 _1116_ (.X(_0409_),
    .B(_0408_),
    .A(net139));
 sg13g2_a21oi_1 _1117_ (.A1(_0400_),
    .A2(_0401_),
    .Y(_0410_),
    .B1(_0402_));
 sg13g2_nor2_1 _1118_ (.A(\raster.tscan.right_err[8] ),
    .B(_0410_),
    .Y(_0411_));
 sg13g2_xnor2_1 _1119_ (.Y(_0412_),
    .A(net198),
    .B(_0410_));
 sg13g2_or3_1 _1120_ (.A(\raster.tscan.right_err[7] ),
    .B(\raster.tscan.right_err[8] ),
    .C(_0387_),
    .X(_0413_));
 sg13g2_o21ai_1 _1121_ (.B1(\raster.tscan.right_err[8] ),
    .Y(_0414_),
    .A1(\raster.tscan.right_err[7] ),
    .A2(_0387_));
 sg13g2_a21oi_1 _1122_ (.A1(_0413_),
    .A2(_0414_),
    .Y(_0415_),
    .B1(net134));
 sg13g2_a22oi_1 _1123_ (.Y(_0416_),
    .B1(_0415_),
    .B2(_0311_),
    .A2(_0412_),
    .A1(_0385_));
 sg13g2_and2_1 _1124_ (.A(net125),
    .B(_0416_),
    .X(_0417_));
 sg13g2_a22oi_1 _1125_ (.Y(_0022_),
    .B1(_0409_),
    .B2(_0417_),
    .A2(_0395_),
    .A1(_0087_));
 sg13g2_nand2b_1 _1126_ (.Y(_0418_),
    .B(_0178_),
    .A_N(_0233_));
 sg13g2_a21oi_2 _1127_ (.B1(net177),
    .Y(_0419_),
    .A2(_0167_),
    .A1(net179));
 sg13g2_nor4_1 _1128_ (.A(_0236_),
    .B(_0272_),
    .C(_0385_),
    .D(_0418_),
    .Y(_0420_));
 sg13g2_and2_1 _1129_ (.A(net159),
    .B(\raster.tscan.left_err[0] ),
    .X(_0421_));
 sg13g2_xor2_1 _1130_ (.B(net109),
    .A(net158),
    .X(_0422_));
 sg13g2_nor2_2 _1131_ (.A(net157),
    .B(net137),
    .Y(_0423_));
 sg13g2_o21ai_1 _1132_ (.B1(net142),
    .Y(_0424_),
    .A1(net148),
    .A2(net146));
 sg13g2_a21oi_1 _1133_ (.A1(net171),
    .A2(net109),
    .Y(_0425_),
    .B1(_0424_));
 sg13g2_o21ai_1 _1134_ (.B1(_0425_),
    .Y(_0426_),
    .A1(_0149_),
    .A2(_0183_));
 sg13g2_o21ai_1 _1135_ (.B1(_0426_),
    .Y(_0427_),
    .A1(net142),
    .A2(_0422_));
 sg13g2_nor2_1 _1136_ (.A(net109),
    .B(_0420_),
    .Y(_0428_));
 sg13g2_a21oi_1 _1137_ (.A1(_0420_),
    .A2(_0427_),
    .Y(_0023_),
    .B1(net110));
 sg13g2_nand2_1 _1138_ (.Y(_0429_),
    .A(net121),
    .B(net128));
 sg13g2_or2_1 _1139_ (.X(_0430_),
    .B(net128),
    .A(_0228_));
 sg13g2_xnor2_1 _1140_ (.Y(_0431_),
    .A(_0098_),
    .B(_0245_));
 sg13g2_nor2_1 _1141_ (.A(net141),
    .B(_0431_),
    .Y(_0432_));
 sg13g2_o21ai_1 _1142_ (.B1(_0429_),
    .Y(_0024_),
    .A1(_0430_),
    .A2(_0432_));
 sg13g2_a21oi_1 _1143_ (.A1(net148),
    .A2(_0228_),
    .Y(_0433_),
    .B1(net129));
 sg13g2_xnor2_1 _1144_ (.Y(_0434_),
    .A(net215),
    .B(net144));
 sg13g2_a21oi_1 _1145_ (.A1(_0254_),
    .A2(_0434_),
    .Y(_0435_),
    .B1(net141));
 sg13g2_o21ai_1 _1146_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0254_),
    .A2(_0434_));
 sg13g2_a22oi_1 _1147_ (.Y(_0025_),
    .B1(_0433_),
    .B2(_0436_),
    .A2(net128),
    .A1(_0100_));
 sg13g2_nor2b_2 _1148_ (.A(_0235_),
    .B_N(_0179_),
    .Y(_0437_));
 sg13g2_o21ai_1 _1149_ (.B1(_0252_),
    .Y(_0438_),
    .A1(_0253_),
    .A2(_0255_));
 sg13g2_nor2_1 _1150_ (.A(net141),
    .B(_0256_),
    .Y(_0439_));
 sg13g2_nand2_1 _1151_ (.Y(_0440_),
    .A(_0438_),
    .B(_0439_));
 sg13g2_a22oi_1 _1152_ (.Y(_0026_),
    .B1(_0437_),
    .B2(_0440_),
    .A2(net128),
    .A1(_0102_));
 sg13g2_a21o_1 _1153_ (.A2(net144),
    .A1(\raster.tscan.left_x[4] ),
    .B1(_0256_),
    .X(_0441_));
 sg13g2_a21oi_1 _1154_ (.A1(_0251_),
    .A2(_0441_),
    .Y(_0442_),
    .B1(net141));
 sg13g2_o21ai_1 _1155_ (.B1(_0442_),
    .Y(_0443_),
    .A1(_0251_),
    .A2(_0441_));
 sg13g2_a22oi_1 _1156_ (.Y(_0444_),
    .B1(_0437_),
    .B2(_0443_),
    .A2(net128),
    .A1(net200));
 sg13g2_inv_1 _1157_ (.Y(_0027_),
    .A(net201));
 sg13g2_o21ai_1 _1158_ (.B1(_0260_),
    .Y(_0445_),
    .A1(_0257_),
    .A2(_0263_));
 sg13g2_nor3_1 _1159_ (.A(_0257_),
    .B(_0260_),
    .C(_0263_),
    .Y(_0446_));
 sg13g2_nor2_1 _1160_ (.A(_0111_),
    .B(_0446_),
    .Y(_0447_));
 sg13g2_a221oi_1 _1161_ (.B2(_0447_),
    .C1(net129),
    .B1(_0445_),
    .A1(net160),
    .Y(_0448_),
    .A2(_0228_));
 sg13g2_a21oi_1 _1162_ (.A1(_0103_),
    .A2(net129),
    .Y(_0028_),
    .B1(_0448_));
 sg13g2_nand2_1 _1163_ (.Y(_0449_),
    .A(net189),
    .B(net129));
 sg13g2_nand2_1 _1164_ (.Y(_0450_),
    .A(_0259_),
    .B(_0445_));
 sg13g2_xor2_1 _1165_ (.B(_0450_),
    .A(_0258_),
    .X(_0451_));
 sg13g2_nor2_1 _1166_ (.A(net142),
    .B(_0451_),
    .Y(_0452_));
 sg13g2_o21ai_1 _1167_ (.B1(_0449_),
    .Y(_0029_),
    .A1(_0430_),
    .A2(_0452_));
 sg13g2_nand3_1 _1168_ (.B(_0261_),
    .C(_0265_),
    .A(_0250_),
    .Y(_0453_));
 sg13g2_nand3_1 _1169_ (.B(_0266_),
    .C(_0453_),
    .A(net137),
    .Y(_0454_));
 sg13g2_a22oi_1 _1170_ (.Y(_0030_),
    .B1(_0433_),
    .B2(_0454_),
    .A2(net129),
    .A1(_0104_));
 sg13g2_o21ai_1 _1171_ (.B1(net158),
    .Y(_0455_),
    .A1(net177),
    .A2(net179));
 sg13g2_and2_1 _1172_ (.A(_0314_),
    .B(_0455_),
    .X(_0456_));
 sg13g2_nand2_1 _1173_ (.Y(_0457_),
    .A(_0330_),
    .B(_0455_));
 sg13g2_and2_1 _1174_ (.A(net168),
    .B(_0457_),
    .X(_0458_));
 sg13g2_nor2_1 _1175_ (.A(net161),
    .B(_0331_),
    .Y(_0459_));
 sg13g2_nand2_1 _1176_ (.Y(_0460_),
    .A(\raster.tscan.left_err[4] ),
    .B(_0459_));
 sg13g2_and2_1 _1177_ (.A(\raster.tscan.left_err[3] ),
    .B(_0456_),
    .X(_0461_));
 sg13g2_nand3_1 _1178_ (.B(net162),
    .C(_0303_),
    .A(\raster.tscan.left_err[2] ),
    .Y(_0462_));
 sg13g2_a21oi_1 _1179_ (.A1(_0149_),
    .A2(_0455_),
    .Y(_0463_),
    .B1(_0093_));
 sg13g2_nand3_1 _1180_ (.B(_0149_),
    .C(_0455_),
    .A(_0093_),
    .Y(_0464_));
 sg13g2_nor2b_1 _1181_ (.A(_0463_),
    .B_N(_0464_),
    .Y(_0465_));
 sg13g2_a21oi_1 _1182_ (.A1(_0421_),
    .A2(_0464_),
    .Y(_0466_),
    .B1(_0463_));
 sg13g2_a21o_1 _1183_ (.A2(_0303_),
    .A1(net162),
    .B1(\raster.tscan.left_err[2] ),
    .X(_0467_));
 sg13g2_nand2_1 _1184_ (.Y(_0468_),
    .A(_0462_),
    .B(_0467_));
 sg13g2_o21ai_1 _1185_ (.B1(_0462_),
    .Y(_0469_),
    .A1(_0466_),
    .A2(_0468_));
 sg13g2_xnor2_1 _1186_ (.Y(_0470_),
    .A(_0094_),
    .B(_0456_));
 sg13g2_a21oi_1 _1187_ (.A1(_0469_),
    .A2(_0470_),
    .Y(_0471_),
    .B1(_0461_));
 sg13g2_xnor2_1 _1188_ (.Y(_0472_),
    .A(\raster.tscan.left_err[4] ),
    .B(_0459_));
 sg13g2_o21ai_1 _1189_ (.B1(_0460_),
    .Y(_0473_),
    .A1(_0471_),
    .A2(_0472_));
 sg13g2_xor2_1 _1190_ (.B(_0457_),
    .A(net168),
    .X(_0474_));
 sg13g2_a21oi_2 _1191_ (.B1(_0458_),
    .Y(_0475_),
    .A2(_0474_),
    .A1(_0473_));
 sg13g2_nand2_1 _1192_ (.Y(_0476_),
    .A(\raster.tscan.left_err[6] ),
    .B(net161));
 sg13g2_nand2_1 _1193_ (.Y(_0477_),
    .A(net159),
    .B(\raster.tscan.left_err[6] ));
 sg13g2_xor2_1 _1194_ (.B(\raster.tscan.left_err[6] ),
    .A(net159),
    .X(_0478_));
 sg13g2_o21ai_1 _1195_ (.B1(_0476_),
    .Y(_0479_),
    .A1(net161),
    .A2(_0478_));
 sg13g2_nand2_1 _1196_ (.Y(_0480_),
    .A(\raster.tscan.left_err[7] ),
    .B(_0455_));
 sg13g2_xnor2_1 _1197_ (.Y(_0481_),
    .A(net197),
    .B(_0455_));
 sg13g2_or2_1 _1198_ (.X(_0482_),
    .B(_0481_),
    .A(_0479_));
 sg13g2_o21ai_1 _1199_ (.B1(\raster.tscan.left_err[6] ),
    .Y(_0483_),
    .A1(net159),
    .A2(net161));
 sg13g2_nand2_1 _1200_ (.Y(_0484_),
    .A(_0480_),
    .B(_0483_));
 sg13g2_o21ai_1 _1201_ (.B1(_0484_),
    .Y(_0485_),
    .A1(\raster.tscan.left_err[7] ),
    .A2(_0455_));
 sg13g2_o21ai_1 _1202_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_0475_),
    .A2(_0482_));
 sg13g2_a21oi_1 _1203_ (.A1(net172),
    .A2(net162),
    .Y(_0487_),
    .B1(_0486_));
 sg13g2_mux2_1 _1204_ (.A0(net162),
    .A1(_0486_),
    .S(_0097_),
    .X(_0488_));
 sg13g2_o21ai_1 _1205_ (.B1(_0234_),
    .Y(_0489_),
    .A1(_0487_),
    .A2(_0488_));
 sg13g2_nand2_1 _1206_ (.Y(_0490_),
    .A(_0178_),
    .B(_0273_));
 sg13g2_nor2_1 _1207_ (.A(net148),
    .B(_0096_),
    .Y(_0491_));
 sg13g2_nor2_1 _1208_ (.A(net159),
    .B(\raster.tscan.left_err[7] ),
    .Y(_0492_));
 sg13g2_nand2_1 _1209_ (.Y(_0493_),
    .A(net158),
    .B(\raster.tscan.left_err[3] ));
 sg13g2_nor2_1 _1210_ (.A(net158),
    .B(\raster.tscan.left_err[3] ),
    .Y(_0494_));
 sg13g2_xor2_1 _1211_ (.B(\raster.tscan.left_err[3] ),
    .A(net158),
    .X(_0495_));
 sg13g2_nor2_1 _1212_ (.A(\raster.tscan.left_err[1] ),
    .B(\raster.tscan.left_err[2] ),
    .Y(_0496_));
 sg13g2_o21ai_1 _1213_ (.B1(_0493_),
    .Y(_0497_),
    .A1(_0494_),
    .A2(_0496_));
 sg13g2_and2_1 _1214_ (.A(\raster.tscan.left_err[4] ),
    .B(_0497_),
    .X(_0498_));
 sg13g2_nand2_1 _1215_ (.Y(_0499_),
    .A(net168),
    .B(_0498_));
 sg13g2_nand3_1 _1216_ (.B(_0478_),
    .C(_0498_),
    .A(\raster.tscan.left_err[5] ),
    .Y(_0500_));
 sg13g2_a21oi_1 _1217_ (.A1(_0477_),
    .A2(_0500_),
    .Y(_0501_),
    .B1(_0492_));
 sg13g2_nor3_1 _1218_ (.A(\raster.tscan.left_err[8] ),
    .B(_0491_),
    .C(_0501_),
    .Y(_0502_));
 sg13g2_and2_1 _1219_ (.A(net205),
    .B(_0502_),
    .X(_0503_));
 sg13g2_o21ai_1 _1220_ (.B1(_0419_),
    .Y(_0504_),
    .A1(_0083_),
    .A2(_0503_));
 sg13g2_or2_1 _1221_ (.X(_0505_),
    .B(_0492_),
    .A(_0491_));
 sg13g2_inv_1 _1222_ (.Y(_0506_),
    .A(_0505_));
 sg13g2_nand2_1 _1223_ (.Y(_0507_),
    .A(net148),
    .B(net168));
 sg13g2_xor2_1 _1224_ (.B(net168),
    .A(net159),
    .X(_0508_));
 sg13g2_and2_1 _1225_ (.A(net158),
    .B(\raster.tscan.left_err[2] ),
    .X(_0509_));
 sg13g2_xor2_1 _1226_ (.B(\raster.tscan.left_err[2] ),
    .A(net158),
    .X(_0510_));
 sg13g2_a21oi_1 _1227_ (.A1(\raster.tscan.left_err[1] ),
    .A2(_0510_),
    .Y(_0511_),
    .B1(_0509_));
 sg13g2_a21o_1 _1228_ (.A2(_0510_),
    .A1(\raster.tscan.left_err[1] ),
    .B1(_0509_),
    .X(_0512_));
 sg13g2_a21oi_1 _1229_ (.A1(_0094_),
    .A2(_0511_),
    .Y(_0513_),
    .B1(_0095_));
 sg13g2_o21ai_1 _1230_ (.B1(\raster.tscan.left_err[4] ),
    .Y(_0514_),
    .A1(\raster.tscan.left_err[3] ),
    .A2(_0512_));
 sg13g2_o21ai_1 _1231_ (.B1(_0507_),
    .Y(_0515_),
    .A1(_0508_),
    .A2(_0514_));
 sg13g2_o21ai_1 _1232_ (.B1(_0506_),
    .Y(_0516_),
    .A1(\raster.tscan.left_err[6] ),
    .A2(_0515_));
 sg13g2_o21ai_1 _1233_ (.B1(_0502_),
    .Y(_0517_),
    .A1(net172),
    .A2(_0516_));
 sg13g2_a221oi_1 _1234_ (.B2(_0084_),
    .C1(net136),
    .B1(_0517_),
    .A1(_0503_),
    .Y(_0518_),
    .A2(_0516_));
 sg13g2_a21oi_1 _1235_ (.A1(_0504_),
    .A2(_0518_),
    .Y(_0519_),
    .B1(_0490_));
 sg13g2_a22oi_1 _1236_ (.Y(_0031_),
    .B1(_0519_),
    .B2(_0489_),
    .A2(_0490_),
    .A1(_0084_));
 sg13g2_nor2_1 _1237_ (.A(_0230_),
    .B(_0231_),
    .Y(_0520_));
 sg13g2_nand3b_1 _1238_ (.B(_0274_),
    .C(_0520_),
    .Y(_0521_),
    .A_N(_0181_));
 sg13g2_a21oi_2 _1239_ (.B1(_0521_),
    .Y(_0522_),
    .A2(_0236_),
    .A1(_0156_));
 sg13g2_a21o_2 _1240_ (.A2(_0236_),
    .A1(_0156_),
    .B1(_0521_),
    .X(_0523_));
 sg13g2_nor2_2 _1241_ (.A(_0228_),
    .B(net127),
    .Y(_0524_));
 sg13g2_nand2_1 _1242_ (.Y(_0525_),
    .A(net175),
    .B(net194));
 sg13g2_nor2_1 _1243_ (.A(net175),
    .B(\raster.tscan.right_x[2] ),
    .Y(_0526_));
 sg13g2_xnor2_1 _1244_ (.Y(_0527_),
    .A(net175),
    .B(net194));
 sg13g2_and2_1 _1245_ (.A(net175),
    .B(net108),
    .X(_0528_));
 sg13g2_xor2_1 _1246_ (.B(net108),
    .A(net177),
    .X(_0529_));
 sg13g2_a21oi_1 _1247_ (.A1(net92),
    .A2(_0529_),
    .Y(_0530_),
    .B1(_0528_));
 sg13g2_a21oi_1 _1248_ (.A1(_0527_),
    .A2(_0530_),
    .Y(_0531_),
    .B1(net141));
 sg13g2_o21ai_1 _1249_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0527_),
    .A2(_0530_));
 sg13g2_a22oi_1 _1250_ (.Y(_0032_),
    .B1(_0524_),
    .B2(_0532_),
    .A2(net127),
    .A1(_0088_));
 sg13g2_nor2_1 _1251_ (.A(net141),
    .B(net127),
    .Y(_0533_));
 sg13g2_nand2_2 _1252_ (.Y(_0534_),
    .A(net137),
    .B(_0522_));
 sg13g2_o21ai_1 _1253_ (.B1(_0525_),
    .Y(_0535_),
    .A1(_0526_),
    .A2(_0530_));
 sg13g2_nand2_1 _1254_ (.Y(_0536_),
    .A(net175),
    .B(net209));
 sg13g2_xor2_1 _1255_ (.B(net209),
    .A(net175),
    .X(_0537_));
 sg13g2_xnor2_1 _1256_ (.Y(_0538_),
    .A(_0535_),
    .B(_0537_));
 sg13g2_a22oi_1 _1257_ (.Y(_0539_),
    .B1(_0423_),
    .B2(net179),
    .A2(_0228_),
    .A1(net160));
 sg13g2_nor2_1 _1258_ (.A(net127),
    .B(_0539_),
    .Y(_0540_));
 sg13g2_nand3_1 _1259_ (.B(_0423_),
    .C(_0522_),
    .A(net213),
    .Y(_0541_));
 sg13g2_a221oi_1 _1260_ (.B2(_0538_),
    .C1(_0540_),
    .B1(_0533_),
    .A1(_0089_),
    .Y(_0033_),
    .A2(net127));
 sg13g2_xnor2_1 _1261_ (.Y(_0542_),
    .A(net175),
    .B(\raster.tscan.right_x[4] ));
 sg13g2_o21ai_1 _1262_ (.B1(_0535_),
    .Y(_0543_),
    .A1(net175),
    .A2(\raster.tscan.right_x[3] ));
 sg13g2_nand3_1 _1263_ (.B(_0542_),
    .C(_0543_),
    .A(_0536_),
    .Y(_0544_));
 sg13g2_a21o_2 _1264_ (.A2(_0543_),
    .A1(_0536_),
    .B1(_0542_),
    .X(_0545_));
 sg13g2_nand4_1 _1265_ (.B(_0522_),
    .C(_0544_),
    .A(net137),
    .Y(_0546_),
    .D(_0545_));
 sg13g2_nand2_1 _1266_ (.Y(_0547_),
    .A(\raster.tscan.right_x[4] ),
    .B(net126));
 sg13g2_nand3_1 _1267_ (.B(_0546_),
    .C(_0547_),
    .A(_0541_),
    .Y(_0034_));
 sg13g2_xnor2_1 _1268_ (.Y(_0548_),
    .A(net176),
    .B(net183));
 sg13g2_o21ai_1 _1269_ (.B1(_0545_),
    .Y(_0549_),
    .A1(_0081_),
    .A2(_0090_));
 sg13g2_xnor2_1 _1270_ (.Y(_0550_),
    .A(_0548_),
    .B(_0549_));
 sg13g2_nand2_1 _1271_ (.Y(_0551_),
    .A(net138),
    .B(_0550_));
 sg13g2_a22oi_1 _1272_ (.Y(_0035_),
    .B1(_0524_),
    .B2(_0551_),
    .A2(net127),
    .A1(_0091_));
 sg13g2_nor2_1 _1273_ (.A(_0423_),
    .B(net126),
    .Y(_0552_));
 sg13g2_nand2_1 _1274_ (.Y(_0553_),
    .A(net176),
    .B(\raster.tscan.right_x[6] ));
 sg13g2_xnor2_1 _1275_ (.Y(_0554_),
    .A(net176),
    .B(\raster.tscan.right_x[6] ));
 sg13g2_o21ai_1 _1276_ (.B1(net176),
    .Y(_0555_),
    .A1(\raster.tscan.right_x[4] ),
    .A2(\raster.tscan.right_x[5] ));
 sg13g2_nor2_1 _1277_ (.A(_0545_),
    .B(_0548_),
    .Y(_0556_));
 sg13g2_nor2b_1 _1278_ (.A(_0556_),
    .B_N(_0555_),
    .Y(_0557_));
 sg13g2_xor2_1 _1279_ (.B(_0557_),
    .A(_0554_),
    .X(_0558_));
 sg13g2_nor2_1 _1280_ (.A(net140),
    .B(_0558_),
    .Y(_0559_));
 sg13g2_nor3_1 _1281_ (.A(_0423_),
    .B(net126),
    .C(_0559_),
    .Y(_0560_));
 sg13g2_a21o_1 _1282_ (.A2(net126),
    .A1(net203),
    .B1(_0560_),
    .X(_0036_));
 sg13g2_and2_1 _1283_ (.A(net227),
    .B(net126),
    .X(_0561_));
 sg13g2_xnor2_1 _1284_ (.Y(_0562_),
    .A(net176),
    .B(\raster.tscan.right_x[7] ));
 sg13g2_o21ai_1 _1285_ (.B1(_0553_),
    .Y(_0563_),
    .A1(_0554_),
    .A2(_0557_));
 sg13g2_o21ai_1 _1286_ (.B1(net138),
    .Y(_0564_),
    .A1(_0562_),
    .A2(_0563_));
 sg13g2_a21o_1 _1287_ (.A2(_0563_),
    .A1(_0562_),
    .B1(_0564_),
    .X(_0565_));
 sg13g2_a21o_1 _1288_ (.A2(_0565_),
    .A1(_0524_),
    .B1(_0561_),
    .X(_0037_));
 sg13g2_nor2_1 _1289_ (.A(_0081_),
    .B(_0092_),
    .Y(_0566_));
 sg13g2_nand2_1 _1290_ (.Y(_0567_),
    .A(_0081_),
    .B(_0092_));
 sg13g2_nand2b_1 _1291_ (.Y(_0568_),
    .B(_0567_),
    .A_N(_0566_));
 sg13g2_nor4_1 _1292_ (.A(_0545_),
    .B(_0548_),
    .C(_0554_),
    .D(_0562_),
    .Y(_0569_));
 sg13g2_o21ai_1 _1293_ (.B1(net176),
    .Y(_0570_),
    .A1(\raster.tscan.right_x[6] ),
    .A2(\raster.tscan.right_x[7] ));
 sg13g2_nand3b_1 _1294_ (.B(_0570_),
    .C(_0555_),
    .Y(_0571_),
    .A_N(_0569_));
 sg13g2_xnor2_1 _1295_ (.Y(_0572_),
    .A(_0568_),
    .B(_0571_));
 sg13g2_nand2_1 _1296_ (.Y(_0573_),
    .A(net137),
    .B(_0572_));
 sg13g2_a22oi_1 _1297_ (.Y(_0038_),
    .B1(_0552_),
    .B2(_0573_),
    .A2(net126),
    .A1(_0092_));
 sg13g2_nand2_1 _1298_ (.Y(_0574_),
    .A(net191),
    .B(net134));
 sg13g2_a21o_1 _1299_ (.A2(_0408_),
    .A1(net145),
    .B1(_0574_),
    .X(_0575_));
 sg13g2_xor2_1 _1300_ (.B(_0411_),
    .A(net191),
    .X(_0576_));
 sg13g2_xnor2_1 _1301_ (.Y(_0577_),
    .A(\raster.tscan.right_err[9] ),
    .B(_0413_));
 sg13g2_and2_1 _1302_ (.A(_0311_),
    .B(_0577_),
    .X(_0578_));
 sg13g2_a22oi_1 _1303_ (.Y(_0579_),
    .B1(_0578_),
    .B2(net140),
    .A2(_0576_),
    .A1(_0385_));
 sg13g2_and2_1 _1304_ (.A(_0275_),
    .B(_0579_),
    .X(_0580_));
 sg13g2_nor2_1 _1305_ (.A(net191),
    .B(_0275_),
    .Y(_0581_));
 sg13g2_a21oi_1 _1306_ (.A1(_0575_),
    .A2(_0580_),
    .Y(_0039_),
    .B1(_0581_));
 sg13g2_or3_1 _1307_ (.A(_0170_),
    .B(_0272_),
    .C(_0418_),
    .X(_0582_));
 sg13g2_xnor2_1 _1308_ (.Y(_0583_),
    .A(_0421_),
    .B(_0465_));
 sg13g2_a21o_1 _1309_ (.A2(_0218_),
    .A1(_0177_),
    .B1(net228),
    .X(_0584_));
 sg13g2_a21oi_1 _1310_ (.A1(_0182_),
    .A2(_0303_),
    .Y(_0585_),
    .B1(net135));
 sg13g2_a22oi_1 _1311_ (.Y(_0586_),
    .B1(_0584_),
    .B2(_0585_),
    .A2(_0583_),
    .A1(net134));
 sg13g2_mux2_1 _1312_ (.A0(_0586_),
    .A1(net228),
    .S(net122),
    .X(_0040_));
 sg13g2_xnor2_1 _1313_ (.Y(_0587_),
    .A(_0466_),
    .B(_0468_));
 sg13g2_nand2_1 _1314_ (.Y(_0588_),
    .A(net135),
    .B(_0587_));
 sg13g2_xnor2_1 _1315_ (.Y(_0589_),
    .A(\raster.tscan.left_err[1] ),
    .B(_0510_));
 sg13g2_xnor2_1 _1316_ (.Y(_0590_),
    .A(\raster.tscan.left_err[1] ),
    .B(\raster.tscan.left_err[2] ));
 sg13g2_a221oi_1 _1317_ (.B2(net171),
    .C1(_0318_),
    .B1(_0590_),
    .A1(_0182_),
    .Y(_0591_),
    .A2(_0314_));
 sg13g2_o21ai_1 _1318_ (.B1(_0591_),
    .Y(_0592_),
    .A1(_0419_),
    .A2(_0589_));
 sg13g2_and2_1 _1319_ (.A(_0588_),
    .B(_0592_),
    .X(_0593_));
 sg13g2_mux2_1 _1320_ (.A0(_0593_),
    .A1(net220),
    .S(net122),
    .X(_0041_));
 sg13g2_xnor2_1 _1321_ (.Y(_0594_),
    .A(_0469_),
    .B(_0470_));
 sg13g2_nand2_1 _1322_ (.Y(_0595_),
    .A(net135),
    .B(_0594_));
 sg13g2_xnor2_1 _1323_ (.Y(_0596_),
    .A(net222),
    .B(_0511_));
 sg13g2_xnor2_1 _1324_ (.Y(_0597_),
    .A(_0495_),
    .B(_0496_));
 sg13g2_a221oi_1 _1325_ (.B2(net171),
    .C1(net135),
    .B1(_0597_),
    .A1(_0182_),
    .Y(_0598_),
    .A2(_0332_));
 sg13g2_o21ai_1 _1326_ (.B1(_0598_),
    .Y(_0599_),
    .A1(_0419_),
    .A2(_0596_));
 sg13g2_a21oi_1 _1327_ (.A1(_0595_),
    .A2(_0599_),
    .Y(_0600_),
    .B1(net122));
 sg13g2_a21oi_1 _1328_ (.A1(_0094_),
    .A2(net122),
    .Y(_0042_),
    .B1(_0600_));
 sg13g2_xnor2_1 _1329_ (.Y(_0601_),
    .A(_0471_),
    .B(_0472_));
 sg13g2_nor3_1 _1330_ (.A(\raster.tscan.left_err[3] ),
    .B(\raster.tscan.left_err[4] ),
    .C(_0512_),
    .Y(_0602_));
 sg13g2_nor3_1 _1331_ (.A(_0419_),
    .B(_0513_),
    .C(_0602_),
    .Y(_0603_));
 sg13g2_nor3_1 _1332_ (.A(_0082_),
    .B(_0167_),
    .C(_0330_),
    .Y(_0604_));
 sg13g2_nor2_1 _1333_ (.A(\raster.tscan.left_err[4] ),
    .B(_0497_),
    .Y(_0605_));
 sg13g2_nor3_1 _1334_ (.A(_0083_),
    .B(_0498_),
    .C(_0605_),
    .Y(_0606_));
 sg13g2_nor4_1 _1335_ (.A(_0424_),
    .B(_0603_),
    .C(_0604_),
    .D(_0606_),
    .Y(_0607_));
 sg13g2_a21oi_1 _1336_ (.A1(net135),
    .A2(_0601_),
    .Y(_0608_),
    .B1(_0607_));
 sg13g2_mux2_1 _1337_ (.A0(_0608_),
    .A1(net221),
    .S(net122),
    .X(_0043_));
 sg13g2_xnor2_1 _1338_ (.Y(_0609_),
    .A(_0473_),
    .B(_0474_));
 sg13g2_xnor2_1 _1339_ (.Y(_0610_),
    .A(_0508_),
    .B(_0513_));
 sg13g2_nand2b_1 _1340_ (.Y(_0611_),
    .B(_0610_),
    .A_N(_0419_));
 sg13g2_a21oi_1 _1341_ (.A1(net168),
    .A2(_0498_),
    .Y(_0612_),
    .B1(_0083_));
 sg13g2_o21ai_1 _1342_ (.B1(_0612_),
    .Y(_0613_),
    .A1(net168),
    .A2(_0498_));
 sg13g2_nand2b_1 _1343_ (.Y(_0614_),
    .B(_0613_),
    .A_N(_0289_));
 sg13g2_a21oi_1 _1344_ (.A1(net158),
    .A2(_0182_),
    .Y(_0615_),
    .B1(_0614_));
 sg13g2_a221oi_1 _1345_ (.B2(_0615_),
    .C1(net123),
    .B1(_0611_),
    .A1(net136),
    .Y(_0616_),
    .A2(_0609_));
 sg13g2_a21o_1 _1346_ (.A2(net122),
    .A1(net168),
    .B1(_0616_),
    .X(_0044_));
 sg13g2_xnor2_1 _1347_ (.Y(_0617_),
    .A(_0475_),
    .B(_0479_));
 sg13g2_xnor2_1 _1348_ (.Y(_0618_),
    .A(\raster.tscan.left_err[6] ),
    .B(_0515_));
 sg13g2_xnor2_1 _1349_ (.Y(_0619_),
    .A(_0478_),
    .B(_0499_));
 sg13g2_a221oi_1 _1350_ (.B2(net172),
    .C1(_0318_),
    .B1(_0619_),
    .A1(net161),
    .Y(_0620_),
    .A2(_0618_));
 sg13g2_a22oi_1 _1351_ (.Y(_0621_),
    .B1(_0620_),
    .B2(_0183_),
    .A2(_0617_),
    .A1(net136));
 sg13g2_mux2_1 _1352_ (.A0(_0621_),
    .A1(net226),
    .S(net122),
    .X(_0045_));
 sg13g2_o21ai_1 _1353_ (.B1(_0483_),
    .Y(_0622_),
    .A1(_0475_),
    .A2(_0479_));
 sg13g2_xnor2_1 _1354_ (.Y(_0623_),
    .A(_0481_),
    .B(_0622_));
 sg13g2_nand2_1 _1355_ (.Y(_0624_),
    .A(net135),
    .B(_0623_));
 sg13g2_nor3_1 _1356_ (.A(\raster.tscan.left_err[6] ),
    .B(_0506_),
    .C(_0515_),
    .Y(_0625_));
 sg13g2_nor2_1 _1357_ (.A(_0219_),
    .B(_0625_),
    .Y(_0626_));
 sg13g2_a21oi_1 _1358_ (.A1(_0477_),
    .A2(_0500_),
    .Y(_0627_),
    .B1(_0505_));
 sg13g2_nand3_1 _1359_ (.B(_0500_),
    .C(_0505_),
    .A(_0477_),
    .Y(_0628_));
 sg13g2_nor2_1 _1360_ (.A(_0083_),
    .B(_0627_),
    .Y(_0629_));
 sg13g2_a22oi_1 _1361_ (.Y(_0630_),
    .B1(_0628_),
    .B2(_0629_),
    .A2(_0626_),
    .A1(_0516_));
 sg13g2_nand2_1 _1362_ (.Y(_0631_),
    .A(_0183_),
    .B(_0630_));
 sg13g2_a21oi_1 _1363_ (.A1(net142),
    .A2(_0631_),
    .Y(_0632_),
    .B1(net122));
 sg13g2_a22oi_1 _1364_ (.Y(_0046_),
    .B1(_0624_),
    .B2(_0632_),
    .A2(net123),
    .A1(_0096_));
 sg13g2_xnor2_1 _1365_ (.Y(_0633_),
    .A(_0097_),
    .B(_0219_));
 sg13g2_o21ai_1 _1366_ (.B1(net136),
    .Y(_0634_),
    .A1(_0486_),
    .A2(_0633_));
 sg13g2_a21o_1 _1367_ (.A2(_0633_),
    .A1(_0486_),
    .B1(_0634_),
    .X(_0635_));
 sg13g2_nand2b_1 _1368_ (.Y(_0636_),
    .B(_0516_),
    .A_N(_0491_));
 sg13g2_xnor2_1 _1369_ (.Y(_0637_),
    .A(\raster.tscan.left_err[8] ),
    .B(_0636_));
 sg13g2_o21ai_1 _1370_ (.B1(\raster.tscan.left_err[8] ),
    .Y(_0638_),
    .A1(_0491_),
    .A2(_0501_));
 sg13g2_nand2b_1 _1371_ (.Y(_0639_),
    .B(_0638_),
    .A_N(_0502_));
 sg13g2_a22oi_1 _1372_ (.Y(_0640_),
    .B1(_0639_),
    .B2(net172),
    .A2(_0637_),
    .A1(net161));
 sg13g2_nand2_1 _1373_ (.Y(_0641_),
    .A(_0183_),
    .B(_0640_));
 sg13g2_a21oi_1 _1374_ (.A1(net142),
    .A2(_0641_),
    .Y(_0642_),
    .B1(net123));
 sg13g2_a22oi_1 _1375_ (.Y(_0047_),
    .B1(_0635_),
    .B2(_0642_),
    .A2(net123),
    .A1(_0097_));
 sg13g2_and3_1 _1376_ (.X(_0643_),
    .A(net219),
    .B(net185),
    .C(net118));
 sg13g2_and2_1 _1377_ (.A(net223),
    .B(_0643_),
    .X(_0644_));
 sg13g2_nand2_1 _1378_ (.Y(_0645_),
    .A(net231),
    .B(_0644_));
 sg13g2_nor3_1 _1379_ (.A(\raster.hpos[5] ),
    .B(\raster.hpos[7] ),
    .C(net167),
    .Y(_0646_));
 sg13g2_nand3_1 _1380_ (.B(net166),
    .C(_0646_),
    .A(\raster.hpos[9] ),
    .Y(_0647_));
 sg13g2_nor2_1 _1381_ (.A(_0645_),
    .B(_0647_),
    .Y(_0648_));
 sg13g2_nor2b_1 _1382_ (.A(_0648_),
    .B_N(net1),
    .Y(_0649_));
 sg13g2_nand2b_2 _1383_ (.Y(_0650_),
    .B(net180),
    .A_N(_0648_));
 sg13g2_nor2_1 _1384_ (.A(net185),
    .B(_0650_),
    .Y(_0048_));
 sg13g2_xnor2_1 _1385_ (.Y(_0651_),
    .A(net219),
    .B(net185));
 sg13g2_nor2_1 _1386_ (.A(_0650_),
    .B(_0651_),
    .Y(_0049_));
 sg13g2_a21oi_1 _1387_ (.A1(\raster.hpos[1] ),
    .A2(\raster.hpos[0] ),
    .Y(_0652_),
    .B1(net118));
 sg13g2_nor3_1 _1388_ (.A(_0643_),
    .B(_0650_),
    .C(net119),
    .Y(_0050_));
 sg13g2_o21ai_1 _1389_ (.B1(net1),
    .Y(_0653_),
    .A1(net223),
    .A2(_0643_));
 sg13g2_nor2_1 _1390_ (.A(_0644_),
    .B(_0653_),
    .Y(_0051_));
 sg13g2_o21ai_1 _1391_ (.B1(net1),
    .Y(_0654_),
    .A1(net231),
    .A2(_0644_));
 sg13g2_nor2b_1 _1392_ (.A(_0654_),
    .B_N(_0645_),
    .Y(_0052_));
 sg13g2_a21oi_1 _1393_ (.A1(\raster.hpos[4] ),
    .A2(_0644_),
    .Y(_0655_),
    .B1(net112));
 sg13g2_nor2_1 _1394_ (.A(_0076_),
    .B(_0645_),
    .Y(_0656_));
 sg13g2_nor3_1 _1395_ (.A(_0650_),
    .B(net113),
    .C(_0656_),
    .Y(_0053_));
 sg13g2_nor2_1 _1396_ (.A(net167),
    .B(_0656_),
    .Y(_0657_));
 sg13g2_and2_1 _1397_ (.A(net167),
    .B(_0656_),
    .X(_0658_));
 sg13g2_nor3_1 _1398_ (.A(_0650_),
    .B(_0657_),
    .C(_0658_),
    .Y(_0054_));
 sg13g2_and2_1 _1399_ (.A(net224),
    .B(_0658_),
    .X(_0659_));
 sg13g2_o21ai_1 _1400_ (.B1(net132),
    .Y(_0660_),
    .A1(net224),
    .A2(_0658_));
 sg13g2_nor2_1 _1401_ (.A(_0659_),
    .B(net225),
    .Y(_0055_));
 sg13g2_and2_1 _1402_ (.A(net166),
    .B(_0659_),
    .X(_0661_));
 sg13g2_o21ai_1 _1403_ (.B1(net132),
    .Y(_0662_),
    .A1(net166),
    .A2(_0659_));
 sg13g2_nor2_1 _1404_ (.A(_0661_),
    .B(_0662_),
    .Y(_0056_));
 sg13g2_a21oi_1 _1405_ (.A1(net230),
    .A2(_0661_),
    .Y(_0663_),
    .B1(_0650_));
 sg13g2_o21ai_1 _1406_ (.B1(_0663_),
    .Y(_0664_),
    .A1(net230),
    .A2(_0661_));
 sg13g2_inv_1 _1407_ (.Y(_0057_),
    .A(_0664_));
 sg13g2_nand2_1 _1408_ (.Y(_0665_),
    .A(net92),
    .B(net127));
 sg13g2_o21ai_1 _1409_ (.B1(_0665_),
    .Y(_0058_),
    .A1(net92),
    .A2(_0534_));
 sg13g2_nand2_1 _1410_ (.Y(_0666_),
    .A(net108),
    .B(net126));
 sg13g2_xnor2_1 _1411_ (.Y(_0667_),
    .A(net92),
    .B(_0529_));
 sg13g2_o21ai_1 _1412_ (.B1(_0666_),
    .Y(_0059_),
    .A1(_0534_),
    .A2(_0667_));
 sg13g2_nand2_1 _1413_ (.Y(_0668_),
    .A(net101),
    .B(net126));
 sg13g2_a21oi_1 _1414_ (.A1(_0567_),
    .A2(_0571_),
    .Y(_0669_),
    .B1(_0566_));
 sg13g2_xnor2_1 _1415_ (.Y(_0670_),
    .A(net176),
    .B(net101));
 sg13g2_xnor2_1 _1416_ (.Y(_0671_),
    .A(_0669_),
    .B(_0670_));
 sg13g2_o21ai_1 _1417_ (.B1(_0668_),
    .Y(_0060_),
    .A1(_0534_),
    .A2(_0671_));
 sg13g2_nand2_1 _1418_ (.Y(_0672_),
    .A(net180),
    .B(_0648_));
 sg13g2_nor4_1 _1419_ (.A(\raster.hvsync_gen.vpos[6] ),
    .B(\raster.hvsync_gen.vpos[7] ),
    .C(\raster.hvsync_gen.vpos[8] ),
    .D(_0080_),
    .Y(_0673_));
 sg13g2_nand3_1 _1420_ (.B(\raster.hvsync_gen.vpos[3] ),
    .C(_0147_),
    .A(\raster.hvsync_gen.vpos[2] ),
    .Y(_0674_));
 sg13g2_nor3_1 _1421_ (.A(\raster.hvsync_gen.vpos[4] ),
    .B(\raster.hvsync_gen.vpos[5] ),
    .C(_0674_),
    .Y(_0675_));
 sg13g2_a21o_2 _1422_ (.A2(_0675_),
    .A1(_0673_),
    .B1(_0672_),
    .X(_0676_));
 sg13g2_nor2b_1 _1423_ (.A(net89),
    .B_N(net130),
    .Y(_0677_));
 sg13g2_a21oi_1 _1424_ (.A1(net89),
    .A2(_0650_),
    .Y(_0061_),
    .B1(_0677_));
 sg13g2_nand2_1 _1425_ (.Y(_0678_),
    .A(net93),
    .B(net131));
 sg13g2_o21ai_1 _1426_ (.B1(_0678_),
    .Y(_0062_),
    .A1(_0148_),
    .A2(_0672_));
 sg13g2_nand2_1 _1427_ (.Y(_0679_),
    .A(net99),
    .B(net131));
 sg13g2_o21ai_1 _1428_ (.B1(_0679_),
    .Y(_0063_),
    .A1(_0138_),
    .A2(net130));
 sg13g2_nand2_1 _1429_ (.Y(_0680_),
    .A(net188),
    .B(net131));
 sg13g2_o21ai_1 _1430_ (.B1(_0680_),
    .Y(_0064_),
    .A1(_0133_),
    .A2(net130));
 sg13g2_nand2_1 _1431_ (.Y(_0681_),
    .A(net163),
    .B(net131));
 sg13g2_o21ai_1 _1432_ (.B1(_0681_),
    .Y(_0065_),
    .A1(_0141_),
    .A2(net130));
 sg13g2_nand2_1 _1433_ (.Y(_0682_),
    .A(net193),
    .B(net131));
 sg13g2_o21ai_1 _1434_ (.B1(_0682_),
    .Y(_0066_),
    .A1(_0127_),
    .A2(net130));
 sg13g2_nand2_1 _1435_ (.Y(_0683_),
    .A(net182),
    .B(net131));
 sg13g2_o21ai_1 _1436_ (.B1(_0683_),
    .Y(_0067_),
    .A1(_0128_),
    .A2(net130));
 sg13g2_nand2_1 _1437_ (.Y(_0684_),
    .A(net103),
    .B(net131));
 sg13g2_o21ai_1 _1438_ (.B1(_0684_),
    .Y(_0068_),
    .A1(_0146_),
    .A2(net130));
 sg13g2_nand2_1 _1439_ (.Y(_0685_),
    .A(net104),
    .B(net131));
 sg13g2_o21ai_1 _1440_ (.B1(_0685_),
    .Y(_0069_),
    .A1(_0124_),
    .A2(net130));
 sg13g2_nand2_1 _1441_ (.Y(_0686_),
    .A(net95),
    .B(net132));
 sg13g2_o21ai_1 _1442_ (.B1(_0686_),
    .Y(_0070_),
    .A1(_0174_),
    .A2(_0676_));
 sg13g2_dfrbpq_2 _1443_ (.RESET_B(net180),
    .D(_0010_),
    .Q(_0009_),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1444_ (.RESET_B(net180),
    .D(net91),
    .Q(\raster.tscan.state[1] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1445_ (.RESET_B(net180),
    .D(_0001_),
    .Q(\raster.tscan.state[2] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_1 _1446_ (.RESET_B(net180),
    .D(_0002_),
    .Q(\raster.tscan.state[3] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1447_ (.RESET_B(net33),
    .D(_0011_),
    .Q(\raster.tscan.left_x[0] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _1448_ (.RESET_B(net31),
    .D(net117),
    .Q(\raster.tscan.left_x[2] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1449_ (.RESET_B(net29),
    .D(net107),
    .Q(\raster.tscan.left_x[9] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _1450_ (.RESET_B(net27),
    .D(_0014_),
    .Q(\raster.tscan.right_err[0] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1451_ (.RESET_B(net26),
    .D(_0015_),
    .Q(\raster.tscan.right_err[1] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1452_ (.RESET_B(net25),
    .D(_0016_),
    .Q(\raster.tscan.right_err[2] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1453_ (.RESET_B(net24),
    .D(_0017_),
    .Q(\raster.tscan.right_err[3] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1454_ (.RESET_B(net23),
    .D(_0018_),
    .Q(\raster.tscan.right_err[4] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1455_ (.RESET_B(net22),
    .D(_0019_),
    .Q(\raster.tscan.right_err[5] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _1456_ (.RESET_B(net21),
    .D(_0020_),
    .Q(\raster.tscan.right_err[6] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1457_ (.RESET_B(net20),
    .D(_0021_),
    .Q(\raster.tscan.right_err[7] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1458_ (.RESET_B(net80),
    .D(net199),
    .Q(\raster.tscan.right_err[8] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1459_ (.RESET_B(net79),
    .D(net111),
    .Q(\raster.tscan.left_err[0] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1460_ (.RESET_B(net78),
    .D(net181),
    .Q(\raster.tscan.left_x[1] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1461_ (.RESET_B(net77),
    .D(_0025_),
    .Q(\raster.tscan.left_x[3] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1462_ (.RESET_B(net76),
    .D(net212),
    .Q(\raster.tscan.left_x[4] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1463_ (.RESET_B(net75),
    .D(_0027_),
    .Q(\raster.tscan.left_x[5] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1464_ (.RESET_B(net74),
    .D(net208),
    .Q(\raster.tscan.left_x[6] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1465_ (.RESET_B(net73),
    .D(net190),
    .Q(\raster.tscan.left_x[7] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1466_ (.RESET_B(net72),
    .D(_0030_),
    .Q(\raster.tscan.left_x[8] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_1 _1467_ (.RESET_B(net71),
    .D(net206),
    .Q(\raster.tscan.left_err[9] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _1468_ (.RESET_B(net70),
    .D(net195),
    .Q(\raster.tscan.right_x[2] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1469_ (.RESET_B(net69),
    .D(net210),
    .Q(\raster.tscan.right_x[3] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1470_ (.RESET_B(net68),
    .D(net214),
    .Q(\raster.tscan.right_x[4] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1471_ (.RESET_B(net67),
    .D(net184),
    .Q(\raster.tscan.right_x[5] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1472_ (.RESET_B(net66),
    .D(_0036_),
    .Q(\raster.tscan.right_x[6] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1473_ (.RESET_B(net65),
    .D(_0037_),
    .Q(\raster.tscan.right_x[7] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_1 _1474_ (.RESET_B(net64),
    .D(net187),
    .Q(\raster.tscan.right_x[8] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1475_ (.RESET_B(net63),
    .D(net192),
    .Q(\raster.tscan.right_err[9] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _1476_ (.RESET_B(net62),
    .D(_0040_),
    .Q(\raster.tscan.left_err[1] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _1477_ (.RESET_B(net61),
    .D(_0041_),
    .Q(\raster.tscan.left_err[2] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1478_ (.RESET_B(net60),
    .D(_0042_),
    .Q(\raster.tscan.left_err[3] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _1479_ (.RESET_B(net59),
    .D(_0043_),
    .Q(\raster.tscan.left_err[4] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _1480_ (.RESET_B(net58),
    .D(_0044_),
    .Q(\raster.tscan.left_err[5] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1481_ (.RESET_B(net57),
    .D(_0045_),
    .Q(\raster.tscan.left_err[6] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1482_ (.RESET_B(net56),
    .D(_0046_),
    .Q(\raster.tscan.left_err[7] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1483_ (.RESET_B(net55),
    .D(_0047_),
    .Q(\raster.tscan.left_err[8] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _1484_ (.RESET_B(net54),
    .D(_0048_),
    .Q(\raster.hpos[0] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _1485_ (.RESET_B(net53),
    .D(_0049_),
    .Q(\raster.hpos[1] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1486_ (.RESET_B(net52),
    .D(net120),
    .Q(\raster.hpos[2] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _1487_ (.RESET_B(net51),
    .D(_0051_),
    .Q(\raster.hpos[3] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1488_ (.RESET_B(net50),
    .D(_0052_),
    .Q(\raster.hpos[4] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _1489_ (.RESET_B(net49),
    .D(net114),
    .Q(\raster.hpos[5] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _1490_ (.RESET_B(net48),
    .D(_0054_),
    .Q(\raster.hpos[6] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1491_ (.RESET_B(net47),
    .D(_0055_),
    .Q(\raster.hpos[7] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_1 _1492_ (.RESET_B(net46),
    .D(_0056_),
    .Q(\raster.hpos[8] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1493_ (.RESET_B(net45),
    .D(_0057_),
    .Q(\raster.hpos[9] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _1494_ (.RESET_B(net44),
    .D(_0058_),
    .Q(\raster.tscan.right_x[0] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1495_ (.RESET_B(net42),
    .D(_0059_),
    .Q(\raster.tscan.right_x[1] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _1496_ (.RESET_B(net81),
    .D(net102),
    .Q(\raster.tscan.right_x[9] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _1497_ (.RESET_B(net40),
    .D(net100),
    .Q(\raster.hvsync_gen.vsync ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1498_ (.RESET_B(net38),
    .D(_0061_),
    .Q(\raster.hvsync_gen.vpos[0] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1499_ (.RESET_B(net36),
    .D(net94),
    .Q(\raster.hvsync_gen.vpos[1] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1500_ (.RESET_B(net34),
    .D(_0063_),
    .Q(\raster.hvsync_gen.vpos[2] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1501_ (.RESET_B(net30),
    .D(_0064_),
    .Q(\raster.hvsync_gen.vpos[3] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _1502_ (.RESET_B(net43),
    .D(_0065_),
    .Q(\raster.hvsync_gen.vpos[4] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1503_ (.RESET_B(net39),
    .D(_0066_),
    .Q(\raster.hvsync_gen.vpos[5] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1504_ (.RESET_B(net35),
    .D(_0067_),
    .Q(\raster.hvsync_gen.vpos[6] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _1505_ (.RESET_B(net28),
    .D(_0068_),
    .Q(\raster.hvsync_gen.vpos[7] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _1506_ (.RESET_B(net37),
    .D(net105),
    .Q(\raster.hvsync_gen.vpos[8] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _1507_ (.RESET_B(net82),
    .D(net96),
    .Q(\raster.hvsync_gen.vpos[9] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _1508_ (.RESET_B(net83),
    .D(net88),
    .Q(hsync),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _1509_ (.RESET_B(net84),
    .D(net147),
    .Q(\raster.frame_counter[0] ),
    .CLK(\raster.hvsync_gen.vsync ));
 sg13g2_dfrbpq_2 _1510_ (.RESET_B(net85),
    .D(_0005_),
    .Q(\raster.frame_counter[1] ),
    .CLK(\raster.hvsync_gen.vsync ));
 sg13g2_dfrbpq_1 _1511_ (.RESET_B(net86),
    .D(_0006_),
    .Q(\raster.frame_counter[2] ),
    .CLK(\raster.hvsync_gen.vsync ));
 sg13g2_dfrbpq_1 _1512_ (.RESET_B(net32),
    .D(_0007_),
    .Q(\raster.frame_counter[3] ),
    .CLK(\raster.hvsync_gen.vsync ));
 sg13g2_dfrbpq_2 _1513_ (.RESET_B(net41),
    .D(_0008_),
    .Q(\raster.frame_counter[4] ),
    .CLK(\raster.hvsync_gen.vsync ));
 sg13g2_tiehi _1456__21 (.L_HI(net21));
 sg13g2_tiehi _1455__22 (.L_HI(net22));
 sg13g2_tiehi _1454__23 (.L_HI(net23));
 sg13g2_tiehi _1453__24 (.L_HI(net24));
 sg13g2_tiehi _1452__25 (.L_HI(net25));
 sg13g2_tiehi _1451__26 (.L_HI(net26));
 sg13g2_tiehi _1450__27 (.L_HI(net27));
 sg13g2_tiehi _1505__28 (.L_HI(net28));
 sg13g2_tiehi _1449__29 (.L_HI(net29));
 sg13g2_tiehi _1501__30 (.L_HI(net30));
 sg13g2_tiehi _1448__31 (.L_HI(net31));
 sg13g2_tiehi _1512__32 (.L_HI(net32));
 sg13g2_tiehi _1447__33 (.L_HI(net33));
 sg13g2_tiehi _1500__34 (.L_HI(net34));
 sg13g2_tiehi _1504__35 (.L_HI(net35));
 sg13g2_tiehi _1499__36 (.L_HI(net36));
 sg13g2_tiehi _1506__37 (.L_HI(net37));
 sg13g2_tiehi _1498__38 (.L_HI(net38));
 sg13g2_tiehi _1503__39 (.L_HI(net39));
 sg13g2_tiehi _1497__40 (.L_HI(net40));
 sg13g2_tiehi _1513__41 (.L_HI(net41));
 sg13g2_tiehi _1495__42 (.L_HI(net42));
 sg13g2_tiehi _1502__43 (.L_HI(net43));
 sg13g2_tiehi _1494__44 (.L_HI(net44));
 sg13g2_tiehi _1493__45 (.L_HI(net45));
 sg13g2_tiehi _1492__46 (.L_HI(net46));
 sg13g2_tiehi _1491__47 (.L_HI(net47));
 sg13g2_tiehi _1490__48 (.L_HI(net48));
 sg13g2_tiehi _1489__49 (.L_HI(net49));
 sg13g2_tiehi _1488__50 (.L_HI(net50));
 sg13g2_tiehi _1487__51 (.L_HI(net51));
 sg13g2_tiehi _1486__52 (.L_HI(net52));
 sg13g2_tiehi _1485__53 (.L_HI(net53));
 sg13g2_tiehi _1484__54 (.L_HI(net54));
 sg13g2_tiehi _1483__55 (.L_HI(net55));
 sg13g2_tiehi _1482__56 (.L_HI(net56));
 sg13g2_tiehi _1481__57 (.L_HI(net57));
 sg13g2_tiehi _1480__58 (.L_HI(net58));
 sg13g2_tiehi _1479__59 (.L_HI(net59));
 sg13g2_tiehi _1478__60 (.L_HI(net60));
 sg13g2_tiehi _1477__61 (.L_HI(net61));
 sg13g2_tiehi _1476__62 (.L_HI(net62));
 sg13g2_tiehi _1475__63 (.L_HI(net63));
 sg13g2_tiehi _1474__64 (.L_HI(net64));
 sg13g2_tiehi _1473__65 (.L_HI(net65));
 sg13g2_tiehi _1472__66 (.L_HI(net66));
 sg13g2_tiehi _1471__67 (.L_HI(net67));
 sg13g2_tiehi _1470__68 (.L_HI(net68));
 sg13g2_tiehi _1469__69 (.L_HI(net69));
 sg13g2_tiehi _1468__70 (.L_HI(net70));
 sg13g2_tiehi _1467__71 (.L_HI(net71));
 sg13g2_tiehi _1466__72 (.L_HI(net72));
 sg13g2_tiehi _1465__73 (.L_HI(net73));
 sg13g2_tiehi _1464__74 (.L_HI(net74));
 sg13g2_tiehi _1463__75 (.L_HI(net75));
 sg13g2_tiehi _1462__76 (.L_HI(net76));
 sg13g2_tiehi _1461__77 (.L_HI(net77));
 sg13g2_tiehi _1460__78 (.L_HI(net78));
 sg13g2_tiehi _1459__79 (.L_HI(net79));
 sg13g2_tiehi _1458__80 (.L_HI(net80));
 sg13g2_tiehi _1496__81 (.L_HI(net81));
 sg13g2_tiehi _1507__82 (.L_HI(net82));
 sg13g2_tiehi _1508__83 (.L_HI(net83));
 sg13g2_tiehi _1509__84 (.L_HI(net84));
 sg13g2_tiehi _1510__85 (.L_HI(net85));
 sg13g2_tiehi _1511__86 (.L_HI(net86));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_tomolt_rasterizer_3 (.L_LO(net3));
 sg13g2_tielo tt_um_tomolt_rasterizer_4 (.L_LO(net4));
 sg13g2_tielo tt_um_tomolt_rasterizer_5 (.L_LO(net5));
 sg13g2_tielo tt_um_tomolt_rasterizer_6 (.L_LO(net6));
 sg13g2_tielo tt_um_tomolt_rasterizer_7 (.L_LO(net7));
 sg13g2_tielo tt_um_tomolt_rasterizer_8 (.L_LO(net8));
 sg13g2_tielo tt_um_tomolt_rasterizer_9 (.L_LO(net9));
 sg13g2_tielo tt_um_tomolt_rasterizer_10 (.L_LO(net10));
 sg13g2_tielo tt_um_tomolt_rasterizer_11 (.L_LO(net11));
 sg13g2_tielo tt_um_tomolt_rasterizer_12 (.L_LO(net12));
 sg13g2_tielo tt_um_tomolt_rasterizer_13 (.L_LO(net13));
 sg13g2_tielo tt_um_tomolt_rasterizer_14 (.L_LO(net14));
 sg13g2_tielo tt_um_tomolt_rasterizer_15 (.L_LO(net15));
 sg13g2_tielo tt_um_tomolt_rasterizer_16 (.L_LO(net16));
 sg13g2_tielo tt_um_tomolt_rasterizer_17 (.L_LO(net17));
 sg13g2_tielo tt_um_tomolt_rasterizer_18 (.L_LO(net18));
 sg13g2_tielo tt_um_tomolt_rasterizer_19 (.L_LO(net19));
 sg13g2_tiehi _1457__20 (.L_HI(net20));
 sg13g2_buf_1 _1599_ (.A(uo_out[4]),
    .X(uo_out[0]));
 sg13g2_buf_1 _1600_ (.A(uo_out[5]),
    .X(uo_out[1]));
 sg13g2_buf_1 _1601_ (.A(\raster.hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _1602_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout122 (.A(_0582_),
    .X(net122));
 sg13g2_buf_1 fanout123 (.A(_0582_),
    .X(net123));
 sg13g2_buf_8 fanout124 (.A(net125),
    .X(net124));
 sg13g2_buf_8 fanout125 (.A(_0276_),
    .X(net125));
 sg13g2_buf_8 fanout126 (.A(_0523_),
    .X(net126));
 sg13g2_buf_8 fanout127 (.A(_0523_),
    .X(net127));
 sg13g2_buf_8 fanout128 (.A(_0237_),
    .X(net128));
 sg13g2_buf_1 fanout129 (.A(_0237_),
    .X(net129));
 sg13g2_buf_8 fanout130 (.A(_0676_),
    .X(net130));
 sg13g2_buf_8 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(_0649_),
    .X(net132));
 sg13g2_buf_8 fanout133 (.A(net134),
    .X(net133));
 sg13g2_buf_8 fanout134 (.A(net138),
    .X(net134));
 sg13g2_buf_8 fanout135 (.A(net137),
    .X(net135));
 sg13g2_buf_1 fanout136 (.A(net137),
    .X(net136));
 sg13g2_buf_8 fanout137 (.A(net138),
    .X(net137));
 sg13g2_buf_8 fanout138 (.A(_0112_),
    .X(net138));
 sg13g2_buf_8 fanout139 (.A(net140),
    .X(net139));
 sg13g2_buf_8 fanout140 (.A(_0111_),
    .X(net140));
 sg13g2_buf_8 fanout141 (.A(net142),
    .X(net141));
 sg13g2_buf_8 fanout142 (.A(_0111_),
    .X(net142));
 sg13g2_buf_8 fanout143 (.A(net144),
    .X(net143));
 sg13g2_buf_8 fanout144 (.A(_0239_),
    .X(net144));
 sg13g2_buf_8 fanout145 (.A(_0222_),
    .X(net145));
 sg13g2_buf_1 fanout146 (.A(_0222_),
    .X(net146));
 sg13g2_buf_8 fanout147 (.A(\raster.geometry[14] ),
    .X(net147));
 sg13g2_buf_8 fanout148 (.A(\raster.geometry[14] ),
    .X(net148));
 sg13g2_buf_8 fanout149 (.A(net150),
    .X(net149));
 sg13g2_buf_8 fanout150 (.A(\raster.frame_counter[3] ),
    .X(net150));
 sg13g2_buf_8 fanout151 (.A(\raster.frame_counter[2] ),
    .X(net151));
 sg13g2_buf_8 fanout152 (.A(net154),
    .X(net152));
 sg13g2_buf_1 fanout153 (.A(net154),
    .X(net153));
 sg13g2_buf_1 fanout154 (.A(\raster.frame_counter[0] ),
    .X(net154));
 sg13g2_buf_8 fanout155 (.A(net157),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(net157),
    .X(net156));
 sg13g2_buf_1 fanout157 (.A(\raster.frame_counter[0] ),
    .X(net157));
 sg13g2_buf_8 fanout158 (.A(net159),
    .X(net158));
 sg13g2_buf_8 fanout159 (.A(net160),
    .X(net159));
 sg13g2_buf_8 fanout160 (.A(\raster.frame_counter[0] ),
    .X(net160));
 sg13g2_buf_8 fanout161 (.A(_0220_),
    .X(net161));
 sg13g2_buf_8 fanout162 (.A(_0219_),
    .X(net162));
 sg13g2_buf_8 fanout163 (.A(net232),
    .X(net163));
 sg13g2_buf_8 fanout164 (.A(net93),
    .X(net164));
 sg13g2_buf_8 fanout165 (.A(net89),
    .X(net165));
 sg13g2_buf_8 fanout166 (.A(net87),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(net236),
    .X(net167));
 sg13g2_buf_8 fanout168 (.A(net233),
    .X(net168));
 sg13g2_buf_8 fanout169 (.A(net237),
    .X(net169));
 sg13g2_buf_8 fanout170 (.A(net235),
    .X(net170));
 sg13g2_buf_8 fanout171 (.A(net115),
    .X(net171));
 sg13g2_buf_1 fanout172 (.A(\raster.tscan.state[3] ),
    .X(net172));
 sg13g2_buf_8 fanout173 (.A(net174),
    .X(net173));
 sg13g2_buf_8 fanout174 (.A(net178),
    .X(net174));
 sg13g2_buf_8 fanout175 (.A(net176),
    .X(net175));
 sg13g2_buf_8 fanout176 (.A(net177),
    .X(net176));
 sg13g2_buf_8 fanout177 (.A(net178),
    .X(net177));
 sg13g2_buf_8 fanout178 (.A(net234),
    .X(net178));
 sg13g2_buf_8 fanout179 (.A(net213),
    .X(net179));
 sg13g2_buf_8 fanout180 (.A(net1),
    .X(net180));
 sg13g2_buf_2 input1 (.A(rst_n),
    .X(net1));
 sg13g2_tielo tt_um_tomolt_rasterizer_2 (.L_LO(net2));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_2_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_4_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_4_12_0_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\raster.hpos[8] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0003_),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold3 (.A(\raster.hvsync_gen.vpos[0] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0009_),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0000_),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold6 (.A(\raster.tscan.right_x[0] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold7 (.A(\raster.hvsync_gen.vpos[1] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold8 (.A(_0062_),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold9 (.A(\raster.hvsync_gen.vpos[9] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0070_),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold11 (.A(\raster.tscan.right_err[0] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0281_),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold13 (.A(\raster.hvsync_gen.vpos[2] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0004_),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold15 (.A(\raster.tscan.right_x[9] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0060_),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold17 (.A(\raster.hvsync_gen.vpos[7] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold18 (.A(\raster.hvsync_gen.vpos[8] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0069_),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold20 (.A(\raster.tscan.left_x[9] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0013_),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold22 (.A(\raster.tscan.right_x[1] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold23 (.A(\raster.tscan.left_err[0] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold24 (.A(_0428_),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0023_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold26 (.A(\raster.hpos[5] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold27 (.A(_0655_),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0053_),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold29 (.A(\raster.tscan.state[3] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold30 (.A(\raster.tscan.left_x[2] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0012_),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold32 (.A(\raster.hpos[2] ),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold33 (.A(_0652_),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0050_),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold35 (.A(\raster.tscan.left_x[1] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0024_),
    .X(net181));
 sg13g2_dlygate4sd3_1 hold37 (.A(\raster.hvsync_gen.vpos[6] ),
    .X(net182));
 sg13g2_dlygate4sd3_1 hold38 (.A(\raster.tscan.right_x[5] ),
    .X(net183));
 sg13g2_dlygate4sd3_1 hold39 (.A(_0035_),
    .X(net184));
 sg13g2_dlygate4sd3_1 hold40 (.A(\raster.hpos[0] ),
    .X(net185));
 sg13g2_dlygate4sd3_1 hold41 (.A(\raster.tscan.right_x[8] ),
    .X(net186));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0038_),
    .X(net187));
 sg13g2_dlygate4sd3_1 hold43 (.A(\raster.hvsync_gen.vpos[3] ),
    .X(net188));
 sg13g2_dlygate4sd3_1 hold44 (.A(\raster.tscan.left_x[7] ),
    .X(net189));
 sg13g2_dlygate4sd3_1 hold45 (.A(_0029_),
    .X(net190));
 sg13g2_dlygate4sd3_1 hold46 (.A(\raster.tscan.right_err[9] ),
    .X(net191));
 sg13g2_dlygate4sd3_1 hold47 (.A(_0039_),
    .X(net192));
 sg13g2_dlygate4sd3_1 hold48 (.A(\raster.hvsync_gen.vpos[5] ),
    .X(net193));
 sg13g2_dlygate4sd3_1 hold49 (.A(\raster.tscan.right_x[2] ),
    .X(net194));
 sg13g2_dlygate4sd3_1 hold50 (.A(_0032_),
    .X(net195));
 sg13g2_dlygate4sd3_1 hold51 (.A(\raster.tscan.right_err[6] ),
    .X(net196));
 sg13g2_dlygate4sd3_1 hold52 (.A(\raster.tscan.left_err[7] ),
    .X(net197));
 sg13g2_dlygate4sd3_1 hold53 (.A(\raster.tscan.right_err[8] ),
    .X(net198));
 sg13g2_dlygate4sd3_1 hold54 (.A(_0022_),
    .X(net199));
 sg13g2_dlygate4sd3_1 hold55 (.A(\raster.tscan.left_x[5] ),
    .X(net200));
 sg13g2_dlygate4sd3_1 hold56 (.A(_0444_),
    .X(net201));
 sg13g2_dlygate4sd3_1 hold57 (.A(\raster.tscan.left_err[8] ),
    .X(net202));
 sg13g2_dlygate4sd3_1 hold58 (.A(\raster.tscan.right_x[6] ),
    .X(net203));
 sg13g2_dlygate4sd3_1 hold59 (.A(\raster.tscan.right_err[5] ),
    .X(net204));
 sg13g2_dlygate4sd3_1 hold60 (.A(\raster.tscan.left_err[9] ),
    .X(net205));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0031_),
    .X(net206));
 sg13g2_dlygate4sd3_1 hold62 (.A(\raster.tscan.left_x[6] ),
    .X(net207));
 sg13g2_dlygate4sd3_1 hold63 (.A(_0028_),
    .X(net208));
 sg13g2_dlygate4sd3_1 hold64 (.A(\raster.tscan.right_x[3] ),
    .X(net209));
 sg13g2_dlygate4sd3_1 hold65 (.A(_0033_),
    .X(net210));
 sg13g2_dlygate4sd3_1 hold66 (.A(\raster.tscan.left_x[4] ),
    .X(net211));
 sg13g2_dlygate4sd3_1 hold67 (.A(_0026_),
    .X(net212));
 sg13g2_dlygate4sd3_1 hold68 (.A(\raster.tscan.state[1] ),
    .X(net213));
 sg13g2_dlygate4sd3_1 hold69 (.A(_0034_),
    .X(net214));
 sg13g2_dlygate4sd3_1 hold70 (.A(\raster.tscan.left_x[3] ),
    .X(net215));
 sg13g2_dlygate4sd3_1 hold71 (.A(\raster.tscan.right_err[4] ),
    .X(net216));
 sg13g2_dlygate4sd3_1 hold72 (.A(\raster.tscan.left_x[8] ),
    .X(net217));
 sg13g2_dlygate4sd3_1 hold73 (.A(\raster.tscan.right_err[1] ),
    .X(net218));
 sg13g2_dlygate4sd3_1 hold74 (.A(\raster.hpos[1] ),
    .X(net219));
 sg13g2_dlygate4sd3_1 hold75 (.A(\raster.tscan.left_err[2] ),
    .X(net220));
 sg13g2_dlygate4sd3_1 hold76 (.A(\raster.tscan.left_err[4] ),
    .X(net221));
 sg13g2_dlygate4sd3_1 hold77 (.A(\raster.tscan.left_err[3] ),
    .X(net222));
 sg13g2_dlygate4sd3_1 hold78 (.A(\raster.hpos[3] ),
    .X(net223));
 sg13g2_dlygate4sd3_1 hold79 (.A(\raster.hpos[7] ),
    .X(net224));
 sg13g2_dlygate4sd3_1 hold80 (.A(_0660_),
    .X(net225));
 sg13g2_dlygate4sd3_1 hold81 (.A(\raster.tscan.left_err[6] ),
    .X(net226));
 sg13g2_dlygate4sd3_1 hold82 (.A(\raster.tscan.right_x[7] ),
    .X(net227));
 sg13g2_dlygate4sd3_1 hold83 (.A(\raster.tscan.left_err[1] ),
    .X(net228));
 sg13g2_dlygate4sd3_1 hold84 (.A(\raster.tscan.left_x[0] ),
    .X(net229));
 sg13g2_dlygate4sd3_1 hold85 (.A(\raster.hpos[9] ),
    .X(net230));
 sg13g2_dlygate4sd3_1 hold86 (.A(\raster.hpos[4] ),
    .X(net231));
 sg13g2_dlygate4sd3_1 hold87 (.A(\raster.hvsync_gen.vpos[4] ),
    .X(net232));
 sg13g2_dlygate4sd3_1 hold88 (.A(\raster.tscan.left_err[5] ),
    .X(net233));
 sg13g2_dlygate4sd3_1 hold89 (.A(\raster.tscan.state[2] ),
    .X(net234));
 sg13g2_dlygate4sd3_1 hold90 (.A(\raster.tscan.right_err[2] ),
    .X(net235));
 sg13g2_dlygate4sd3_1 hold91 (.A(\raster.hpos[6] ),
    .X(net236));
 sg13g2_dlygate4sd3_1 hold92 (.A(\raster.tscan.right_err[3] ),
    .X(net237));
 sg13g2_dlygate4sd3_1 hold93 (.A(\raster.tscan.right_err[7] ),
    .X(net238));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_67 ();
 sg13g2_decap_8 FILLER_7_74 ();
 sg13g2_decap_8 FILLER_7_90 ();
 sg13g2_decap_8 FILLER_7_97 ();
 sg13g2_decap_8 FILLER_7_104 ();
 sg13g2_decap_8 FILLER_7_111 ();
 sg13g2_decap_8 FILLER_7_118 ();
 sg13g2_decap_8 FILLER_7_125 ();
 sg13g2_decap_4 FILLER_7_132 ();
 sg13g2_fill_2 FILLER_7_136 ();
 sg13g2_fill_2 FILLER_7_142 ();
 sg13g2_decap_8 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_160 ();
 sg13g2_fill_2 FILLER_7_167 ();
 sg13g2_fill_1 FILLER_7_169 ();
 sg13g2_decap_8 FILLER_7_198 ();
 sg13g2_decap_4 FILLER_7_205 ();
 sg13g2_fill_2 FILLER_7_209 ();
 sg13g2_decap_8 FILLER_7_220 ();
 sg13g2_decap_8 FILLER_7_227 ();
 sg13g2_decap_8 FILLER_7_234 ();
 sg13g2_decap_8 FILLER_7_241 ();
 sg13g2_decap_8 FILLER_7_248 ();
 sg13g2_decap_8 FILLER_7_255 ();
 sg13g2_decap_8 FILLER_7_262 ();
 sg13g2_decap_8 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_276 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_fill_1 FILLER_8_56 ();
 sg13g2_fill_1 FILLER_8_85 ();
 sg13g2_decap_4 FILLER_8_103 ();
 sg13g2_fill_2 FILLER_8_120 ();
 sg13g2_fill_1 FILLER_8_122 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_fill_2 FILLER_8_173 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_229 ();
 sg13g2_decap_4 FILLER_8_236 ();
 sg13g2_fill_2 FILLER_8_240 ();
 sg13g2_decap_8 FILLER_8_246 ();
 sg13g2_fill_2 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_4 FILLER_8_403 ();
 sg13g2_fill_2 FILLER_8_407 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_4 FILLER_9_63 ();
 sg13g2_fill_2 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_fill_2 FILLER_9_81 ();
 sg13g2_fill_1 FILLER_9_83 ();
 sg13g2_decap_4 FILLER_9_105 ();
 sg13g2_fill_2 FILLER_9_122 ();
 sg13g2_fill_1 FILLER_9_124 ();
 sg13g2_fill_2 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_4 FILLER_9_154 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_fill_1 FILLER_9_169 ();
 sg13g2_fill_1 FILLER_9_180 ();
 sg13g2_fill_2 FILLER_9_191 ();
 sg13g2_decap_4 FILLER_9_216 ();
 sg13g2_fill_1 FILLER_9_220 ();
 sg13g2_decap_8 FILLER_9_225 ();
 sg13g2_decap_4 FILLER_9_232 ();
 sg13g2_fill_1 FILLER_9_236 ();
 sg13g2_fill_2 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_267 ();
 sg13g2_decap_8 FILLER_9_272 ();
 sg13g2_decap_8 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_286 ();
 sg13g2_decap_8 FILLER_9_293 ();
 sg13g2_decap_8 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_4 FILLER_10_28 ();
 sg13g2_fill_2 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_87 ();
 sg13g2_decap_4 FILLER_10_98 ();
 sg13g2_decap_4 FILLER_10_106 ();
 sg13g2_fill_2 FILLER_10_110 ();
 sg13g2_decap_8 FILLER_10_117 ();
 sg13g2_decap_4 FILLER_10_124 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_fill_1 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_174 ();
 sg13g2_decap_8 FILLER_10_181 ();
 sg13g2_fill_1 FILLER_10_188 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_4 FILLER_10_212 ();
 sg13g2_decap_4 FILLER_10_244 ();
 sg13g2_fill_1 FILLER_10_248 ();
 sg13g2_fill_1 FILLER_10_262 ();
 sg13g2_decap_4 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_330 ();
 sg13g2_decap_8 FILLER_10_337 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_358 ();
 sg13g2_decap_8 FILLER_10_365 ();
 sg13g2_decap_8 FILLER_10_372 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_8 FILLER_10_393 ();
 sg13g2_decap_8 FILLER_10_400 ();
 sg13g2_fill_2 FILLER_10_407 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_41 ();
 sg13g2_decap_8 FILLER_11_48 ();
 sg13g2_decap_8 FILLER_11_79 ();
 sg13g2_decap_4 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_decap_4 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_147 ();
 sg13g2_fill_2 FILLER_11_153 ();
 sg13g2_fill_1 FILLER_11_155 ();
 sg13g2_decap_4 FILLER_11_178 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_fill_2 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_267 ();
 sg13g2_fill_2 FILLER_11_274 ();
 sg13g2_decap_4 FILLER_11_295 ();
 sg13g2_fill_1 FILLER_11_299 ();
 sg13g2_fill_1 FILLER_11_304 ();
 sg13g2_decap_4 FILLER_11_314 ();
 sg13g2_fill_2 FILLER_11_318 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_32 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_103 ();
 sg13g2_decap_8 FILLER_12_122 ();
 sg13g2_decap_4 FILLER_12_129 ();
 sg13g2_fill_1 FILLER_12_133 ();
 sg13g2_decap_4 FILLER_12_143 ();
 sg13g2_fill_1 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_fill_2 FILLER_12_161 ();
 sg13g2_fill_1 FILLER_12_163 ();
 sg13g2_decap_4 FILLER_12_173 ();
 sg13g2_fill_2 FILLER_12_177 ();
 sg13g2_decap_8 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_236 ();
 sg13g2_decap_4 FILLER_12_243 ();
 sg13g2_decap_8 FILLER_12_260 ();
 sg13g2_decap_4 FILLER_12_267 ();
 sg13g2_fill_2 FILLER_12_271 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_decap_4 FILLER_12_330 ();
 sg13g2_fill_2 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_4 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_376 ();
 sg13g2_decap_8 FILLER_12_383 ();
 sg13g2_decap_8 FILLER_12_390 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_4 FILLER_12_404 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_37 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_128 ();
 sg13g2_fill_2 FILLER_13_156 ();
 sg13g2_decap_4 FILLER_13_163 ();
 sg13g2_fill_2 FILLER_13_167 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_fill_1 FILLER_13_189 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_fill_1 FILLER_13_224 ();
 sg13g2_fill_1 FILLER_13_234 ();
 sg13g2_decap_4 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_274 ();
 sg13g2_decap_4 FILLER_13_299 ();
 sg13g2_fill_1 FILLER_13_303 ();
 sg13g2_fill_1 FILLER_13_314 ();
 sg13g2_decap_4 FILLER_13_353 ();
 sg13g2_decap_8 FILLER_13_395 ();
 sg13g2_decap_8 FILLER_13_402 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_38 ();
 sg13g2_decap_8 FILLER_14_45 ();
 sg13g2_decap_4 FILLER_14_52 ();
 sg13g2_fill_1 FILLER_14_56 ();
 sg13g2_fill_2 FILLER_14_81 ();
 sg13g2_fill_1 FILLER_14_83 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_fill_2 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_121 ();
 sg13g2_decap_8 FILLER_14_128 ();
 sg13g2_decap_8 FILLER_14_135 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_decap_8 FILLER_14_149 ();
 sg13g2_fill_2 FILLER_14_156 ();
 sg13g2_fill_1 FILLER_14_158 ();
 sg13g2_fill_2 FILLER_14_197 ();
 sg13g2_fill_2 FILLER_14_205 ();
 sg13g2_decap_4 FILLER_14_212 ();
 sg13g2_fill_2 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_decap_4 FILLER_14_248 ();
 sg13g2_fill_2 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_272 ();
 sg13g2_decap_4 FILLER_14_290 ();
 sg13g2_fill_2 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_4 FILLER_14_331 ();
 sg13g2_fill_2 FILLER_14_335 ();
 sg13g2_decap_4 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_357 ();
 sg13g2_decap_4 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_4 FILLER_15_69 ();
 sg13g2_decap_4 FILLER_15_98 ();
 sg13g2_decap_4 FILLER_15_118 ();
 sg13g2_fill_2 FILLER_15_135 ();
 sg13g2_fill_1 FILLER_15_137 ();
 sg13g2_decap_4 FILLER_15_143 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_175 ();
 sg13g2_fill_1 FILLER_15_191 ();
 sg13g2_fill_2 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_209 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_4 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_235 ();
 sg13g2_fill_2 FILLER_15_241 ();
 sg13g2_fill_2 FILLER_15_248 ();
 sg13g2_decap_4 FILLER_15_271 ();
 sg13g2_fill_1 FILLER_15_275 ();
 sg13g2_decap_4 FILLER_15_301 ();
 sg13g2_fill_2 FILLER_15_305 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_fill_2 FILLER_15_348 ();
 sg13g2_fill_1 FILLER_15_350 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_fill_1 FILLER_15_372 ();
 sg13g2_decap_8 FILLER_15_394 ();
 sg13g2_decap_8 FILLER_15_401 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_4 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_43 ();
 sg13g2_decap_4 FILLER_16_50 ();
 sg13g2_fill_2 FILLER_16_54 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_84 ();
 sg13g2_decap_4 FILLER_16_101 ();
 sg13g2_fill_2 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_120 ();
 sg13g2_fill_2 FILLER_16_127 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_161 ();
 sg13g2_fill_2 FILLER_16_189 ();
 sg13g2_fill_1 FILLER_16_210 ();
 sg13g2_decap_4 FILLER_16_228 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_fill_2 FILLER_16_255 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_decap_8 FILLER_16_267 ();
 sg13g2_decap_8 FILLER_16_274 ();
 sg13g2_decap_4 FILLER_16_281 ();
 sg13g2_fill_1 FILLER_16_285 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_fill_1 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_313 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_decap_4 FILLER_16_327 ();
 sg13g2_fill_2 FILLER_16_331 ();
 sg13g2_decap_4 FILLER_16_352 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_decap_4 FILLER_16_372 ();
 sg13g2_fill_2 FILLER_16_376 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_4 FILLER_17_28 ();
 sg13g2_fill_2 FILLER_17_32 ();
 sg13g2_fill_2 FILLER_17_62 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_decap_8 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_85 ();
 sg13g2_decap_4 FILLER_17_103 ();
 sg13g2_fill_1 FILLER_17_107 ();
 sg13g2_decap_4 FILLER_17_123 ();
 sg13g2_fill_1 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_197 ();
 sg13g2_decap_8 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_211 ();
 sg13g2_decap_8 FILLER_17_222 ();
 sg13g2_fill_1 FILLER_17_229 ();
 sg13g2_decap_8 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_261 ();
 sg13g2_fill_1 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_275 ();
 sg13g2_fill_2 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_295 ();
 sg13g2_decap_4 FILLER_17_311 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_fill_2 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_373 ();
 sg13g2_fill_1 FILLER_17_380 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_4 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_111 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_decap_4 FILLER_18_119 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_decap_8 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_165 ();
 sg13g2_fill_1 FILLER_18_167 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_decap_8 FILLER_18_248 ();
 sg13g2_fill_1 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_275 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_fill_2 FILLER_18_348 ();
 sg13g2_fill_1 FILLER_18_350 ();
 sg13g2_fill_2 FILLER_18_356 ();
 sg13g2_fill_1 FILLER_18_358 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_fill_1 FILLER_18_375 ();
 sg13g2_decap_4 FILLER_18_381 ();
 sg13g2_fill_2 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_391 ();
 sg13g2_decap_8 FILLER_18_398 ();
 sg13g2_decap_4 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_4 FILLER_19_42 ();
 sg13g2_fill_2 FILLER_19_46 ();
 sg13g2_decap_4 FILLER_19_76 ();
 sg13g2_fill_1 FILLER_19_80 ();
 sg13g2_decap_4 FILLER_19_142 ();
 sg13g2_fill_2 FILLER_19_146 ();
 sg13g2_fill_1 FILLER_19_175 ();
 sg13g2_decap_4 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_251 ();
 sg13g2_fill_2 FILLER_19_258 ();
 sg13g2_fill_1 FILLER_19_260 ();
 sg13g2_decap_4 FILLER_19_272 ();
 sg13g2_decap_4 FILLER_19_317 ();
 sg13g2_fill_1 FILLER_19_321 ();
 sg13g2_fill_2 FILLER_19_365 ();
 sg13g2_decap_4 FILLER_19_388 ();
 sg13g2_fill_1 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_402 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_4 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_57 ();
 sg13g2_decap_4 FILLER_20_64 ();
 sg13g2_fill_2 FILLER_20_68 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_fill_2 FILLER_20_81 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_4 FILLER_20_147 ();
 sg13g2_fill_2 FILLER_20_151 ();
 sg13g2_decap_4 FILLER_20_157 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_fill_2 FILLER_20_172 ();
 sg13g2_fill_1 FILLER_20_174 ();
 sg13g2_decap_8 FILLER_20_192 ();
 sg13g2_decap_4 FILLER_20_199 ();
 sg13g2_decap_4 FILLER_20_209 ();
 sg13g2_fill_2 FILLER_20_213 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_4 FILLER_20_231 ();
 sg13g2_fill_1 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_240 ();
 sg13g2_fill_2 FILLER_20_247 ();
 sg13g2_decap_4 FILLER_20_259 ();
 sg13g2_fill_1 FILLER_20_263 ();
 sg13g2_fill_2 FILLER_20_276 ();
 sg13g2_decap_4 FILLER_20_310 ();
 sg13g2_fill_1 FILLER_20_314 ();
 sg13g2_fill_1 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_fill_1 FILLER_20_375 ();
 sg13g2_fill_1 FILLER_20_380 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_fill_2 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_44 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_4 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_100 ();
 sg13g2_decap_8 FILLER_21_143 ();
 sg13g2_decap_4 FILLER_21_150 ();
 sg13g2_fill_2 FILLER_21_154 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_decap_4 FILLER_21_192 ();
 sg13g2_decap_4 FILLER_21_204 ();
 sg13g2_fill_2 FILLER_21_259 ();
 sg13g2_fill_1 FILLER_21_261 ();
 sg13g2_fill_2 FILLER_21_276 ();
 sg13g2_fill_1 FILLER_21_278 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_decap_8 FILLER_21_398 ();
 sg13g2_decap_4 FILLER_21_405 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_fill_2 FILLER_22_86 ();
 sg13g2_decap_4 FILLER_22_92 ();
 sg13g2_fill_2 FILLER_22_96 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_decap_4 FILLER_22_110 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_decap_4 FILLER_22_151 ();
 sg13g2_decap_4 FILLER_22_181 ();
 sg13g2_decap_8 FILLER_22_198 ();
 sg13g2_fill_1 FILLER_22_205 ();
 sg13g2_decap_4 FILLER_22_214 ();
 sg13g2_fill_1 FILLER_22_218 ();
 sg13g2_fill_2 FILLER_22_241 ();
 sg13g2_fill_2 FILLER_22_252 ();
 sg13g2_fill_1 FILLER_22_277 ();
 sg13g2_decap_4 FILLER_22_282 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_372 ();
 sg13g2_decap_8 FILLER_22_379 ();
 sg13g2_fill_1 FILLER_22_386 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_49 ();
 sg13g2_fill_2 FILLER_23_53 ();
 sg13g2_fill_2 FILLER_23_111 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_decap_8 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_157 ();
 sg13g2_fill_1 FILLER_23_164 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_fill_2 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_178 ();
 sg13g2_fill_1 FILLER_23_213 ();
 sg13g2_fill_1 FILLER_23_252 ();
 sg13g2_decap_4 FILLER_23_279 ();
 sg13g2_fill_1 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_301 ();
 sg13g2_fill_2 FILLER_23_309 ();
 sg13g2_fill_1 FILLER_23_339 ();
 sg13g2_fill_2 FILLER_23_353 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_377 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_4 FILLER_24_35 ();
 sg13g2_fill_2 FILLER_24_39 ();
 sg13g2_fill_1 FILLER_24_69 ();
 sg13g2_fill_2 FILLER_24_97 ();
 sg13g2_fill_1 FILLER_24_99 ();
 sg13g2_fill_2 FILLER_24_104 ();
 sg13g2_decap_8 FILLER_24_115 ();
 sg13g2_decap_8 FILLER_24_122 ();
 sg13g2_decap_8 FILLER_24_134 ();
 sg13g2_decap_8 FILLER_24_141 ();
 sg13g2_decap_4 FILLER_24_148 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_fill_2 FILLER_24_178 ();
 sg13g2_fill_1 FILLER_24_180 ();
 sg13g2_decap_4 FILLER_24_187 ();
 sg13g2_fill_2 FILLER_24_191 ();
 sg13g2_fill_1 FILLER_24_200 ();
 sg13g2_decap_4 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_266 ();
 sg13g2_decap_8 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_fill_1 FILLER_24_301 ();
 sg13g2_fill_1 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_311 ();
 sg13g2_decap_8 FILLER_24_318 ();
 sg13g2_fill_2 FILLER_24_348 ();
 sg13g2_fill_1 FILLER_24_350 ();
 sg13g2_fill_2 FILLER_24_382 ();
 sg13g2_fill_1 FILLER_24_398 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_4 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_50 ();
 sg13g2_decap_4 FILLER_25_55 ();
 sg13g2_fill_2 FILLER_25_59 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_fill_2 FILLER_25_96 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_fill_2 FILLER_25_118 ();
 sg13g2_fill_2 FILLER_25_126 ();
 sg13g2_fill_1 FILLER_25_128 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_4 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_272 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_fill_2 FILLER_25_282 ();
 sg13g2_fill_1 FILLER_25_296 ();
 sg13g2_decap_4 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_329 ();
 sg13g2_decap_4 FILLER_25_334 ();
 sg13g2_decap_4 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_4 FILLER_26_42 ();
 sg13g2_fill_2 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_76 ();
 sg13g2_fill_1 FILLER_26_96 ();
 sg13g2_decap_4 FILLER_26_132 ();
 sg13g2_fill_1 FILLER_26_136 ();
 sg13g2_decap_4 FILLER_26_148 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_4 FILLER_26_174 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_187 ();
 sg13g2_decap_8 FILLER_26_194 ();
 sg13g2_fill_1 FILLER_26_201 ();
 sg13g2_decap_4 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_215 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_2 FILLER_26_264 ();
 sg13g2_decap_4 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_351 ();
 sg13g2_decap_4 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_fill_2 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_4 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_53 ();
 sg13g2_decap_8 FILLER_27_58 ();
 sg13g2_decap_4 FILLER_27_65 ();
 sg13g2_fill_1 FILLER_27_95 ();
 sg13g2_fill_1 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_151 ();
 sg13g2_fill_1 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_fill_1 FILLER_27_192 ();
 sg13g2_decap_4 FILLER_27_217 ();
 sg13g2_decap_4 FILLER_27_225 ();
 sg13g2_fill_2 FILLER_27_229 ();
 sg13g2_decap_4 FILLER_27_244 ();
 sg13g2_fill_1 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_fill_2 FILLER_27_270 ();
 sg13g2_fill_1 FILLER_27_280 ();
 sg13g2_fill_2 FILLER_27_302 ();
 sg13g2_fill_2 FILLER_27_344 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_fill_1 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_fill_1 FILLER_27_391 ();
 sg13g2_decap_8 FILLER_27_398 ();
 sg13g2_decap_4 FILLER_27_405 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_4 FILLER_28_42 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_decap_4 FILLER_28_75 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_96 ();
 sg13g2_fill_2 FILLER_28_108 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_decap_4 FILLER_28_121 ();
 sg13g2_fill_1 FILLER_28_125 ();
 sg13g2_fill_2 FILLER_28_131 ();
 sg13g2_fill_1 FILLER_28_133 ();
 sg13g2_fill_2 FILLER_28_146 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_fill_2 FILLER_28_190 ();
 sg13g2_decap_4 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_200 ();
 sg13g2_fill_2 FILLER_28_217 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_decap_8 FILLER_28_262 ();
 sg13g2_decap_4 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_decap_4 FILLER_28_375 ();
 sg13g2_fill_2 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_62 ();
 sg13g2_decap_8 FILLER_29_69 ();
 sg13g2_fill_1 FILLER_29_90 ();
 sg13g2_decap_8 FILLER_29_120 ();
 sg13g2_fill_2 FILLER_29_139 ();
 sg13g2_fill_1 FILLER_29_141 ();
 sg13g2_fill_1 FILLER_29_169 ();
 sg13g2_fill_1 FILLER_29_224 ();
 sg13g2_fill_1 FILLER_29_259 ();
 sg13g2_decap_4 FILLER_29_268 ();
 sg13g2_fill_2 FILLER_29_272 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_fill_2 FILLER_29_289 ();
 sg13g2_fill_1 FILLER_29_291 ();
 sg13g2_fill_2 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_303 ();
 sg13g2_fill_1 FILLER_29_331 ();
 sg13g2_decap_4 FILLER_29_356 ();
 sg13g2_fill_1 FILLER_29_360 ();
 sg13g2_fill_2 FILLER_29_366 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_fill_1 FILLER_29_380 ();
 sg13g2_decap_8 FILLER_29_400 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_4 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_108 ();
 sg13g2_decap_8 FILLER_30_115 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_fill_2 FILLER_30_140 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_fill_1 FILLER_30_156 ();
 sg13g2_fill_2 FILLER_30_166 ();
 sg13g2_fill_2 FILLER_30_198 ();
 sg13g2_decap_4 FILLER_30_217 ();
 sg13g2_fill_2 FILLER_30_221 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_decap_4 FILLER_30_261 ();
 sg13g2_fill_2 FILLER_30_265 ();
 sg13g2_fill_2 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_339 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_fill_2 FILLER_31_127 ();
 sg13g2_fill_2 FILLER_31_166 ();
 sg13g2_fill_1 FILLER_31_188 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_4 FILLER_31_245 ();
 sg13g2_fill_1 FILLER_31_249 ();
 sg13g2_fill_2 FILLER_31_263 ();
 sg13g2_decap_8 FILLER_31_268 ();
 sg13g2_fill_2 FILLER_31_275 ();
 sg13g2_fill_1 FILLER_31_277 ();
 sg13g2_decap_4 FILLER_31_282 ();
 sg13g2_fill_2 FILLER_31_286 ();
 sg13g2_decap_8 FILLER_31_296 ();
 sg13g2_decap_4 FILLER_31_303 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_316 ();
 sg13g2_fill_2 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_333 ();
 sg13g2_decap_4 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_350 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_390 ();
 sg13g2_decap_4 FILLER_31_404 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_fill_1 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_86 ();
 sg13g2_decap_8 FILLER_32_93 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_151 ();
 sg13g2_decap_4 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_decap_4 FILLER_32_203 ();
 sg13g2_fill_1 FILLER_32_207 ();
 sg13g2_fill_1 FILLER_32_212 ();
 sg13g2_fill_2 FILLER_32_223 ();
 sg13g2_fill_2 FILLER_32_241 ();
 sg13g2_decap_8 FILLER_32_258 ();
 sg13g2_decap_4 FILLER_32_265 ();
 sg13g2_fill_2 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_319 ();
 sg13g2_fill_1 FILLER_32_341 ();
 sg13g2_fill_2 FILLER_32_364 ();
 sg13g2_fill_1 FILLER_32_366 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_135 ();
 sg13g2_fill_1 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_fill_2 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_231 ();
 sg13g2_fill_1 FILLER_33_235 ();
 sg13g2_fill_2 FILLER_33_249 ();
 sg13g2_decap_4 FILLER_33_254 ();
 sg13g2_fill_2 FILLER_33_258 ();
 sg13g2_decap_4 FILLER_33_302 ();
 sg13g2_fill_2 FILLER_33_313 ();
 sg13g2_decap_4 FILLER_33_320 ();
 sg13g2_decap_8 FILLER_33_340 ();
 sg13g2_fill_2 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_349 ();
 sg13g2_fill_2 FILLER_33_380 ();
 sg13g2_fill_1 FILLER_33_382 ();
 sg13g2_fill_1 FILLER_33_396 ();
 sg13g2_fill_2 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_112 ();
 sg13g2_fill_1 FILLER_34_144 ();
 sg13g2_decap_4 FILLER_34_182 ();
 sg13g2_fill_1 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_decap_8 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_243 ();
 sg13g2_decap_4 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_258 ();
 sg13g2_fill_2 FILLER_34_262 ();
 sg13g2_decap_8 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_284 ();
 sg13g2_fill_2 FILLER_34_298 ();
 sg13g2_fill_1 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_310 ();
 sg13g2_decap_4 FILLER_34_316 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_fill_2 FILLER_34_349 ();
 sg13g2_fill_1 FILLER_34_351 ();
 sg13g2_fill_2 FILLER_34_365 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_125 ();
 sg13g2_decap_8 FILLER_35_141 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_decap_8 FILLER_35_152 ();
 sg13g2_decap_8 FILLER_35_159 ();
 sg13g2_fill_2 FILLER_35_166 ();
 sg13g2_fill_1 FILLER_35_172 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_decap_4 FILLER_35_206 ();
 sg13g2_fill_1 FILLER_35_210 ();
 sg13g2_fill_1 FILLER_35_227 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_322 ();
 sg13g2_fill_1 FILLER_35_324 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_fill_2 FILLER_36_154 ();
 sg13g2_decap_4 FILLER_36_178 ();
 sg13g2_decap_8 FILLER_36_191 ();
 sg13g2_decap_4 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_36_202 ();
 sg13g2_decap_8 FILLER_36_233 ();
 sg13g2_fill_2 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_255 ();
 sg13g2_fill_1 FILLER_36_261 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_2 FILLER_36_314 ();
 sg13g2_fill_1 FILLER_36_316 ();
 sg13g2_fill_2 FILLER_36_324 ();
 sg13g2_fill_1 FILLER_36_326 ();
 sg13g2_fill_1 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_fill_1 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_405 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_4 FILLER_37_147 ();
 sg13g2_fill_2 FILLER_37_151 ();
 sg13g2_fill_2 FILLER_37_190 ();
 sg13g2_decap_4 FILLER_37_196 ();
 sg13g2_fill_2 FILLER_37_200 ();
 sg13g2_decap_4 FILLER_37_232 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_280 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_2 FILLER_37_360 ();
 sg13g2_fill_1 FILLER_37_362 ();
 sg13g2_decap_4 FILLER_37_367 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_4 FILLER_37_403 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_decap_4 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_fill_2 FILLER_38_172 ();
 sg13g2_fill_1 FILLER_38_174 ();
 sg13g2_fill_2 FILLER_38_206 ();
 sg13g2_fill_1 FILLER_38_208 ();
 sg13g2_fill_2 FILLER_38_272 ();
 sg13g2_fill_1 FILLER_38_274 ();
 sg13g2_fill_2 FILLER_38_307 ();
 sg13g2_fill_1 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_386 ();
 sg13g2_decap_8 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_407 ();
 assign uio_oe[0] = net2;
 assign uio_oe[1] = net3;
 assign uio_oe[2] = net4;
 assign uio_oe[3] = net5;
 assign uio_oe[4] = net6;
 assign uio_oe[5] = net7;
 assign uio_oe[6] = net8;
 assign uio_oe[7] = net9;
 assign uio_out[0] = net10;
 assign uio_out[1] = net11;
 assign uio_out[2] = net12;
 assign uio_out[3] = net13;
 assign uio_out[4] = net14;
 assign uio_out[5] = net15;
 assign uio_out[6] = net16;
 assign uio_out[7] = net17;
 assign uo_out[2] = net18;
 assign uo_out[6] = net19;
endmodule
