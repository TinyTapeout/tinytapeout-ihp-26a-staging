module tt_um_wedgetail_tester (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire clk_regs;
 wire \dpll.clk8x_fout ;
 wire \dpll.clk_fout ;
 wire \dpll.id_decrement ;
 wire \dpll.id_decrement_done ;
 wire \dpll.id_increment ;
 wire \dpll.id_increment_done ;
 wire \dpll.id_out ;
 wire \dpll.k_count[0] ;
 wire \dpll.k_count[1] ;
 wire \dpll.k_count[2] ;
 wire \dpll.k_count[3] ;
 wire \dpll.k_count[4] ;
 wire \dpll.k_count[5] ;
 wire \dpll.k_count[6] ;
 wire \dpll.k_count[7] ;
 wire \dpll.k_count_borrow ;
 wire \dpll.k_count_carry ;
 wire \dpll.n_count[0] ;
 wire \dpll.n_count[1] ;
 wire \dpll.n_count[2] ;
 wire \dpll.n_count[4] ;
 wire \dpll.n_count[5] ;
 wire \mod_ro_128.fabric[0] ;
 wire \mod_ro_128.fabric[100] ;
 wire \mod_ro_128.fabric[101] ;
 wire \mod_ro_128.fabric[102] ;
 wire \mod_ro_128.fabric[103] ;
 wire \mod_ro_128.fabric[104] ;
 wire \mod_ro_128.fabric[105] ;
 wire \mod_ro_128.fabric[106] ;
 wire \mod_ro_128.fabric[107] ;
 wire \mod_ro_128.fabric[108] ;
 wire \mod_ro_128.fabric[109] ;
 wire \mod_ro_128.fabric[10] ;
 wire \mod_ro_128.fabric[110] ;
 wire \mod_ro_128.fabric[111] ;
 wire \mod_ro_128.fabric[112] ;
 wire \mod_ro_128.fabric[113] ;
 wire \mod_ro_128.fabric[114] ;
 wire \mod_ro_128.fabric[115] ;
 wire \mod_ro_128.fabric[116] ;
 wire \mod_ro_128.fabric[117] ;
 wire \mod_ro_128.fabric[118] ;
 wire \mod_ro_128.fabric[119] ;
 wire \mod_ro_128.fabric[11] ;
 wire \mod_ro_128.fabric[120] ;
 wire \mod_ro_128.fabric[121] ;
 wire \mod_ro_128.fabric[122] ;
 wire \mod_ro_128.fabric[123] ;
 wire \mod_ro_128.fabric[124] ;
 wire \mod_ro_128.fabric[125] ;
 wire \mod_ro_128.fabric[126] ;
 wire \mod_ro_128.fabric[127] ;
 wire \mod_ro_128.fabric[128] ;
 wire \mod_ro_128.fabric[12] ;
 wire \mod_ro_128.fabric[13] ;
 wire \mod_ro_128.fabric[14] ;
 wire \mod_ro_128.fabric[15] ;
 wire \mod_ro_128.fabric[16] ;
 wire \mod_ro_128.fabric[17] ;
 wire \mod_ro_128.fabric[18] ;
 wire \mod_ro_128.fabric[19] ;
 wire \mod_ro_128.fabric[1] ;
 wire \mod_ro_128.fabric[20] ;
 wire \mod_ro_128.fabric[21] ;
 wire \mod_ro_128.fabric[22] ;
 wire \mod_ro_128.fabric[23] ;
 wire \mod_ro_128.fabric[24] ;
 wire \mod_ro_128.fabric[25] ;
 wire \mod_ro_128.fabric[26] ;
 wire \mod_ro_128.fabric[27] ;
 wire \mod_ro_128.fabric[28] ;
 wire \mod_ro_128.fabric[29] ;
 wire \mod_ro_128.fabric[2] ;
 wire \mod_ro_128.fabric[30] ;
 wire \mod_ro_128.fabric[31] ;
 wire \mod_ro_128.fabric[32] ;
 wire \mod_ro_128.fabric[33] ;
 wire \mod_ro_128.fabric[34] ;
 wire \mod_ro_128.fabric[35] ;
 wire \mod_ro_128.fabric[36] ;
 wire \mod_ro_128.fabric[37] ;
 wire \mod_ro_128.fabric[38] ;
 wire \mod_ro_128.fabric[39] ;
 wire \mod_ro_128.fabric[3] ;
 wire \mod_ro_128.fabric[40] ;
 wire \mod_ro_128.fabric[41] ;
 wire \mod_ro_128.fabric[42] ;
 wire \mod_ro_128.fabric[43] ;
 wire \mod_ro_128.fabric[44] ;
 wire \mod_ro_128.fabric[45] ;
 wire \mod_ro_128.fabric[46] ;
 wire \mod_ro_128.fabric[47] ;
 wire \mod_ro_128.fabric[48] ;
 wire \mod_ro_128.fabric[49] ;
 wire \mod_ro_128.fabric[4] ;
 wire \mod_ro_128.fabric[50] ;
 wire \mod_ro_128.fabric[51] ;
 wire \mod_ro_128.fabric[52] ;
 wire \mod_ro_128.fabric[53] ;
 wire \mod_ro_128.fabric[54] ;
 wire \mod_ro_128.fabric[55] ;
 wire \mod_ro_128.fabric[56] ;
 wire \mod_ro_128.fabric[57] ;
 wire \mod_ro_128.fabric[58] ;
 wire \mod_ro_128.fabric[59] ;
 wire \mod_ro_128.fabric[5] ;
 wire \mod_ro_128.fabric[60] ;
 wire \mod_ro_128.fabric[61] ;
 wire \mod_ro_128.fabric[62] ;
 wire \mod_ro_128.fabric[63] ;
 wire \mod_ro_128.fabric[64] ;
 wire \mod_ro_128.fabric[65] ;
 wire \mod_ro_128.fabric[66] ;
 wire \mod_ro_128.fabric[67] ;
 wire \mod_ro_128.fabric[68] ;
 wire \mod_ro_128.fabric[69] ;
 wire \mod_ro_128.fabric[6] ;
 wire \mod_ro_128.fabric[70] ;
 wire \mod_ro_128.fabric[71] ;
 wire \mod_ro_128.fabric[72] ;
 wire \mod_ro_128.fabric[73] ;
 wire \mod_ro_128.fabric[74] ;
 wire \mod_ro_128.fabric[75] ;
 wire \mod_ro_128.fabric[76] ;
 wire \mod_ro_128.fabric[77] ;
 wire \mod_ro_128.fabric[78] ;
 wire \mod_ro_128.fabric[79] ;
 wire \mod_ro_128.fabric[7] ;
 wire \mod_ro_128.fabric[80] ;
 wire \mod_ro_128.fabric[81] ;
 wire \mod_ro_128.fabric[82] ;
 wire \mod_ro_128.fabric[83] ;
 wire \mod_ro_128.fabric[84] ;
 wire \mod_ro_128.fabric[85] ;
 wire \mod_ro_128.fabric[86] ;
 wire \mod_ro_128.fabric[87] ;
 wire \mod_ro_128.fabric[88] ;
 wire \mod_ro_128.fabric[89] ;
 wire \mod_ro_128.fabric[8] ;
 wire \mod_ro_128.fabric[90] ;
 wire \mod_ro_128.fabric[91] ;
 wire \mod_ro_128.fabric[92] ;
 wire \mod_ro_128.fabric[93] ;
 wire \mod_ro_128.fabric[94] ;
 wire \mod_ro_128.fabric[95] ;
 wire \mod_ro_128.fabric[96] ;
 wire \mod_ro_128.fabric[97] ;
 wire \mod_ro_128.fabric[98] ;
 wire \mod_ro_128.fabric[99] ;
 wire \mod_ro_128.fabric[9] ;
 wire \mod_ro_16.fabric[0] ;
 wire \mod_ro_16.fabric[10] ;
 wire \mod_ro_16.fabric[11] ;
 wire \mod_ro_16.fabric[12] ;
 wire \mod_ro_16.fabric[13] ;
 wire \mod_ro_16.fabric[14] ;
 wire \mod_ro_16.fabric[15] ;
 wire \mod_ro_16.fabric[16] ;
 wire \mod_ro_16.fabric[1] ;
 wire \mod_ro_16.fabric[2] ;
 wire \mod_ro_16.fabric[3] ;
 wire \mod_ro_16.fabric[4] ;
 wire \mod_ro_16.fabric[5] ;
 wire \mod_ro_16.fabric[6] ;
 wire \mod_ro_16.fabric[7] ;
 wire \mod_ro_16.fabric[8] ;
 wire \mod_ro_16.fabric[9] ;
 wire \mod_ro_256.fabric[0] ;
 wire \mod_ro_256.fabric[100] ;
 wire \mod_ro_256.fabric[101] ;
 wire \mod_ro_256.fabric[102] ;
 wire \mod_ro_256.fabric[103] ;
 wire \mod_ro_256.fabric[104] ;
 wire \mod_ro_256.fabric[105] ;
 wire \mod_ro_256.fabric[106] ;
 wire \mod_ro_256.fabric[107] ;
 wire \mod_ro_256.fabric[108] ;
 wire \mod_ro_256.fabric[109] ;
 wire \mod_ro_256.fabric[10] ;
 wire \mod_ro_256.fabric[110] ;
 wire \mod_ro_256.fabric[111] ;
 wire \mod_ro_256.fabric[112] ;
 wire \mod_ro_256.fabric[113] ;
 wire \mod_ro_256.fabric[114] ;
 wire \mod_ro_256.fabric[115] ;
 wire \mod_ro_256.fabric[116] ;
 wire \mod_ro_256.fabric[117] ;
 wire \mod_ro_256.fabric[118] ;
 wire \mod_ro_256.fabric[119] ;
 wire \mod_ro_256.fabric[11] ;
 wire \mod_ro_256.fabric[120] ;
 wire \mod_ro_256.fabric[121] ;
 wire \mod_ro_256.fabric[122] ;
 wire \mod_ro_256.fabric[123] ;
 wire \mod_ro_256.fabric[124] ;
 wire \mod_ro_256.fabric[125] ;
 wire \mod_ro_256.fabric[126] ;
 wire \mod_ro_256.fabric[127] ;
 wire \mod_ro_256.fabric[128] ;
 wire \mod_ro_256.fabric[129] ;
 wire \mod_ro_256.fabric[12] ;
 wire \mod_ro_256.fabric[130] ;
 wire \mod_ro_256.fabric[131] ;
 wire \mod_ro_256.fabric[132] ;
 wire \mod_ro_256.fabric[133] ;
 wire \mod_ro_256.fabric[134] ;
 wire \mod_ro_256.fabric[135] ;
 wire \mod_ro_256.fabric[136] ;
 wire \mod_ro_256.fabric[137] ;
 wire \mod_ro_256.fabric[138] ;
 wire \mod_ro_256.fabric[139] ;
 wire \mod_ro_256.fabric[13] ;
 wire \mod_ro_256.fabric[140] ;
 wire \mod_ro_256.fabric[141] ;
 wire \mod_ro_256.fabric[142] ;
 wire \mod_ro_256.fabric[143] ;
 wire \mod_ro_256.fabric[144] ;
 wire \mod_ro_256.fabric[145] ;
 wire \mod_ro_256.fabric[146] ;
 wire \mod_ro_256.fabric[147] ;
 wire \mod_ro_256.fabric[148] ;
 wire \mod_ro_256.fabric[149] ;
 wire \mod_ro_256.fabric[14] ;
 wire \mod_ro_256.fabric[150] ;
 wire \mod_ro_256.fabric[151] ;
 wire \mod_ro_256.fabric[152] ;
 wire \mod_ro_256.fabric[153] ;
 wire \mod_ro_256.fabric[154] ;
 wire \mod_ro_256.fabric[155] ;
 wire \mod_ro_256.fabric[156] ;
 wire \mod_ro_256.fabric[157] ;
 wire \mod_ro_256.fabric[158] ;
 wire \mod_ro_256.fabric[159] ;
 wire \mod_ro_256.fabric[15] ;
 wire \mod_ro_256.fabric[160] ;
 wire \mod_ro_256.fabric[161] ;
 wire \mod_ro_256.fabric[162] ;
 wire \mod_ro_256.fabric[163] ;
 wire \mod_ro_256.fabric[164] ;
 wire \mod_ro_256.fabric[165] ;
 wire \mod_ro_256.fabric[166] ;
 wire \mod_ro_256.fabric[167] ;
 wire \mod_ro_256.fabric[168] ;
 wire \mod_ro_256.fabric[169] ;
 wire \mod_ro_256.fabric[16] ;
 wire \mod_ro_256.fabric[170] ;
 wire \mod_ro_256.fabric[171] ;
 wire \mod_ro_256.fabric[172] ;
 wire \mod_ro_256.fabric[173] ;
 wire \mod_ro_256.fabric[174] ;
 wire \mod_ro_256.fabric[175] ;
 wire \mod_ro_256.fabric[176] ;
 wire \mod_ro_256.fabric[177] ;
 wire \mod_ro_256.fabric[178] ;
 wire \mod_ro_256.fabric[179] ;
 wire \mod_ro_256.fabric[17] ;
 wire \mod_ro_256.fabric[180] ;
 wire \mod_ro_256.fabric[181] ;
 wire \mod_ro_256.fabric[182] ;
 wire \mod_ro_256.fabric[183] ;
 wire \mod_ro_256.fabric[184] ;
 wire \mod_ro_256.fabric[185] ;
 wire \mod_ro_256.fabric[186] ;
 wire \mod_ro_256.fabric[187] ;
 wire \mod_ro_256.fabric[188] ;
 wire \mod_ro_256.fabric[189] ;
 wire \mod_ro_256.fabric[18] ;
 wire \mod_ro_256.fabric[190] ;
 wire \mod_ro_256.fabric[191] ;
 wire \mod_ro_256.fabric[192] ;
 wire \mod_ro_256.fabric[193] ;
 wire \mod_ro_256.fabric[194] ;
 wire \mod_ro_256.fabric[195] ;
 wire \mod_ro_256.fabric[196] ;
 wire \mod_ro_256.fabric[197] ;
 wire \mod_ro_256.fabric[198] ;
 wire \mod_ro_256.fabric[199] ;
 wire \mod_ro_256.fabric[19] ;
 wire \mod_ro_256.fabric[1] ;
 wire \mod_ro_256.fabric[200] ;
 wire \mod_ro_256.fabric[201] ;
 wire \mod_ro_256.fabric[202] ;
 wire \mod_ro_256.fabric[203] ;
 wire \mod_ro_256.fabric[204] ;
 wire \mod_ro_256.fabric[205] ;
 wire \mod_ro_256.fabric[206] ;
 wire \mod_ro_256.fabric[207] ;
 wire \mod_ro_256.fabric[208] ;
 wire \mod_ro_256.fabric[209] ;
 wire \mod_ro_256.fabric[20] ;
 wire \mod_ro_256.fabric[210] ;
 wire \mod_ro_256.fabric[211] ;
 wire \mod_ro_256.fabric[212] ;
 wire \mod_ro_256.fabric[213] ;
 wire \mod_ro_256.fabric[214] ;
 wire \mod_ro_256.fabric[215] ;
 wire \mod_ro_256.fabric[216] ;
 wire \mod_ro_256.fabric[217] ;
 wire \mod_ro_256.fabric[218] ;
 wire \mod_ro_256.fabric[219] ;
 wire \mod_ro_256.fabric[21] ;
 wire \mod_ro_256.fabric[220] ;
 wire \mod_ro_256.fabric[221] ;
 wire \mod_ro_256.fabric[222] ;
 wire \mod_ro_256.fabric[223] ;
 wire \mod_ro_256.fabric[224] ;
 wire \mod_ro_256.fabric[225] ;
 wire \mod_ro_256.fabric[226] ;
 wire \mod_ro_256.fabric[227] ;
 wire \mod_ro_256.fabric[228] ;
 wire \mod_ro_256.fabric[229] ;
 wire \mod_ro_256.fabric[22] ;
 wire \mod_ro_256.fabric[230] ;
 wire \mod_ro_256.fabric[231] ;
 wire \mod_ro_256.fabric[232] ;
 wire \mod_ro_256.fabric[233] ;
 wire \mod_ro_256.fabric[234] ;
 wire \mod_ro_256.fabric[235] ;
 wire \mod_ro_256.fabric[236] ;
 wire \mod_ro_256.fabric[237] ;
 wire \mod_ro_256.fabric[238] ;
 wire \mod_ro_256.fabric[239] ;
 wire \mod_ro_256.fabric[23] ;
 wire \mod_ro_256.fabric[240] ;
 wire \mod_ro_256.fabric[241] ;
 wire \mod_ro_256.fabric[242] ;
 wire \mod_ro_256.fabric[243] ;
 wire \mod_ro_256.fabric[244] ;
 wire \mod_ro_256.fabric[245] ;
 wire \mod_ro_256.fabric[246] ;
 wire \mod_ro_256.fabric[247] ;
 wire \mod_ro_256.fabric[248] ;
 wire \mod_ro_256.fabric[249] ;
 wire \mod_ro_256.fabric[24] ;
 wire \mod_ro_256.fabric[250] ;
 wire \mod_ro_256.fabric[251] ;
 wire \mod_ro_256.fabric[252] ;
 wire \mod_ro_256.fabric[253] ;
 wire \mod_ro_256.fabric[254] ;
 wire \mod_ro_256.fabric[255] ;
 wire \mod_ro_256.fabric[256] ;
 wire \mod_ro_256.fabric[25] ;
 wire \mod_ro_256.fabric[26] ;
 wire \mod_ro_256.fabric[27] ;
 wire \mod_ro_256.fabric[28] ;
 wire \mod_ro_256.fabric[29] ;
 wire \mod_ro_256.fabric[2] ;
 wire \mod_ro_256.fabric[30] ;
 wire \mod_ro_256.fabric[31] ;
 wire \mod_ro_256.fabric[32] ;
 wire \mod_ro_256.fabric[33] ;
 wire \mod_ro_256.fabric[34] ;
 wire \mod_ro_256.fabric[35] ;
 wire \mod_ro_256.fabric[36] ;
 wire \mod_ro_256.fabric[37] ;
 wire \mod_ro_256.fabric[38] ;
 wire \mod_ro_256.fabric[39] ;
 wire \mod_ro_256.fabric[3] ;
 wire \mod_ro_256.fabric[40] ;
 wire \mod_ro_256.fabric[41] ;
 wire \mod_ro_256.fabric[42] ;
 wire \mod_ro_256.fabric[43] ;
 wire \mod_ro_256.fabric[44] ;
 wire \mod_ro_256.fabric[45] ;
 wire \mod_ro_256.fabric[46] ;
 wire \mod_ro_256.fabric[47] ;
 wire \mod_ro_256.fabric[48] ;
 wire \mod_ro_256.fabric[49] ;
 wire \mod_ro_256.fabric[4] ;
 wire \mod_ro_256.fabric[50] ;
 wire \mod_ro_256.fabric[51] ;
 wire \mod_ro_256.fabric[52] ;
 wire \mod_ro_256.fabric[53] ;
 wire \mod_ro_256.fabric[54] ;
 wire \mod_ro_256.fabric[55] ;
 wire \mod_ro_256.fabric[56] ;
 wire \mod_ro_256.fabric[57] ;
 wire \mod_ro_256.fabric[58] ;
 wire \mod_ro_256.fabric[59] ;
 wire \mod_ro_256.fabric[5] ;
 wire \mod_ro_256.fabric[60] ;
 wire \mod_ro_256.fabric[61] ;
 wire \mod_ro_256.fabric[62] ;
 wire \mod_ro_256.fabric[63] ;
 wire \mod_ro_256.fabric[64] ;
 wire \mod_ro_256.fabric[65] ;
 wire \mod_ro_256.fabric[66] ;
 wire \mod_ro_256.fabric[67] ;
 wire \mod_ro_256.fabric[68] ;
 wire \mod_ro_256.fabric[69] ;
 wire \mod_ro_256.fabric[6] ;
 wire \mod_ro_256.fabric[70] ;
 wire \mod_ro_256.fabric[71] ;
 wire \mod_ro_256.fabric[72] ;
 wire \mod_ro_256.fabric[73] ;
 wire \mod_ro_256.fabric[74] ;
 wire \mod_ro_256.fabric[75] ;
 wire \mod_ro_256.fabric[76] ;
 wire \mod_ro_256.fabric[77] ;
 wire \mod_ro_256.fabric[78] ;
 wire \mod_ro_256.fabric[79] ;
 wire \mod_ro_256.fabric[7] ;
 wire \mod_ro_256.fabric[80] ;
 wire \mod_ro_256.fabric[81] ;
 wire \mod_ro_256.fabric[82] ;
 wire \mod_ro_256.fabric[83] ;
 wire \mod_ro_256.fabric[84] ;
 wire \mod_ro_256.fabric[85] ;
 wire \mod_ro_256.fabric[86] ;
 wire \mod_ro_256.fabric[87] ;
 wire \mod_ro_256.fabric[88] ;
 wire \mod_ro_256.fabric[89] ;
 wire \mod_ro_256.fabric[8] ;
 wire \mod_ro_256.fabric[90] ;
 wire \mod_ro_256.fabric[91] ;
 wire \mod_ro_256.fabric[92] ;
 wire \mod_ro_256.fabric[93] ;
 wire \mod_ro_256.fabric[94] ;
 wire \mod_ro_256.fabric[95] ;
 wire \mod_ro_256.fabric[96] ;
 wire \mod_ro_256.fabric[97] ;
 wire \mod_ro_256.fabric[98] ;
 wire \mod_ro_256.fabric[99] ;
 wire \mod_ro_256.fabric[9] ;
 wire \mod_ro_31.fabric[0] ;
 wire \mod_ro_31.fabric[10] ;
 wire \mod_ro_31.fabric[11] ;
 wire \mod_ro_31.fabric[12] ;
 wire \mod_ro_31.fabric[13] ;
 wire \mod_ro_31.fabric[14] ;
 wire \mod_ro_31.fabric[15] ;
 wire \mod_ro_31.fabric[16] ;
 wire \mod_ro_31.fabric[17] ;
 wire \mod_ro_31.fabric[18] ;
 wire \mod_ro_31.fabric[19] ;
 wire \mod_ro_31.fabric[1] ;
 wire \mod_ro_31.fabric[20] ;
 wire \mod_ro_31.fabric[21] ;
 wire \mod_ro_31.fabric[22] ;
 wire \mod_ro_31.fabric[23] ;
 wire \mod_ro_31.fabric[24] ;
 wire \mod_ro_31.fabric[25] ;
 wire \mod_ro_31.fabric[26] ;
 wire \mod_ro_31.fabric[27] ;
 wire \mod_ro_31.fabric[28] ;
 wire \mod_ro_31.fabric[29] ;
 wire \mod_ro_31.fabric[2] ;
 wire \mod_ro_31.fabric[30] ;
 wire \mod_ro_31.fabric[31] ;
 wire \mod_ro_31.fabric[3] ;
 wire \mod_ro_31.fabric[4] ;
 wire \mod_ro_31.fabric[5] ;
 wire \mod_ro_31.fabric[6] ;
 wire \mod_ro_31.fabric[7] ;
 wire \mod_ro_31.fabric[8] ;
 wire \mod_ro_31.fabric[9] ;
 wire \mod_ro_32_1.fabric[0] ;
 wire \mod_ro_32_1.fabric[10] ;
 wire \mod_ro_32_1.fabric[11] ;
 wire \mod_ro_32_1.fabric[12] ;
 wire \mod_ro_32_1.fabric[13] ;
 wire \mod_ro_32_1.fabric[14] ;
 wire \mod_ro_32_1.fabric[15] ;
 wire \mod_ro_32_1.fabric[16] ;
 wire \mod_ro_32_1.fabric[17] ;
 wire \mod_ro_32_1.fabric[18] ;
 wire \mod_ro_32_1.fabric[19] ;
 wire \mod_ro_32_1.fabric[1] ;
 wire \mod_ro_32_1.fabric[20] ;
 wire \mod_ro_32_1.fabric[21] ;
 wire \mod_ro_32_1.fabric[22] ;
 wire \mod_ro_32_1.fabric[23] ;
 wire \mod_ro_32_1.fabric[24] ;
 wire \mod_ro_32_1.fabric[25] ;
 wire \mod_ro_32_1.fabric[26] ;
 wire \mod_ro_32_1.fabric[27] ;
 wire \mod_ro_32_1.fabric[28] ;
 wire \mod_ro_32_1.fabric[29] ;
 wire \mod_ro_32_1.fabric[2] ;
 wire \mod_ro_32_1.fabric[30] ;
 wire \mod_ro_32_1.fabric[31] ;
 wire \mod_ro_32_1.fabric[32] ;
 wire \mod_ro_32_1.fabric[3] ;
 wire \mod_ro_32_1.fabric[4] ;
 wire \mod_ro_32_1.fabric[5] ;
 wire \mod_ro_32_1.fabric[6] ;
 wire \mod_ro_32_1.fabric[7] ;
 wire \mod_ro_32_1.fabric[8] ;
 wire \mod_ro_32_1.fabric[9] ;
 wire \mod_ro_32_2.fabric[0] ;
 wire \mod_ro_32_2.fabric[10] ;
 wire \mod_ro_32_2.fabric[11] ;
 wire \mod_ro_32_2.fabric[12] ;
 wire \mod_ro_32_2.fabric[13] ;
 wire \mod_ro_32_2.fabric[14] ;
 wire \mod_ro_32_2.fabric[15] ;
 wire \mod_ro_32_2.fabric[16] ;
 wire \mod_ro_32_2.fabric[17] ;
 wire \mod_ro_32_2.fabric[18] ;
 wire \mod_ro_32_2.fabric[19] ;
 wire \mod_ro_32_2.fabric[1] ;
 wire \mod_ro_32_2.fabric[20] ;
 wire \mod_ro_32_2.fabric[21] ;
 wire \mod_ro_32_2.fabric[22] ;
 wire \mod_ro_32_2.fabric[23] ;
 wire \mod_ro_32_2.fabric[24] ;
 wire \mod_ro_32_2.fabric[25] ;
 wire \mod_ro_32_2.fabric[26] ;
 wire \mod_ro_32_2.fabric[27] ;
 wire \mod_ro_32_2.fabric[28] ;
 wire \mod_ro_32_2.fabric[29] ;
 wire \mod_ro_32_2.fabric[2] ;
 wire \mod_ro_32_2.fabric[30] ;
 wire \mod_ro_32_2.fabric[31] ;
 wire \mod_ro_32_2.fabric[32] ;
 wire \mod_ro_32_2.fabric[3] ;
 wire \mod_ro_32_2.fabric[4] ;
 wire \mod_ro_32_2.fabric[5] ;
 wire \mod_ro_32_2.fabric[6] ;
 wire \mod_ro_32_2.fabric[7] ;
 wire \mod_ro_32_2.fabric[8] ;
 wire \mod_ro_32_2.fabric[9] ;
 wire \mod_ro_32_raw.fabric[0] ;
 wire \mod_ro_32_raw.fabric[10] ;
 wire \mod_ro_32_raw.fabric[11] ;
 wire \mod_ro_32_raw.fabric[12] ;
 wire \mod_ro_32_raw.fabric[13] ;
 wire \mod_ro_32_raw.fabric[14] ;
 wire \mod_ro_32_raw.fabric[15] ;
 wire \mod_ro_32_raw.fabric[16] ;
 wire \mod_ro_32_raw.fabric[17] ;
 wire \mod_ro_32_raw.fabric[18] ;
 wire \mod_ro_32_raw.fabric[19] ;
 wire \mod_ro_32_raw.fabric[1] ;
 wire \mod_ro_32_raw.fabric[20] ;
 wire \mod_ro_32_raw.fabric[21] ;
 wire \mod_ro_32_raw.fabric[22] ;
 wire \mod_ro_32_raw.fabric[23] ;
 wire \mod_ro_32_raw.fabric[24] ;
 wire \mod_ro_32_raw.fabric[25] ;
 wire \mod_ro_32_raw.fabric[26] ;
 wire \mod_ro_32_raw.fabric[27] ;
 wire \mod_ro_32_raw.fabric[28] ;
 wire \mod_ro_32_raw.fabric[29] ;
 wire \mod_ro_32_raw.fabric[2] ;
 wire \mod_ro_32_raw.fabric[30] ;
 wire \mod_ro_32_raw.fabric[31] ;
 wire \mod_ro_32_raw.fabric[32] ;
 wire \mod_ro_32_raw.fabric[3] ;
 wire \mod_ro_32_raw.fabric[4] ;
 wire \mod_ro_32_raw.fabric[5] ;
 wire \mod_ro_32_raw.fabric[6] ;
 wire \mod_ro_32_raw.fabric[7] ;
 wire \mod_ro_32_raw.fabric[8] ;
 wire \mod_ro_32_raw.fabric[9] ;
 wire \mod_ro_64.fabric[0] ;
 wire \mod_ro_64.fabric[10] ;
 wire \mod_ro_64.fabric[11] ;
 wire \mod_ro_64.fabric[12] ;
 wire \mod_ro_64.fabric[13] ;
 wire \mod_ro_64.fabric[14] ;
 wire \mod_ro_64.fabric[15] ;
 wire \mod_ro_64.fabric[16] ;
 wire \mod_ro_64.fabric[17] ;
 wire \mod_ro_64.fabric[18] ;
 wire \mod_ro_64.fabric[19] ;
 wire \mod_ro_64.fabric[1] ;
 wire \mod_ro_64.fabric[20] ;
 wire \mod_ro_64.fabric[21] ;
 wire \mod_ro_64.fabric[22] ;
 wire \mod_ro_64.fabric[23] ;
 wire \mod_ro_64.fabric[24] ;
 wire \mod_ro_64.fabric[25] ;
 wire \mod_ro_64.fabric[26] ;
 wire \mod_ro_64.fabric[27] ;
 wire \mod_ro_64.fabric[28] ;
 wire \mod_ro_64.fabric[29] ;
 wire \mod_ro_64.fabric[2] ;
 wire \mod_ro_64.fabric[30] ;
 wire \mod_ro_64.fabric[31] ;
 wire \mod_ro_64.fabric[32] ;
 wire \mod_ro_64.fabric[33] ;
 wire \mod_ro_64.fabric[34] ;
 wire \mod_ro_64.fabric[35] ;
 wire \mod_ro_64.fabric[36] ;
 wire \mod_ro_64.fabric[37] ;
 wire \mod_ro_64.fabric[38] ;
 wire \mod_ro_64.fabric[39] ;
 wire \mod_ro_64.fabric[3] ;
 wire \mod_ro_64.fabric[40] ;
 wire \mod_ro_64.fabric[41] ;
 wire \mod_ro_64.fabric[42] ;
 wire \mod_ro_64.fabric[43] ;
 wire \mod_ro_64.fabric[44] ;
 wire \mod_ro_64.fabric[45] ;
 wire \mod_ro_64.fabric[46] ;
 wire \mod_ro_64.fabric[47] ;
 wire \mod_ro_64.fabric[48] ;
 wire \mod_ro_64.fabric[49] ;
 wire \mod_ro_64.fabric[4] ;
 wire \mod_ro_64.fabric[50] ;
 wire \mod_ro_64.fabric[51] ;
 wire \mod_ro_64.fabric[52] ;
 wire \mod_ro_64.fabric[53] ;
 wire \mod_ro_64.fabric[54] ;
 wire \mod_ro_64.fabric[55] ;
 wire \mod_ro_64.fabric[56] ;
 wire \mod_ro_64.fabric[57] ;
 wire \mod_ro_64.fabric[58] ;
 wire \mod_ro_64.fabric[59] ;
 wire \mod_ro_64.fabric[5] ;
 wire \mod_ro_64.fabric[60] ;
 wire \mod_ro_64.fabric[61] ;
 wire \mod_ro_64.fabric[62] ;
 wire \mod_ro_64.fabric[63] ;
 wire \mod_ro_64.fabric[64] ;
 wire \mod_ro_64.fabric[6] ;
 wire \mod_ro_64.fabric[7] ;
 wire \mod_ro_64.fabric[8] ;
 wire \mod_ro_64.fabric[9] ;
 wire mux_out;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_0_clk_regs;
 wire clknet_2_0__leaf_clk_regs;
 wire clknet_2_1__leaf_clk_regs;
 wire clknet_2_2__leaf_clk_regs;
 wire clknet_2_3__leaf_clk_regs;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;

 sg13g2_a21oi_1 _133_ (.A1(\dpll.id_decrement ),
    .A2(net56),
    .Y(_010_),
    .B1(_024_));
 sg13g2_o21ai_1 _134_ (.B1(net18),
    .Y(_025_),
    .A1(\dpll.id_increment ),
    .A2(\dpll.k_count_carry ));
 sg13g2_a21oi_1 _135_ (.A1(\dpll.id_increment ),
    .A2(net54),
    .Y(_011_),
    .B1(_025_));
 sg13g2_xor2_1 _136_ (.B(net4),
    .A(net86),
    .X(_026_));
 sg13g2_and2_1 _137_ (.A(net17),
    .B(_026_),
    .X(_027_));
 sg13g2_nand2_2 _138_ (.Y(_028_),
    .A(net17),
    .B(_026_));
 sg13g2_nor2_2 _139_ (.A(_081_),
    .B(_026_),
    .Y(_029_));
 sg13g2_nand2_1 _140_ (.Y(_030_),
    .A(net79),
    .B(net13));
 sg13g2_o21ai_1 _141_ (.B1(_030_),
    .Y(_012_),
    .A1(net79),
    .A2(_028_));
 sg13g2_nand2_1 _142_ (.Y(_031_),
    .A(net81),
    .B(net13));
 sg13g2_nor2b_1 _143_ (.A(net14),
    .B_N(net81),
    .Y(_032_));
 sg13g2_xnor2_1 _144_ (.Y(_033_),
    .A(net81),
    .B(net14));
 sg13g2_xnor2_1 _145_ (.Y(_034_),
    .A(net79),
    .B(_033_));
 sg13g2_o21ai_1 _146_ (.B1(_031_),
    .Y(_013_),
    .A1(_028_),
    .A2(_034_));
 sg13g2_nand2_1 _147_ (.Y(_035_),
    .A(net89),
    .B(net13));
 sg13g2_a21oi_2 _148_ (.B1(_032_),
    .Y(_036_),
    .A2(_033_),
    .A1(net79));
 sg13g2_nand2_1 _149_ (.Y(_037_),
    .A(net89),
    .B(_078_));
 sg13g2_xor2_1 _150_ (.B(net14),
    .A(net89),
    .X(_038_));
 sg13g2_xnor2_1 _151_ (.Y(_039_),
    .A(_036_),
    .B(_038_));
 sg13g2_o21ai_1 _152_ (.B1(_035_),
    .Y(_014_),
    .A1(_028_),
    .A2(_039_));
 sg13g2_xnor2_1 _153_ (.Y(_040_),
    .A(net90),
    .B(net14));
 sg13g2_o21ai_1 _154_ (.B1(_037_),
    .Y(_041_),
    .A1(_036_),
    .A2(_038_));
 sg13g2_o21ai_1 _155_ (.B1(_027_),
    .Y(_042_),
    .A1(_040_),
    .A2(_041_));
 sg13g2_a21oi_1 _156_ (.A1(_040_),
    .A2(_041_),
    .Y(_043_),
    .B1(_042_));
 sg13g2_a21oi_1 _157_ (.A1(net90),
    .A2(net13),
    .Y(_044_),
    .B1(_043_));
 sg13g2_inv_1 _158_ (.Y(_015_),
    .A(_044_));
 sg13g2_nand2_1 _159_ (.Y(_045_),
    .A(net71),
    .B(net13));
 sg13g2_nand2b_1 _160_ (.Y(_046_),
    .B(_040_),
    .A_N(_038_));
 sg13g2_o21ai_1 _161_ (.B1(_078_),
    .Y(_047_),
    .A1(\dpll.k_count[3] ),
    .A2(\dpll.k_count[2] ));
 sg13g2_o21ai_1 _162_ (.B1(_047_),
    .Y(_048_),
    .A1(_036_),
    .A2(_046_));
 sg13g2_nor2b_1 _163_ (.A(net14),
    .B_N(net71),
    .Y(_049_));
 sg13g2_nand2b_1 _164_ (.Y(_050_),
    .B(net14),
    .A_N(net71));
 sg13g2_nand2b_1 _165_ (.Y(_051_),
    .B(_050_),
    .A_N(_049_));
 sg13g2_xor2_1 _166_ (.B(_051_),
    .A(_048_),
    .X(_052_));
 sg13g2_o21ai_1 _167_ (.B1(_045_),
    .Y(_016_),
    .A1(_028_),
    .A2(_052_));
 sg13g2_nand2_1 _168_ (.Y(_053_),
    .A(net77),
    .B(net13));
 sg13g2_xor2_1 _169_ (.B(net14),
    .A(net77),
    .X(_054_));
 sg13g2_a21oi_1 _170_ (.A1(_048_),
    .A2(_050_),
    .Y(_055_),
    .B1(_049_));
 sg13g2_xnor2_1 _171_ (.Y(_056_),
    .A(_054_),
    .B(_055_));
 sg13g2_o21ai_1 _172_ (.B1(_053_),
    .Y(_017_),
    .A1(_028_),
    .A2(_056_));
 sg13g2_nand2_1 _173_ (.Y(_057_),
    .A(net75),
    .B(_029_));
 sg13g2_nand2_1 _174_ (.Y(_058_),
    .A(\dpll.k_count[6] ),
    .B(_078_));
 sg13g2_xor2_1 _175_ (.B(net15),
    .A(net75),
    .X(_059_));
 sg13g2_nor2_1 _176_ (.A(_051_),
    .B(_054_),
    .Y(_060_));
 sg13g2_a221oi_1 _177_ (.B2(_060_),
    .C1(_049_),
    .B1(_048_),
    .A1(\dpll.k_count[5] ),
    .Y(_061_),
    .A2(_078_));
 sg13g2_xnor2_1 _178_ (.Y(_062_),
    .A(_059_),
    .B(_061_));
 sg13g2_o21ai_1 _179_ (.B1(_057_),
    .Y(_018_),
    .A1(_028_),
    .A2(_062_));
 sg13g2_nand2_1 _180_ (.Y(_063_),
    .A(net73),
    .B(_029_));
 sg13g2_o21ai_1 _181_ (.B1(_058_),
    .Y(_064_),
    .A1(_059_),
    .A2(_061_));
 sg13g2_xnor2_1 _182_ (.Y(_065_),
    .A(net73),
    .B(net15));
 sg13g2_xnor2_1 _183_ (.Y(_066_),
    .A(_064_),
    .B(_065_));
 sg13g2_o21ai_1 _184_ (.B1(_063_),
    .Y(_019_),
    .A1(_028_),
    .A2(_066_));
 sg13g2_nand2_1 _185_ (.Y(_067_),
    .A(_078_),
    .B(net17));
 sg13g2_nor4_1 _186_ (.A(\dpll.k_count[3] ),
    .B(\dpll.k_count[2] ),
    .C(\dpll.k_count[1] ),
    .D(\dpll.k_count[0] ),
    .Y(_068_));
 sg13g2_nor4_1 _187_ (.A(\dpll.k_count[7] ),
    .B(\dpll.k_count[6] ),
    .C(\dpll.k_count[5] ),
    .D(\dpll.k_count[4] ),
    .Y(_069_));
 sg13g2_a21oi_1 _188_ (.A1(_068_),
    .A2(_069_),
    .Y(_070_),
    .B1(_067_));
 sg13g2_a21oi_1 _189_ (.A1(_078_),
    .A2(net18),
    .Y(_071_),
    .B1(net58));
 sg13g2_nor3_1 _190_ (.A(net13),
    .B(_070_),
    .C(net59),
    .Y(_020_));
 sg13g2_nand4_1 _191_ (.B(\dpll.k_count[2] ),
    .C(\dpll.k_count[1] ),
    .A(\dpll.k_count[3] ),
    .Y(_072_),
    .D(\dpll.k_count[0] ));
 sg13g2_nand4_1 _192_ (.B(\dpll.k_count[6] ),
    .C(\dpll.k_count[5] ),
    .A(\dpll.k_count[7] ),
    .Y(_073_),
    .D(\dpll.k_count[4] ));
 sg13g2_nor2_1 _193_ (.A(_072_),
    .B(_073_),
    .Y(_074_));
 sg13g2_nor3_1 _194_ (.A(_078_),
    .B(_081_),
    .C(_074_),
    .Y(_075_));
 sg13g2_a21oi_1 _195_ (.A1(net15),
    .A2(net18),
    .Y(_076_),
    .B1(net64));
 sg13g2_nor3_1 _196_ (.A(net13),
    .B(_075_),
    .C(net65),
    .Y(_021_));
 sg13g2_inv_1 _197_ (.Y(_077_),
    .A(net86));
 sg13g2_inv_4 _198_ (.A(net14),
    .Y(_078_));
 sg13g2_inv_1 _199_ (.Y(_079_),
    .A(net88));
 sg13g2_inv_1 _200_ (.Y(_080_),
    .A(net67));
 sg13g2_inv_4 _201_ (.A(net17),
    .Y(_081_));
 sg13g2_inv_1 _202_ (.Y(_082_),
    .A(\mod_ro_256.fabric[0] ));
 sg13g2_or2_1 _203_ (.X(_083_),
    .B(\mod_ro_32_2.fabric[0] ),
    .A(net3));
 sg13g2_nand2b_1 _204_ (.Y(_084_),
    .B(net3),
    .A_N(\mod_ro_31.fabric[0] ));
 sg13g2_nand3_1 _205_ (.B(_083_),
    .C(_084_),
    .A(net1),
    .Y(_085_));
 sg13g2_a21oi_1 _206_ (.A1(net3),
    .A2(\mod_ro_32_2.fabric[0] ),
    .Y(_086_),
    .B1(\mod_ro_32_1.fabric[0] ));
 sg13g2_nor2_1 _207_ (.A(net1),
    .B(_086_),
    .Y(_087_));
 sg13g2_nor2_1 _208_ (.A(net2),
    .B(_087_),
    .Y(_088_));
 sg13g2_nand2b_1 _209_ (.Y(_089_),
    .B(net3),
    .A_N(\mod_ro_128.fabric[0] ));
 sg13g2_o21ai_1 _210_ (.B1(_089_),
    .Y(_090_),
    .A1(net3),
    .A2(\mod_ro_64.fabric[0] ));
 sg13g2_o21ai_1 _211_ (.B1(net1),
    .Y(_091_),
    .A1(net3),
    .A2(\mod_ro_16.fabric[0] ));
 sg13g2_a21oi_1 _212_ (.A1(net3),
    .A2(_082_),
    .Y(_092_),
    .B1(_091_));
 sg13g2_o21ai_1 _213_ (.B1(net2),
    .Y(_093_),
    .A1(net1),
    .A2(_090_));
 sg13g2_nor2_1 _214_ (.A(_092_),
    .B(_093_),
    .Y(_094_));
 sg13g2_a21oi_1 _215_ (.A1(_085_),
    .A2(_088_),
    .Y(mux_out),
    .B1(_094_));
 sg13g2_nand2_1 _216_ (.Y(_095_),
    .A(net70),
    .B(net16));
 sg13g2_nor2_1 _217_ (.A(net69),
    .B(net16),
    .Y(_096_));
 sg13g2_a21oi_1 _218_ (.A1(net70),
    .A2(net16),
    .Y(_097_),
    .B1(_096_));
 sg13g2_nor2_1 _219_ (.A(_081_),
    .B(_097_),
    .Y(_000_));
 sg13g2_o21ai_1 _220_ (.B1(net17),
    .Y(_098_),
    .A1(net16),
    .A2(\dpll.n_count[0] ));
 sg13g2_a21oi_1 _221_ (.A1(net52),
    .A2(\dpll.n_count[0] ),
    .Y(_001_),
    .B1(_098_));
 sg13g2_a21oi_1 _222_ (.A1(net16),
    .A2(\dpll.n_count[0] ),
    .Y(_099_),
    .B1(net61));
 sg13g2_nand3_1 _223_ (.B(net61),
    .C(net91),
    .A(net16),
    .Y(_100_));
 sg13g2_nand2_1 _224_ (.Y(_101_),
    .A(net18),
    .B(_100_));
 sg13g2_nor2_1 _225_ (.A(net62),
    .B(_101_),
    .Y(_002_));
 sg13g2_or2_1 _226_ (.X(_102_),
    .B(_100_),
    .A(_080_));
 sg13g2_nand2_1 _227_ (.Y(_103_),
    .A(net17),
    .B(_102_));
 sg13g2_a21oi_1 _228_ (.A1(_080_),
    .A2(_100_),
    .Y(_003_),
    .B1(_103_));
 sg13g2_and2_1 _229_ (.A(_079_),
    .B(_102_),
    .X(_104_));
 sg13g2_nor2_2 _230_ (.A(_079_),
    .B(_102_),
    .Y(_105_));
 sg13g2_nor3_1 _231_ (.A(_081_),
    .B(_104_),
    .C(_105_),
    .Y(_004_));
 sg13g2_xnor2_1 _232_ (.Y(_106_),
    .A(net83),
    .B(_105_));
 sg13g2_nor2_1 _233_ (.A(_081_),
    .B(_106_),
    .Y(_005_));
 sg13g2_a21oi_1 _234_ (.A1(net83),
    .A2(_105_),
    .Y(_107_),
    .B1(net15));
 sg13g2_nand3_1 _235_ (.B(net83),
    .C(_105_),
    .A(net15),
    .Y(_108_));
 sg13g2_nand2_1 _236_ (.Y(_109_),
    .A(net17),
    .B(_108_));
 sg13g2_nor2_1 _237_ (.A(net84),
    .B(_109_),
    .Y(_006_));
 sg13g2_o21ai_1 _238_ (.B1(net17),
    .Y(_110_),
    .A1(_077_),
    .A2(_108_));
 sg13g2_a21oi_1 _239_ (.A1(_077_),
    .A2(_108_),
    .Y(_007_),
    .B1(_110_));
 sg13g2_nand2b_1 _240_ (.Y(_022_),
    .B(net54),
    .A_N(net16));
 sg13g2_a21oi_1 _241_ (.A1(_095_),
    .A2(_022_),
    .Y(_008_),
    .B1(_081_));
 sg13g2_nor2b_1 _242_ (.A(net56),
    .B_N(net16),
    .Y(_023_));
 sg13g2_nor3_1 _243_ (.A(_081_),
    .B(_096_),
    .C(_023_),
    .Y(_009_));
 sg13g2_o21ai_1 _244_ (.B1(net18),
    .Y(_024_),
    .A1(\dpll.id_decrement ),
    .A2(\dpll.k_count_borrow ));
 sg13g2_dfrbpq_1 _245_ (.RESET_B(net39),
    .D(_000_),
    .Q(\dpll.id_out ),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _246_ (.RESET_B(net50),
    .D(net53),
    .Q(\dpll.n_count[0] ),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _247_ (.RESET_B(net48),
    .D(net63),
    .Q(\dpll.n_count[1] ),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _248_ (.RESET_B(net46),
    .D(net68),
    .Q(\dpll.n_count[2] ),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _249_ (.RESET_B(net44),
    .D(_004_),
    .Q(\dpll.clk8x_fout ),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _250_ (.RESET_B(net42),
    .D(_005_),
    .Q(\dpll.n_count[4] ),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _251_ (.RESET_B(net40),
    .D(net85),
    .Q(\dpll.n_count[5] ),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_dfrbpq_1 _252_ (.RESET_B(net38),
    .D(net87),
    .Q(\dpll.clk_fout ),
    .CLK(clknet_2_0__leaf_clk_regs));
 sg13g2_dfrbpq_1 _253_ (.RESET_B(net36),
    .D(_008_),
    .Q(\dpll.id_increment_done ),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_dfrbpq_1 _254_ (.RESET_B(net34),
    .D(_009_),
    .Q(\dpll.id_decrement_done ),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _255_ (.RESET_B(net32),
    .D(net57),
    .Q(\dpll.id_decrement ),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _256_ (.RESET_B(net30),
    .D(net55),
    .Q(\dpll.id_increment ),
    .CLK(clknet_2_3__leaf_clk_regs));
 sg13g2_dfrbpq_2 _257_ (.RESET_B(net49),
    .D(net80),
    .Q(\dpll.k_count[0] ),
    .CLK(clknet_2_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _258_ (.RESET_B(net45),
    .D(net82),
    .Q(\dpll.k_count[1] ),
    .CLK(clknet_2_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _259_ (.RESET_B(net41),
    .D(_014_),
    .Q(\dpll.k_count[2] ),
    .CLK(clknet_2_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _260_ (.RESET_B(net37),
    .D(_015_),
    .Q(\dpll.k_count[3] ),
    .CLK(clknet_2_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _261_ (.RESET_B(net33),
    .D(net72),
    .Q(\dpll.k_count[4] ),
    .CLK(clknet_2_0__leaf_clk_regs));
 sg13g2_dfrbpq_2 _262_ (.RESET_B(net51),
    .D(net78),
    .Q(\dpll.k_count[5] ),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _263_ (.RESET_B(net43),
    .D(net76),
    .Q(\dpll.k_count[6] ),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_dfrbpq_2 _264_ (.RESET_B(net35),
    .D(net74),
    .Q(\dpll.k_count[7] ),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _265_ (.RESET_B(net47),
    .D(net60),
    .Q(\dpll.k_count_borrow ),
    .CLK(clknet_2_2__leaf_clk_regs));
 sg13g2_dfrbpq_1 _266_ (.RESET_B(net31),
    .D(net66),
    .Q(\dpll.k_count_carry ),
    .CLK(clknet_2_1__leaf_clk_regs));
 sg13g2_tiehi _266__25 (.L_HI(net31));
 sg13g2_tiehi _255__26 (.L_HI(net32));
 sg13g2_tiehi _261__27 (.L_HI(net33));
 sg13g2_tiehi _254__28 (.L_HI(net34));
 sg13g2_tiehi _264__29 (.L_HI(net35));
 sg13g2_tiehi _253__30 (.L_HI(net36));
 sg13g2_tiehi _260__31 (.L_HI(net37));
 sg13g2_tiehi _252__32 (.L_HI(net38));
 sg13g2_tiehi _245__33 (.L_HI(net39));
 sg13g2_tiehi _251__34 (.L_HI(net40));
 sg13g2_tiehi _259__35 (.L_HI(net41));
 sg13g2_tiehi _250__36 (.L_HI(net42));
 sg13g2_tiehi _263__37 (.L_HI(net43));
 sg13g2_tiehi _249__38 (.L_HI(net44));
 sg13g2_tiehi _258__39 (.L_HI(net45));
 sg13g2_tiehi _248__40 (.L_HI(net46));
 sg13g2_tiehi _265__41 (.L_HI(net47));
 sg13g2_tiehi _247__42 (.L_HI(net48));
 sg13g2_tiehi _257__43 (.L_HI(net49));
 sg13g2_tiehi _246__44 (.L_HI(net50));
 sg13g2_tiehi _262__45 (.L_HI(net51));
 sg13g2_buf_8 clkbuf_regs_0_clk (.A(clk),
    .X(clk_regs));
 sg13g2_tielo tt_um_wedgetail_tester_6 (.L_LO(net6));
 sg13g2_tielo tt_um_wedgetail_tester_7 (.L_LO(net7));
 sg13g2_tielo tt_um_wedgetail_tester_8 (.L_LO(net8));
 sg13g2_tielo tt_um_wedgetail_tester_9 (.L_LO(net9));
 sg13g2_tielo tt_um_wedgetail_tester_10 (.L_LO(net10));
 sg13g2_tielo tt_um_wedgetail_tester_11 (.L_LO(net11));
 sg13g2_tielo tt_um_wedgetail_tester_12 (.L_LO(net12));
 sg13g2_tielo tt_um_wedgetail_tester_13 (.L_LO(net19));
 sg13g2_tielo tt_um_wedgetail_tester_14 (.L_LO(net20));
 sg13g2_tielo tt_um_wedgetail_tester_15 (.L_LO(net21));
 sg13g2_tielo tt_um_wedgetail_tester_16 (.L_LO(net22));
 sg13g2_tielo tt_um_wedgetail_tester_17 (.L_LO(net23));
 sg13g2_tielo tt_um_wedgetail_tester_18 (.L_LO(net24));
 sg13g2_tielo tt_um_wedgetail_tester_19 (.L_LO(net25));
 sg13g2_tielo tt_um_wedgetail_tester_20 (.L_LO(net26));
 sg13g2_tielo tt_um_wedgetail_tester_21 (.L_LO(net27));
 sg13g2_tielo tt_um_wedgetail_tester_22 (.L_LO(net28));
 sg13g2_tielo tt_um_wedgetail_tester_23 (.L_LO(net29));
 sg13g2_tiehi _256__24 (.L_HI(net30));
 sg13g2_buf_1 _308_ (.A(mux_out),
    .X(uo_out[0]));
 sg13g2_buf_1 _309_ (.A(clknet_1_0__leaf_clk),
    .X(uo_out[1]));
 sg13g2_buf_1 _310_ (.A(\mod_ro_32_raw.fabric[0] ),
    .X(uo_out[2]));
 sg13g2_buf_1 _311_ (.A(\dpll.clk_fout ),
    .X(uo_out[3]));
 sg13g2_buf_1 _312_ (.A(\dpll.clk8x_fout ),
    .X(uo_out[4]));
 sg13g2_inv_1 \mod_ro_128.feedback  (.Y(\mod_ro_128.fabric[0] ),
    .A(\mod_ro_128.fabric[128] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[0].inv  (.Y(\mod_ro_128.fabric[1] ),
    .A(\mod_ro_128.fabric[0] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[100].inv  (.Y(\mod_ro_128.fabric[101] ),
    .A(\mod_ro_128.fabric[100] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[101].inv  (.Y(\mod_ro_128.fabric[102] ),
    .A(\mod_ro_128.fabric[101] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[102].inv  (.Y(\mod_ro_128.fabric[103] ),
    .A(\mod_ro_128.fabric[102] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[103].inv  (.Y(\mod_ro_128.fabric[104] ),
    .A(\mod_ro_128.fabric[103] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[104].inv  (.Y(\mod_ro_128.fabric[105] ),
    .A(\mod_ro_128.fabric[104] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[105].inv  (.Y(\mod_ro_128.fabric[106] ),
    .A(\mod_ro_128.fabric[105] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[106].inv  (.Y(\mod_ro_128.fabric[107] ),
    .A(\mod_ro_128.fabric[106] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[107].inv  (.Y(\mod_ro_128.fabric[108] ),
    .A(\mod_ro_128.fabric[107] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[108].inv  (.Y(\mod_ro_128.fabric[109] ),
    .A(\mod_ro_128.fabric[108] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[109].inv  (.Y(\mod_ro_128.fabric[110] ),
    .A(\mod_ro_128.fabric[109] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[10].inv  (.Y(\mod_ro_128.fabric[11] ),
    .A(\mod_ro_128.fabric[10] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[110].inv  (.Y(\mod_ro_128.fabric[111] ),
    .A(\mod_ro_128.fabric[110] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[111].inv  (.Y(\mod_ro_128.fabric[112] ),
    .A(\mod_ro_128.fabric[111] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[112].inv  (.Y(\mod_ro_128.fabric[113] ),
    .A(\mod_ro_128.fabric[112] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[113].inv  (.Y(\mod_ro_128.fabric[114] ),
    .A(\mod_ro_128.fabric[113] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[114].inv  (.Y(\mod_ro_128.fabric[115] ),
    .A(\mod_ro_128.fabric[114] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[115].inv  (.Y(\mod_ro_128.fabric[116] ),
    .A(\mod_ro_128.fabric[115] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[116].inv  (.Y(\mod_ro_128.fabric[117] ),
    .A(\mod_ro_128.fabric[116] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[117].inv  (.Y(\mod_ro_128.fabric[118] ),
    .A(\mod_ro_128.fabric[117] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[118].inv  (.Y(\mod_ro_128.fabric[119] ),
    .A(\mod_ro_128.fabric[118] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[119].inv  (.Y(\mod_ro_128.fabric[120] ),
    .A(\mod_ro_128.fabric[119] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[11].inv  (.Y(\mod_ro_128.fabric[12] ),
    .A(\mod_ro_128.fabric[11] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[120].inv  (.Y(\mod_ro_128.fabric[121] ),
    .A(\mod_ro_128.fabric[120] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[121].inv  (.Y(\mod_ro_128.fabric[122] ),
    .A(\mod_ro_128.fabric[121] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[122].inv  (.Y(\mod_ro_128.fabric[123] ),
    .A(\mod_ro_128.fabric[122] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[123].inv  (.Y(\mod_ro_128.fabric[124] ),
    .A(\mod_ro_128.fabric[123] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[124].inv  (.Y(\mod_ro_128.fabric[125] ),
    .A(\mod_ro_128.fabric[124] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[125].inv  (.Y(\mod_ro_128.fabric[126] ),
    .A(\mod_ro_128.fabric[125] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[126].inv  (.Y(\mod_ro_128.fabric[127] ),
    .A(\mod_ro_128.fabric[126] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[127].inv  (.Y(\mod_ro_128.fabric[128] ),
    .A(\mod_ro_128.fabric[127] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[12].inv  (.Y(\mod_ro_128.fabric[13] ),
    .A(\mod_ro_128.fabric[12] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[13].inv  (.Y(\mod_ro_128.fabric[14] ),
    .A(\mod_ro_128.fabric[13] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[14].inv  (.Y(\mod_ro_128.fabric[15] ),
    .A(\mod_ro_128.fabric[14] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[15].inv  (.Y(\mod_ro_128.fabric[16] ),
    .A(\mod_ro_128.fabric[15] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[16].inv  (.Y(\mod_ro_128.fabric[17] ),
    .A(\mod_ro_128.fabric[16] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[17].inv  (.Y(\mod_ro_128.fabric[18] ),
    .A(\mod_ro_128.fabric[17] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[18].inv  (.Y(\mod_ro_128.fabric[19] ),
    .A(\mod_ro_128.fabric[18] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[19].inv  (.Y(\mod_ro_128.fabric[20] ),
    .A(\mod_ro_128.fabric[19] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[1].inv  (.Y(\mod_ro_128.fabric[2] ),
    .A(\mod_ro_128.fabric[1] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[20].inv  (.Y(\mod_ro_128.fabric[21] ),
    .A(\mod_ro_128.fabric[20] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[21].inv  (.Y(\mod_ro_128.fabric[22] ),
    .A(\mod_ro_128.fabric[21] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[22].inv  (.Y(\mod_ro_128.fabric[23] ),
    .A(\mod_ro_128.fabric[22] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[23].inv  (.Y(\mod_ro_128.fabric[24] ),
    .A(\mod_ro_128.fabric[23] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[24].inv  (.Y(\mod_ro_128.fabric[25] ),
    .A(\mod_ro_128.fabric[24] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[25].inv  (.Y(\mod_ro_128.fabric[26] ),
    .A(\mod_ro_128.fabric[25] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[26].inv  (.Y(\mod_ro_128.fabric[27] ),
    .A(\mod_ro_128.fabric[26] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[27].inv  (.Y(\mod_ro_128.fabric[28] ),
    .A(\mod_ro_128.fabric[27] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[28].inv  (.Y(\mod_ro_128.fabric[29] ),
    .A(\mod_ro_128.fabric[28] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[29].inv  (.Y(\mod_ro_128.fabric[30] ),
    .A(\mod_ro_128.fabric[29] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[2].inv  (.Y(\mod_ro_128.fabric[3] ),
    .A(\mod_ro_128.fabric[2] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[30].inv  (.Y(\mod_ro_128.fabric[31] ),
    .A(\mod_ro_128.fabric[30] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[31].inv  (.Y(\mod_ro_128.fabric[32] ),
    .A(\mod_ro_128.fabric[31] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[32].inv  (.Y(\mod_ro_128.fabric[33] ),
    .A(\mod_ro_128.fabric[32] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[33].inv  (.Y(\mod_ro_128.fabric[34] ),
    .A(\mod_ro_128.fabric[33] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[34].inv  (.Y(\mod_ro_128.fabric[35] ),
    .A(\mod_ro_128.fabric[34] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[35].inv  (.Y(\mod_ro_128.fabric[36] ),
    .A(\mod_ro_128.fabric[35] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[36].inv  (.Y(\mod_ro_128.fabric[37] ),
    .A(\mod_ro_128.fabric[36] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[37].inv  (.Y(\mod_ro_128.fabric[38] ),
    .A(\mod_ro_128.fabric[37] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[38].inv  (.Y(\mod_ro_128.fabric[39] ),
    .A(\mod_ro_128.fabric[38] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[39].inv  (.Y(\mod_ro_128.fabric[40] ),
    .A(\mod_ro_128.fabric[39] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[3].inv  (.Y(\mod_ro_128.fabric[4] ),
    .A(\mod_ro_128.fabric[3] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[40].inv  (.Y(\mod_ro_128.fabric[41] ),
    .A(\mod_ro_128.fabric[40] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[41].inv  (.Y(\mod_ro_128.fabric[42] ),
    .A(\mod_ro_128.fabric[41] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[42].inv  (.Y(\mod_ro_128.fabric[43] ),
    .A(\mod_ro_128.fabric[42] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[43].inv  (.Y(\mod_ro_128.fabric[44] ),
    .A(\mod_ro_128.fabric[43] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[44].inv  (.Y(\mod_ro_128.fabric[45] ),
    .A(\mod_ro_128.fabric[44] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[45].inv  (.Y(\mod_ro_128.fabric[46] ),
    .A(\mod_ro_128.fabric[45] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[46].inv  (.Y(\mod_ro_128.fabric[47] ),
    .A(\mod_ro_128.fabric[46] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[47].inv  (.Y(\mod_ro_128.fabric[48] ),
    .A(\mod_ro_128.fabric[47] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[48].inv  (.Y(\mod_ro_128.fabric[49] ),
    .A(\mod_ro_128.fabric[48] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[49].inv  (.Y(\mod_ro_128.fabric[50] ),
    .A(\mod_ro_128.fabric[49] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[4].inv  (.Y(\mod_ro_128.fabric[5] ),
    .A(\mod_ro_128.fabric[4] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[50].inv  (.Y(\mod_ro_128.fabric[51] ),
    .A(\mod_ro_128.fabric[50] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[51].inv  (.Y(\mod_ro_128.fabric[52] ),
    .A(\mod_ro_128.fabric[51] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[52].inv  (.Y(\mod_ro_128.fabric[53] ),
    .A(\mod_ro_128.fabric[52] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[53].inv  (.Y(\mod_ro_128.fabric[54] ),
    .A(\mod_ro_128.fabric[53] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[54].inv  (.Y(\mod_ro_128.fabric[55] ),
    .A(\mod_ro_128.fabric[54] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[55].inv  (.Y(\mod_ro_128.fabric[56] ),
    .A(\mod_ro_128.fabric[55] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[56].inv  (.Y(\mod_ro_128.fabric[57] ),
    .A(\mod_ro_128.fabric[56] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[57].inv  (.Y(\mod_ro_128.fabric[58] ),
    .A(\mod_ro_128.fabric[57] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[58].inv  (.Y(\mod_ro_128.fabric[59] ),
    .A(\mod_ro_128.fabric[58] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[59].inv  (.Y(\mod_ro_128.fabric[60] ),
    .A(\mod_ro_128.fabric[59] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[5].inv  (.Y(\mod_ro_128.fabric[6] ),
    .A(\mod_ro_128.fabric[5] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[60].inv  (.Y(\mod_ro_128.fabric[61] ),
    .A(\mod_ro_128.fabric[60] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[61].inv  (.Y(\mod_ro_128.fabric[62] ),
    .A(\mod_ro_128.fabric[61] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[62].inv  (.Y(\mod_ro_128.fabric[63] ),
    .A(\mod_ro_128.fabric[62] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[63].inv  (.Y(\mod_ro_128.fabric[64] ),
    .A(\mod_ro_128.fabric[63] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[64].inv  (.Y(\mod_ro_128.fabric[65] ),
    .A(\mod_ro_128.fabric[64] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[65].inv  (.Y(\mod_ro_128.fabric[66] ),
    .A(\mod_ro_128.fabric[65] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[66].inv  (.Y(\mod_ro_128.fabric[67] ),
    .A(\mod_ro_128.fabric[66] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[67].inv  (.Y(\mod_ro_128.fabric[68] ),
    .A(\mod_ro_128.fabric[67] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[68].inv  (.Y(\mod_ro_128.fabric[69] ),
    .A(\mod_ro_128.fabric[68] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[69].inv  (.Y(\mod_ro_128.fabric[70] ),
    .A(\mod_ro_128.fabric[69] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[6].inv  (.Y(\mod_ro_128.fabric[7] ),
    .A(\mod_ro_128.fabric[6] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[70].inv  (.Y(\mod_ro_128.fabric[71] ),
    .A(\mod_ro_128.fabric[70] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[71].inv  (.Y(\mod_ro_128.fabric[72] ),
    .A(\mod_ro_128.fabric[71] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[72].inv  (.Y(\mod_ro_128.fabric[73] ),
    .A(\mod_ro_128.fabric[72] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[73].inv  (.Y(\mod_ro_128.fabric[74] ),
    .A(\mod_ro_128.fabric[73] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[74].inv  (.Y(\mod_ro_128.fabric[75] ),
    .A(\mod_ro_128.fabric[74] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[75].inv  (.Y(\mod_ro_128.fabric[76] ),
    .A(\mod_ro_128.fabric[75] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[76].inv  (.Y(\mod_ro_128.fabric[77] ),
    .A(\mod_ro_128.fabric[76] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[77].inv  (.Y(\mod_ro_128.fabric[78] ),
    .A(\mod_ro_128.fabric[77] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[78].inv  (.Y(\mod_ro_128.fabric[79] ),
    .A(\mod_ro_128.fabric[78] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[79].inv  (.Y(\mod_ro_128.fabric[80] ),
    .A(\mod_ro_128.fabric[79] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[7].inv  (.Y(\mod_ro_128.fabric[8] ),
    .A(\mod_ro_128.fabric[7] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[80].inv  (.Y(\mod_ro_128.fabric[81] ),
    .A(\mod_ro_128.fabric[80] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[81].inv  (.Y(\mod_ro_128.fabric[82] ),
    .A(\mod_ro_128.fabric[81] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[82].inv  (.Y(\mod_ro_128.fabric[83] ),
    .A(\mod_ro_128.fabric[82] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[83].inv  (.Y(\mod_ro_128.fabric[84] ),
    .A(\mod_ro_128.fabric[83] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[84].inv  (.Y(\mod_ro_128.fabric[85] ),
    .A(\mod_ro_128.fabric[84] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[85].inv  (.Y(\mod_ro_128.fabric[86] ),
    .A(\mod_ro_128.fabric[85] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[86].inv  (.Y(\mod_ro_128.fabric[87] ),
    .A(\mod_ro_128.fabric[86] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[87].inv  (.Y(\mod_ro_128.fabric[88] ),
    .A(\mod_ro_128.fabric[87] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[88].inv  (.Y(\mod_ro_128.fabric[89] ),
    .A(\mod_ro_128.fabric[88] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[89].inv  (.Y(\mod_ro_128.fabric[90] ),
    .A(\mod_ro_128.fabric[89] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[8].inv  (.Y(\mod_ro_128.fabric[9] ),
    .A(\mod_ro_128.fabric[8] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[90].inv  (.Y(\mod_ro_128.fabric[91] ),
    .A(\mod_ro_128.fabric[90] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[91].inv  (.Y(\mod_ro_128.fabric[92] ),
    .A(\mod_ro_128.fabric[91] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[92].inv  (.Y(\mod_ro_128.fabric[93] ),
    .A(\mod_ro_128.fabric[92] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[93].inv  (.Y(\mod_ro_128.fabric[94] ),
    .A(\mod_ro_128.fabric[93] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[94].inv  (.Y(\mod_ro_128.fabric[95] ),
    .A(\mod_ro_128.fabric[94] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[95].inv  (.Y(\mod_ro_128.fabric[96] ),
    .A(\mod_ro_128.fabric[95] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[96].inv  (.Y(\mod_ro_128.fabric[97] ),
    .A(\mod_ro_128.fabric[96] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[97].inv  (.Y(\mod_ro_128.fabric[98] ),
    .A(\mod_ro_128.fabric[97] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[98].inv  (.Y(\mod_ro_128.fabric[99] ),
    .A(\mod_ro_128.fabric[98] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[99].inv  (.Y(\mod_ro_128.fabric[100] ),
    .A(\mod_ro_128.fabric[99] ));
 sg13g2_inv_1 \mod_ro_128.osc_gen[9].inv  (.Y(\mod_ro_128.fabric[10] ),
    .A(\mod_ro_128.fabric[9] ));
 sg13g2_inv_1 \mod_ro_16.feedback  (.Y(\mod_ro_16.fabric[0] ),
    .A(\mod_ro_16.fabric[16] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[0].inv  (.Y(\mod_ro_16.fabric[1] ),
    .A(\mod_ro_16.fabric[0] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[10].inv  (.Y(\mod_ro_16.fabric[11] ),
    .A(\mod_ro_16.fabric[10] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[11].inv  (.Y(\mod_ro_16.fabric[12] ),
    .A(\mod_ro_16.fabric[11] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[12].inv  (.Y(\mod_ro_16.fabric[13] ),
    .A(\mod_ro_16.fabric[12] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[13].inv  (.Y(\mod_ro_16.fabric[14] ),
    .A(\mod_ro_16.fabric[13] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[14].inv  (.Y(\mod_ro_16.fabric[15] ),
    .A(\mod_ro_16.fabric[14] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[15].inv  (.Y(\mod_ro_16.fabric[16] ),
    .A(\mod_ro_16.fabric[15] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[1].inv  (.Y(\mod_ro_16.fabric[2] ),
    .A(\mod_ro_16.fabric[1] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[2].inv  (.Y(\mod_ro_16.fabric[3] ),
    .A(\mod_ro_16.fabric[2] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[3].inv  (.Y(\mod_ro_16.fabric[4] ),
    .A(\mod_ro_16.fabric[3] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[4].inv  (.Y(\mod_ro_16.fabric[5] ),
    .A(\mod_ro_16.fabric[4] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[5].inv  (.Y(\mod_ro_16.fabric[6] ),
    .A(\mod_ro_16.fabric[5] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[6].inv  (.Y(\mod_ro_16.fabric[7] ),
    .A(\mod_ro_16.fabric[6] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[7].inv  (.Y(\mod_ro_16.fabric[8] ),
    .A(\mod_ro_16.fabric[7] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[8].inv  (.Y(\mod_ro_16.fabric[9] ),
    .A(\mod_ro_16.fabric[8] ));
 sg13g2_inv_1 \mod_ro_16.osc_gen[9].inv  (.Y(\mod_ro_16.fabric[10] ),
    .A(\mod_ro_16.fabric[9] ));
 sg13g2_inv_1 \mod_ro_256.feedback  (.Y(\mod_ro_256.fabric[0] ),
    .A(\mod_ro_256.fabric[256] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[0].inv  (.Y(\mod_ro_256.fabric[1] ),
    .A(\mod_ro_256.fabric[0] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[100].inv  (.Y(\mod_ro_256.fabric[101] ),
    .A(\mod_ro_256.fabric[100] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[101].inv  (.Y(\mod_ro_256.fabric[102] ),
    .A(\mod_ro_256.fabric[101] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[102].inv  (.Y(\mod_ro_256.fabric[103] ),
    .A(\mod_ro_256.fabric[102] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[103].inv  (.Y(\mod_ro_256.fabric[104] ),
    .A(\mod_ro_256.fabric[103] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[104].inv  (.Y(\mod_ro_256.fabric[105] ),
    .A(\mod_ro_256.fabric[104] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[105].inv  (.Y(\mod_ro_256.fabric[106] ),
    .A(\mod_ro_256.fabric[105] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[106].inv  (.Y(\mod_ro_256.fabric[107] ),
    .A(\mod_ro_256.fabric[106] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[107].inv  (.Y(\mod_ro_256.fabric[108] ),
    .A(\mod_ro_256.fabric[107] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[108].inv  (.Y(\mod_ro_256.fabric[109] ),
    .A(\mod_ro_256.fabric[108] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[109].inv  (.Y(\mod_ro_256.fabric[110] ),
    .A(\mod_ro_256.fabric[109] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[10].inv  (.Y(\mod_ro_256.fabric[11] ),
    .A(\mod_ro_256.fabric[10] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[110].inv  (.Y(\mod_ro_256.fabric[111] ),
    .A(\mod_ro_256.fabric[110] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[111].inv  (.Y(\mod_ro_256.fabric[112] ),
    .A(\mod_ro_256.fabric[111] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[112].inv  (.Y(\mod_ro_256.fabric[113] ),
    .A(\mod_ro_256.fabric[112] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[113].inv  (.Y(\mod_ro_256.fabric[114] ),
    .A(\mod_ro_256.fabric[113] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[114].inv  (.Y(\mod_ro_256.fabric[115] ),
    .A(\mod_ro_256.fabric[114] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[115].inv  (.Y(\mod_ro_256.fabric[116] ),
    .A(\mod_ro_256.fabric[115] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[116].inv  (.Y(\mod_ro_256.fabric[117] ),
    .A(\mod_ro_256.fabric[116] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[117].inv  (.Y(\mod_ro_256.fabric[118] ),
    .A(\mod_ro_256.fabric[117] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[118].inv  (.Y(\mod_ro_256.fabric[119] ),
    .A(\mod_ro_256.fabric[118] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[119].inv  (.Y(\mod_ro_256.fabric[120] ),
    .A(\mod_ro_256.fabric[119] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[11].inv  (.Y(\mod_ro_256.fabric[12] ),
    .A(\mod_ro_256.fabric[11] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[120].inv  (.Y(\mod_ro_256.fabric[121] ),
    .A(\mod_ro_256.fabric[120] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[121].inv  (.Y(\mod_ro_256.fabric[122] ),
    .A(\mod_ro_256.fabric[121] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[122].inv  (.Y(\mod_ro_256.fabric[123] ),
    .A(\mod_ro_256.fabric[122] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[123].inv  (.Y(\mod_ro_256.fabric[124] ),
    .A(\mod_ro_256.fabric[123] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[124].inv  (.Y(\mod_ro_256.fabric[125] ),
    .A(\mod_ro_256.fabric[124] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[125].inv  (.Y(\mod_ro_256.fabric[126] ),
    .A(\mod_ro_256.fabric[125] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[126].inv  (.Y(\mod_ro_256.fabric[127] ),
    .A(\mod_ro_256.fabric[126] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[127].inv  (.Y(\mod_ro_256.fabric[128] ),
    .A(\mod_ro_256.fabric[127] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[128].inv  (.Y(\mod_ro_256.fabric[129] ),
    .A(\mod_ro_256.fabric[128] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[129].inv  (.Y(\mod_ro_256.fabric[130] ),
    .A(\mod_ro_256.fabric[129] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[12].inv  (.Y(\mod_ro_256.fabric[13] ),
    .A(\mod_ro_256.fabric[12] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[130].inv  (.Y(\mod_ro_256.fabric[131] ),
    .A(\mod_ro_256.fabric[130] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[131].inv  (.Y(\mod_ro_256.fabric[132] ),
    .A(\mod_ro_256.fabric[131] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[132].inv  (.Y(\mod_ro_256.fabric[133] ),
    .A(\mod_ro_256.fabric[132] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[133].inv  (.Y(\mod_ro_256.fabric[134] ),
    .A(\mod_ro_256.fabric[133] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[134].inv  (.Y(\mod_ro_256.fabric[135] ),
    .A(\mod_ro_256.fabric[134] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[135].inv  (.Y(\mod_ro_256.fabric[136] ),
    .A(\mod_ro_256.fabric[135] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[136].inv  (.Y(\mod_ro_256.fabric[137] ),
    .A(\mod_ro_256.fabric[136] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[137].inv  (.Y(\mod_ro_256.fabric[138] ),
    .A(\mod_ro_256.fabric[137] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[138].inv  (.Y(\mod_ro_256.fabric[139] ),
    .A(\mod_ro_256.fabric[138] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[139].inv  (.Y(\mod_ro_256.fabric[140] ),
    .A(\mod_ro_256.fabric[139] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[13].inv  (.Y(\mod_ro_256.fabric[14] ),
    .A(\mod_ro_256.fabric[13] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[140].inv  (.Y(\mod_ro_256.fabric[141] ),
    .A(\mod_ro_256.fabric[140] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[141].inv  (.Y(\mod_ro_256.fabric[142] ),
    .A(\mod_ro_256.fabric[141] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[142].inv  (.Y(\mod_ro_256.fabric[143] ),
    .A(\mod_ro_256.fabric[142] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[143].inv  (.Y(\mod_ro_256.fabric[144] ),
    .A(\mod_ro_256.fabric[143] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[144].inv  (.Y(\mod_ro_256.fabric[145] ),
    .A(\mod_ro_256.fabric[144] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[145].inv  (.Y(\mod_ro_256.fabric[146] ),
    .A(\mod_ro_256.fabric[145] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[146].inv  (.Y(\mod_ro_256.fabric[147] ),
    .A(\mod_ro_256.fabric[146] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[147].inv  (.Y(\mod_ro_256.fabric[148] ),
    .A(\mod_ro_256.fabric[147] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[148].inv  (.Y(\mod_ro_256.fabric[149] ),
    .A(\mod_ro_256.fabric[148] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[149].inv  (.Y(\mod_ro_256.fabric[150] ),
    .A(\mod_ro_256.fabric[149] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[14].inv  (.Y(\mod_ro_256.fabric[15] ),
    .A(\mod_ro_256.fabric[14] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[150].inv  (.Y(\mod_ro_256.fabric[151] ),
    .A(\mod_ro_256.fabric[150] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[151].inv  (.Y(\mod_ro_256.fabric[152] ),
    .A(\mod_ro_256.fabric[151] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[152].inv  (.Y(\mod_ro_256.fabric[153] ),
    .A(\mod_ro_256.fabric[152] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[153].inv  (.Y(\mod_ro_256.fabric[154] ),
    .A(\mod_ro_256.fabric[153] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[154].inv  (.Y(\mod_ro_256.fabric[155] ),
    .A(\mod_ro_256.fabric[154] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[155].inv  (.Y(\mod_ro_256.fabric[156] ),
    .A(\mod_ro_256.fabric[155] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[156].inv  (.Y(\mod_ro_256.fabric[157] ),
    .A(\mod_ro_256.fabric[156] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[157].inv  (.Y(\mod_ro_256.fabric[158] ),
    .A(\mod_ro_256.fabric[157] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[158].inv  (.Y(\mod_ro_256.fabric[159] ),
    .A(\mod_ro_256.fabric[158] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[159].inv  (.Y(\mod_ro_256.fabric[160] ),
    .A(\mod_ro_256.fabric[159] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[15].inv  (.Y(\mod_ro_256.fabric[16] ),
    .A(\mod_ro_256.fabric[15] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[160].inv  (.Y(\mod_ro_256.fabric[161] ),
    .A(\mod_ro_256.fabric[160] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[161].inv  (.Y(\mod_ro_256.fabric[162] ),
    .A(\mod_ro_256.fabric[161] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[162].inv  (.Y(\mod_ro_256.fabric[163] ),
    .A(\mod_ro_256.fabric[162] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[163].inv  (.Y(\mod_ro_256.fabric[164] ),
    .A(\mod_ro_256.fabric[163] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[164].inv  (.Y(\mod_ro_256.fabric[165] ),
    .A(\mod_ro_256.fabric[164] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[165].inv  (.Y(\mod_ro_256.fabric[166] ),
    .A(\mod_ro_256.fabric[165] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[166].inv  (.Y(\mod_ro_256.fabric[167] ),
    .A(\mod_ro_256.fabric[166] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[167].inv  (.Y(\mod_ro_256.fabric[168] ),
    .A(\mod_ro_256.fabric[167] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[168].inv  (.Y(\mod_ro_256.fabric[169] ),
    .A(\mod_ro_256.fabric[168] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[169].inv  (.Y(\mod_ro_256.fabric[170] ),
    .A(\mod_ro_256.fabric[169] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[16].inv  (.Y(\mod_ro_256.fabric[17] ),
    .A(\mod_ro_256.fabric[16] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[170].inv  (.Y(\mod_ro_256.fabric[171] ),
    .A(\mod_ro_256.fabric[170] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[171].inv  (.Y(\mod_ro_256.fabric[172] ),
    .A(\mod_ro_256.fabric[171] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[172].inv  (.Y(\mod_ro_256.fabric[173] ),
    .A(\mod_ro_256.fabric[172] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[173].inv  (.Y(\mod_ro_256.fabric[174] ),
    .A(\mod_ro_256.fabric[173] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[174].inv  (.Y(\mod_ro_256.fabric[175] ),
    .A(\mod_ro_256.fabric[174] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[175].inv  (.Y(\mod_ro_256.fabric[176] ),
    .A(\mod_ro_256.fabric[175] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[176].inv  (.Y(\mod_ro_256.fabric[177] ),
    .A(\mod_ro_256.fabric[176] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[177].inv  (.Y(\mod_ro_256.fabric[178] ),
    .A(\mod_ro_256.fabric[177] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[178].inv  (.Y(\mod_ro_256.fabric[179] ),
    .A(\mod_ro_256.fabric[178] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[179].inv  (.Y(\mod_ro_256.fabric[180] ),
    .A(\mod_ro_256.fabric[179] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[17].inv  (.Y(\mod_ro_256.fabric[18] ),
    .A(\mod_ro_256.fabric[17] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[180].inv  (.Y(\mod_ro_256.fabric[181] ),
    .A(\mod_ro_256.fabric[180] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[181].inv  (.Y(\mod_ro_256.fabric[182] ),
    .A(\mod_ro_256.fabric[181] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[182].inv  (.Y(\mod_ro_256.fabric[183] ),
    .A(\mod_ro_256.fabric[182] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[183].inv  (.Y(\mod_ro_256.fabric[184] ),
    .A(\mod_ro_256.fabric[183] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[184].inv  (.Y(\mod_ro_256.fabric[185] ),
    .A(\mod_ro_256.fabric[184] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[185].inv  (.Y(\mod_ro_256.fabric[186] ),
    .A(\mod_ro_256.fabric[185] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[186].inv  (.Y(\mod_ro_256.fabric[187] ),
    .A(\mod_ro_256.fabric[186] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[187].inv  (.Y(\mod_ro_256.fabric[188] ),
    .A(\mod_ro_256.fabric[187] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[188].inv  (.Y(\mod_ro_256.fabric[189] ),
    .A(\mod_ro_256.fabric[188] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[189].inv  (.Y(\mod_ro_256.fabric[190] ),
    .A(\mod_ro_256.fabric[189] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[18].inv  (.Y(\mod_ro_256.fabric[19] ),
    .A(\mod_ro_256.fabric[18] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[190].inv  (.Y(\mod_ro_256.fabric[191] ),
    .A(\mod_ro_256.fabric[190] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[191].inv  (.Y(\mod_ro_256.fabric[192] ),
    .A(\mod_ro_256.fabric[191] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[192].inv  (.Y(\mod_ro_256.fabric[193] ),
    .A(\mod_ro_256.fabric[192] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[193].inv  (.Y(\mod_ro_256.fabric[194] ),
    .A(\mod_ro_256.fabric[193] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[194].inv  (.Y(\mod_ro_256.fabric[195] ),
    .A(\mod_ro_256.fabric[194] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[195].inv  (.Y(\mod_ro_256.fabric[196] ),
    .A(\mod_ro_256.fabric[195] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[196].inv  (.Y(\mod_ro_256.fabric[197] ),
    .A(\mod_ro_256.fabric[196] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[197].inv  (.Y(\mod_ro_256.fabric[198] ),
    .A(\mod_ro_256.fabric[197] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[198].inv  (.Y(\mod_ro_256.fabric[199] ),
    .A(\mod_ro_256.fabric[198] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[199].inv  (.Y(\mod_ro_256.fabric[200] ),
    .A(\mod_ro_256.fabric[199] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[19].inv  (.Y(\mod_ro_256.fabric[20] ),
    .A(\mod_ro_256.fabric[19] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[1].inv  (.Y(\mod_ro_256.fabric[2] ),
    .A(\mod_ro_256.fabric[1] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[200].inv  (.Y(\mod_ro_256.fabric[201] ),
    .A(\mod_ro_256.fabric[200] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[201].inv  (.Y(\mod_ro_256.fabric[202] ),
    .A(\mod_ro_256.fabric[201] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[202].inv  (.Y(\mod_ro_256.fabric[203] ),
    .A(\mod_ro_256.fabric[202] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[203].inv  (.Y(\mod_ro_256.fabric[204] ),
    .A(\mod_ro_256.fabric[203] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[204].inv  (.Y(\mod_ro_256.fabric[205] ),
    .A(\mod_ro_256.fabric[204] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[205].inv  (.Y(\mod_ro_256.fabric[206] ),
    .A(\mod_ro_256.fabric[205] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[206].inv  (.Y(\mod_ro_256.fabric[207] ),
    .A(\mod_ro_256.fabric[206] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[207].inv  (.Y(\mod_ro_256.fabric[208] ),
    .A(\mod_ro_256.fabric[207] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[208].inv  (.Y(\mod_ro_256.fabric[209] ),
    .A(\mod_ro_256.fabric[208] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[209].inv  (.Y(\mod_ro_256.fabric[210] ),
    .A(\mod_ro_256.fabric[209] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[20].inv  (.Y(\mod_ro_256.fabric[21] ),
    .A(\mod_ro_256.fabric[20] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[210].inv  (.Y(\mod_ro_256.fabric[211] ),
    .A(\mod_ro_256.fabric[210] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[211].inv  (.Y(\mod_ro_256.fabric[212] ),
    .A(\mod_ro_256.fabric[211] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[212].inv  (.Y(\mod_ro_256.fabric[213] ),
    .A(\mod_ro_256.fabric[212] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[213].inv  (.Y(\mod_ro_256.fabric[214] ),
    .A(\mod_ro_256.fabric[213] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[214].inv  (.Y(\mod_ro_256.fabric[215] ),
    .A(\mod_ro_256.fabric[214] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[215].inv  (.Y(\mod_ro_256.fabric[216] ),
    .A(\mod_ro_256.fabric[215] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[216].inv  (.Y(\mod_ro_256.fabric[217] ),
    .A(\mod_ro_256.fabric[216] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[217].inv  (.Y(\mod_ro_256.fabric[218] ),
    .A(\mod_ro_256.fabric[217] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[218].inv  (.Y(\mod_ro_256.fabric[219] ),
    .A(\mod_ro_256.fabric[218] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[219].inv  (.Y(\mod_ro_256.fabric[220] ),
    .A(\mod_ro_256.fabric[219] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[21].inv  (.Y(\mod_ro_256.fabric[22] ),
    .A(\mod_ro_256.fabric[21] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[220].inv  (.Y(\mod_ro_256.fabric[221] ),
    .A(\mod_ro_256.fabric[220] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[221].inv  (.Y(\mod_ro_256.fabric[222] ),
    .A(\mod_ro_256.fabric[221] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[222].inv  (.Y(\mod_ro_256.fabric[223] ),
    .A(\mod_ro_256.fabric[222] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[223].inv  (.Y(\mod_ro_256.fabric[224] ),
    .A(\mod_ro_256.fabric[223] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[224].inv  (.Y(\mod_ro_256.fabric[225] ),
    .A(\mod_ro_256.fabric[224] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[225].inv  (.Y(\mod_ro_256.fabric[226] ),
    .A(\mod_ro_256.fabric[225] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[226].inv  (.Y(\mod_ro_256.fabric[227] ),
    .A(\mod_ro_256.fabric[226] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[227].inv  (.Y(\mod_ro_256.fabric[228] ),
    .A(\mod_ro_256.fabric[227] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[228].inv  (.Y(\mod_ro_256.fabric[229] ),
    .A(\mod_ro_256.fabric[228] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[229].inv  (.Y(\mod_ro_256.fabric[230] ),
    .A(\mod_ro_256.fabric[229] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[22].inv  (.Y(\mod_ro_256.fabric[23] ),
    .A(\mod_ro_256.fabric[22] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[230].inv  (.Y(\mod_ro_256.fabric[231] ),
    .A(\mod_ro_256.fabric[230] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[231].inv  (.Y(\mod_ro_256.fabric[232] ),
    .A(\mod_ro_256.fabric[231] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[232].inv  (.Y(\mod_ro_256.fabric[233] ),
    .A(\mod_ro_256.fabric[232] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[233].inv  (.Y(\mod_ro_256.fabric[234] ),
    .A(\mod_ro_256.fabric[233] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[234].inv  (.Y(\mod_ro_256.fabric[235] ),
    .A(\mod_ro_256.fabric[234] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[235].inv  (.Y(\mod_ro_256.fabric[236] ),
    .A(\mod_ro_256.fabric[235] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[236].inv  (.Y(\mod_ro_256.fabric[237] ),
    .A(\mod_ro_256.fabric[236] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[237].inv  (.Y(\mod_ro_256.fabric[238] ),
    .A(\mod_ro_256.fabric[237] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[238].inv  (.Y(\mod_ro_256.fabric[239] ),
    .A(\mod_ro_256.fabric[238] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[239].inv  (.Y(\mod_ro_256.fabric[240] ),
    .A(\mod_ro_256.fabric[239] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[23].inv  (.Y(\mod_ro_256.fabric[24] ),
    .A(\mod_ro_256.fabric[23] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[240].inv  (.Y(\mod_ro_256.fabric[241] ),
    .A(\mod_ro_256.fabric[240] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[241].inv  (.Y(\mod_ro_256.fabric[242] ),
    .A(\mod_ro_256.fabric[241] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[242].inv  (.Y(\mod_ro_256.fabric[243] ),
    .A(\mod_ro_256.fabric[242] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[243].inv  (.Y(\mod_ro_256.fabric[244] ),
    .A(\mod_ro_256.fabric[243] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[244].inv  (.Y(\mod_ro_256.fabric[245] ),
    .A(\mod_ro_256.fabric[244] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[245].inv  (.Y(\mod_ro_256.fabric[246] ),
    .A(\mod_ro_256.fabric[245] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[246].inv  (.Y(\mod_ro_256.fabric[247] ),
    .A(\mod_ro_256.fabric[246] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[247].inv  (.Y(\mod_ro_256.fabric[248] ),
    .A(\mod_ro_256.fabric[247] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[248].inv  (.Y(\mod_ro_256.fabric[249] ),
    .A(\mod_ro_256.fabric[248] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[249].inv  (.Y(\mod_ro_256.fabric[250] ),
    .A(\mod_ro_256.fabric[249] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[24].inv  (.Y(\mod_ro_256.fabric[25] ),
    .A(\mod_ro_256.fabric[24] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[250].inv  (.Y(\mod_ro_256.fabric[251] ),
    .A(\mod_ro_256.fabric[250] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[251].inv  (.Y(\mod_ro_256.fabric[252] ),
    .A(\mod_ro_256.fabric[251] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[252].inv  (.Y(\mod_ro_256.fabric[253] ),
    .A(\mod_ro_256.fabric[252] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[253].inv  (.Y(\mod_ro_256.fabric[254] ),
    .A(\mod_ro_256.fabric[253] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[254].inv  (.Y(\mod_ro_256.fabric[255] ),
    .A(\mod_ro_256.fabric[254] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[255].inv  (.Y(\mod_ro_256.fabric[256] ),
    .A(\mod_ro_256.fabric[255] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[25].inv  (.Y(\mod_ro_256.fabric[26] ),
    .A(\mod_ro_256.fabric[25] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[26].inv  (.Y(\mod_ro_256.fabric[27] ),
    .A(\mod_ro_256.fabric[26] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[27].inv  (.Y(\mod_ro_256.fabric[28] ),
    .A(\mod_ro_256.fabric[27] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[28].inv  (.Y(\mod_ro_256.fabric[29] ),
    .A(\mod_ro_256.fabric[28] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[29].inv  (.Y(\mod_ro_256.fabric[30] ),
    .A(\mod_ro_256.fabric[29] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[2].inv  (.Y(\mod_ro_256.fabric[3] ),
    .A(\mod_ro_256.fabric[2] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[30].inv  (.Y(\mod_ro_256.fabric[31] ),
    .A(\mod_ro_256.fabric[30] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[31].inv  (.Y(\mod_ro_256.fabric[32] ),
    .A(\mod_ro_256.fabric[31] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[32].inv  (.Y(\mod_ro_256.fabric[33] ),
    .A(\mod_ro_256.fabric[32] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[33].inv  (.Y(\mod_ro_256.fabric[34] ),
    .A(\mod_ro_256.fabric[33] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[34].inv  (.Y(\mod_ro_256.fabric[35] ),
    .A(\mod_ro_256.fabric[34] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[35].inv  (.Y(\mod_ro_256.fabric[36] ),
    .A(\mod_ro_256.fabric[35] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[36].inv  (.Y(\mod_ro_256.fabric[37] ),
    .A(\mod_ro_256.fabric[36] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[37].inv  (.Y(\mod_ro_256.fabric[38] ),
    .A(\mod_ro_256.fabric[37] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[38].inv  (.Y(\mod_ro_256.fabric[39] ),
    .A(\mod_ro_256.fabric[38] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[39].inv  (.Y(\mod_ro_256.fabric[40] ),
    .A(\mod_ro_256.fabric[39] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[3].inv  (.Y(\mod_ro_256.fabric[4] ),
    .A(\mod_ro_256.fabric[3] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[40].inv  (.Y(\mod_ro_256.fabric[41] ),
    .A(\mod_ro_256.fabric[40] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[41].inv  (.Y(\mod_ro_256.fabric[42] ),
    .A(\mod_ro_256.fabric[41] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[42].inv  (.Y(\mod_ro_256.fabric[43] ),
    .A(\mod_ro_256.fabric[42] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[43].inv  (.Y(\mod_ro_256.fabric[44] ),
    .A(\mod_ro_256.fabric[43] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[44].inv  (.Y(\mod_ro_256.fabric[45] ),
    .A(\mod_ro_256.fabric[44] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[45].inv  (.Y(\mod_ro_256.fabric[46] ),
    .A(\mod_ro_256.fabric[45] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[46].inv  (.Y(\mod_ro_256.fabric[47] ),
    .A(\mod_ro_256.fabric[46] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[47].inv  (.Y(\mod_ro_256.fabric[48] ),
    .A(\mod_ro_256.fabric[47] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[48].inv  (.Y(\mod_ro_256.fabric[49] ),
    .A(\mod_ro_256.fabric[48] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[49].inv  (.Y(\mod_ro_256.fabric[50] ),
    .A(\mod_ro_256.fabric[49] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[4].inv  (.Y(\mod_ro_256.fabric[5] ),
    .A(\mod_ro_256.fabric[4] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[50].inv  (.Y(\mod_ro_256.fabric[51] ),
    .A(\mod_ro_256.fabric[50] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[51].inv  (.Y(\mod_ro_256.fabric[52] ),
    .A(\mod_ro_256.fabric[51] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[52].inv  (.Y(\mod_ro_256.fabric[53] ),
    .A(\mod_ro_256.fabric[52] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[53].inv  (.Y(\mod_ro_256.fabric[54] ),
    .A(\mod_ro_256.fabric[53] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[54].inv  (.Y(\mod_ro_256.fabric[55] ),
    .A(\mod_ro_256.fabric[54] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[55].inv  (.Y(\mod_ro_256.fabric[56] ),
    .A(\mod_ro_256.fabric[55] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[56].inv  (.Y(\mod_ro_256.fabric[57] ),
    .A(\mod_ro_256.fabric[56] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[57].inv  (.Y(\mod_ro_256.fabric[58] ),
    .A(\mod_ro_256.fabric[57] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[58].inv  (.Y(\mod_ro_256.fabric[59] ),
    .A(\mod_ro_256.fabric[58] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[59].inv  (.Y(\mod_ro_256.fabric[60] ),
    .A(\mod_ro_256.fabric[59] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[5].inv  (.Y(\mod_ro_256.fabric[6] ),
    .A(\mod_ro_256.fabric[5] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[60].inv  (.Y(\mod_ro_256.fabric[61] ),
    .A(\mod_ro_256.fabric[60] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[61].inv  (.Y(\mod_ro_256.fabric[62] ),
    .A(\mod_ro_256.fabric[61] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[62].inv  (.Y(\mod_ro_256.fabric[63] ),
    .A(\mod_ro_256.fabric[62] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[63].inv  (.Y(\mod_ro_256.fabric[64] ),
    .A(\mod_ro_256.fabric[63] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[64].inv  (.Y(\mod_ro_256.fabric[65] ),
    .A(\mod_ro_256.fabric[64] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[65].inv  (.Y(\mod_ro_256.fabric[66] ),
    .A(\mod_ro_256.fabric[65] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[66].inv  (.Y(\mod_ro_256.fabric[67] ),
    .A(\mod_ro_256.fabric[66] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[67].inv  (.Y(\mod_ro_256.fabric[68] ),
    .A(\mod_ro_256.fabric[67] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[68].inv  (.Y(\mod_ro_256.fabric[69] ),
    .A(\mod_ro_256.fabric[68] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[69].inv  (.Y(\mod_ro_256.fabric[70] ),
    .A(\mod_ro_256.fabric[69] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[6].inv  (.Y(\mod_ro_256.fabric[7] ),
    .A(\mod_ro_256.fabric[6] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[70].inv  (.Y(\mod_ro_256.fabric[71] ),
    .A(\mod_ro_256.fabric[70] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[71].inv  (.Y(\mod_ro_256.fabric[72] ),
    .A(\mod_ro_256.fabric[71] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[72].inv  (.Y(\mod_ro_256.fabric[73] ),
    .A(\mod_ro_256.fabric[72] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[73].inv  (.Y(\mod_ro_256.fabric[74] ),
    .A(\mod_ro_256.fabric[73] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[74].inv  (.Y(\mod_ro_256.fabric[75] ),
    .A(\mod_ro_256.fabric[74] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[75].inv  (.Y(\mod_ro_256.fabric[76] ),
    .A(\mod_ro_256.fabric[75] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[76].inv  (.Y(\mod_ro_256.fabric[77] ),
    .A(\mod_ro_256.fabric[76] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[77].inv  (.Y(\mod_ro_256.fabric[78] ),
    .A(\mod_ro_256.fabric[77] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[78].inv  (.Y(\mod_ro_256.fabric[79] ),
    .A(\mod_ro_256.fabric[78] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[79].inv  (.Y(\mod_ro_256.fabric[80] ),
    .A(\mod_ro_256.fabric[79] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[7].inv  (.Y(\mod_ro_256.fabric[8] ),
    .A(\mod_ro_256.fabric[7] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[80].inv  (.Y(\mod_ro_256.fabric[81] ),
    .A(\mod_ro_256.fabric[80] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[81].inv  (.Y(\mod_ro_256.fabric[82] ),
    .A(\mod_ro_256.fabric[81] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[82].inv  (.Y(\mod_ro_256.fabric[83] ),
    .A(\mod_ro_256.fabric[82] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[83].inv  (.Y(\mod_ro_256.fabric[84] ),
    .A(\mod_ro_256.fabric[83] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[84].inv  (.Y(\mod_ro_256.fabric[85] ),
    .A(\mod_ro_256.fabric[84] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[85].inv  (.Y(\mod_ro_256.fabric[86] ),
    .A(\mod_ro_256.fabric[85] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[86].inv  (.Y(\mod_ro_256.fabric[87] ),
    .A(\mod_ro_256.fabric[86] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[87].inv  (.Y(\mod_ro_256.fabric[88] ),
    .A(\mod_ro_256.fabric[87] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[88].inv  (.Y(\mod_ro_256.fabric[89] ),
    .A(\mod_ro_256.fabric[88] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[89].inv  (.Y(\mod_ro_256.fabric[90] ),
    .A(\mod_ro_256.fabric[89] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[8].inv  (.Y(\mod_ro_256.fabric[9] ),
    .A(\mod_ro_256.fabric[8] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[90].inv  (.Y(\mod_ro_256.fabric[91] ),
    .A(\mod_ro_256.fabric[90] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[91].inv  (.Y(\mod_ro_256.fabric[92] ),
    .A(\mod_ro_256.fabric[91] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[92].inv  (.Y(\mod_ro_256.fabric[93] ),
    .A(\mod_ro_256.fabric[92] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[93].inv  (.Y(\mod_ro_256.fabric[94] ),
    .A(\mod_ro_256.fabric[93] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[94].inv  (.Y(\mod_ro_256.fabric[95] ),
    .A(\mod_ro_256.fabric[94] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[95].inv  (.Y(\mod_ro_256.fabric[96] ),
    .A(\mod_ro_256.fabric[95] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[96].inv  (.Y(\mod_ro_256.fabric[97] ),
    .A(\mod_ro_256.fabric[96] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[97].inv  (.Y(\mod_ro_256.fabric[98] ),
    .A(\mod_ro_256.fabric[97] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[98].inv  (.Y(\mod_ro_256.fabric[99] ),
    .A(\mod_ro_256.fabric[98] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[99].inv  (.Y(\mod_ro_256.fabric[100] ),
    .A(\mod_ro_256.fabric[99] ));
 sg13g2_inv_1 \mod_ro_256.osc_gen[9].inv  (.Y(\mod_ro_256.fabric[10] ),
    .A(\mod_ro_256.fabric[9] ));
 sg13g2_inv_1 \mod_ro_31.feedback  (.Y(\mod_ro_31.fabric[0] ),
    .A(\mod_ro_31.fabric[31] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[0].inv  (.Y(\mod_ro_31.fabric[1] ),
    .A(\mod_ro_31.fabric[0] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[10].inv  (.Y(\mod_ro_31.fabric[11] ),
    .A(\mod_ro_31.fabric[10] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[11].inv  (.Y(\mod_ro_31.fabric[12] ),
    .A(\mod_ro_31.fabric[11] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[12].inv  (.Y(\mod_ro_31.fabric[13] ),
    .A(\mod_ro_31.fabric[12] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[13].inv  (.Y(\mod_ro_31.fabric[14] ),
    .A(\mod_ro_31.fabric[13] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[14].inv  (.Y(\mod_ro_31.fabric[15] ),
    .A(\mod_ro_31.fabric[14] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[15].inv  (.Y(\mod_ro_31.fabric[16] ),
    .A(\mod_ro_31.fabric[15] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[16].inv  (.Y(\mod_ro_31.fabric[17] ),
    .A(\mod_ro_31.fabric[16] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[17].inv  (.Y(\mod_ro_31.fabric[18] ),
    .A(\mod_ro_31.fabric[17] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[18].inv  (.Y(\mod_ro_31.fabric[19] ),
    .A(\mod_ro_31.fabric[18] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[19].inv  (.Y(\mod_ro_31.fabric[20] ),
    .A(\mod_ro_31.fabric[19] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[1].inv  (.Y(\mod_ro_31.fabric[2] ),
    .A(\mod_ro_31.fabric[1] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[20].inv  (.Y(\mod_ro_31.fabric[21] ),
    .A(\mod_ro_31.fabric[20] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[21].inv  (.Y(\mod_ro_31.fabric[22] ),
    .A(\mod_ro_31.fabric[21] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[22].inv  (.Y(\mod_ro_31.fabric[23] ),
    .A(\mod_ro_31.fabric[22] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[23].inv  (.Y(\mod_ro_31.fabric[24] ),
    .A(\mod_ro_31.fabric[23] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[24].inv  (.Y(\mod_ro_31.fabric[25] ),
    .A(\mod_ro_31.fabric[24] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[25].inv  (.Y(\mod_ro_31.fabric[26] ),
    .A(\mod_ro_31.fabric[25] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[26].inv  (.Y(\mod_ro_31.fabric[27] ),
    .A(\mod_ro_31.fabric[26] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[27].inv  (.Y(\mod_ro_31.fabric[28] ),
    .A(\mod_ro_31.fabric[27] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[28].inv  (.Y(\mod_ro_31.fabric[29] ),
    .A(\mod_ro_31.fabric[28] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[29].inv  (.Y(\mod_ro_31.fabric[30] ),
    .A(\mod_ro_31.fabric[29] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[2].inv  (.Y(\mod_ro_31.fabric[3] ),
    .A(\mod_ro_31.fabric[2] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[30].inv  (.Y(\mod_ro_31.fabric[31] ),
    .A(\mod_ro_31.fabric[30] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[3].inv  (.Y(\mod_ro_31.fabric[4] ),
    .A(\mod_ro_31.fabric[3] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[4].inv  (.Y(\mod_ro_31.fabric[5] ),
    .A(\mod_ro_31.fabric[4] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[5].inv  (.Y(\mod_ro_31.fabric[6] ),
    .A(\mod_ro_31.fabric[5] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[6].inv  (.Y(\mod_ro_31.fabric[7] ),
    .A(\mod_ro_31.fabric[6] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[7].inv  (.Y(\mod_ro_31.fabric[8] ),
    .A(\mod_ro_31.fabric[7] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[8].inv  (.Y(\mod_ro_31.fabric[9] ),
    .A(\mod_ro_31.fabric[8] ));
 sg13g2_inv_1 \mod_ro_31.osc_gen[9].inv  (.Y(\mod_ro_31.fabric[10] ),
    .A(\mod_ro_31.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_1.feedback  (.Y(\mod_ro_32_1.fabric[0] ),
    .A(\mod_ro_32_1.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[0].inv  (.Y(\mod_ro_32_1.fabric[1] ),
    .A(\mod_ro_32_1.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[10].inv  (.Y(\mod_ro_32_1.fabric[11] ),
    .A(\mod_ro_32_1.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[11].inv  (.Y(\mod_ro_32_1.fabric[12] ),
    .A(\mod_ro_32_1.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[12].inv  (.Y(\mod_ro_32_1.fabric[13] ),
    .A(\mod_ro_32_1.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[13].inv  (.Y(\mod_ro_32_1.fabric[14] ),
    .A(\mod_ro_32_1.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[14].inv  (.Y(\mod_ro_32_1.fabric[15] ),
    .A(\mod_ro_32_1.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[15].inv  (.Y(\mod_ro_32_1.fabric[16] ),
    .A(\mod_ro_32_1.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[16].inv  (.Y(\mod_ro_32_1.fabric[17] ),
    .A(\mod_ro_32_1.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[17].inv  (.Y(\mod_ro_32_1.fabric[18] ),
    .A(\mod_ro_32_1.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[18].inv  (.Y(\mod_ro_32_1.fabric[19] ),
    .A(\mod_ro_32_1.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[19].inv  (.Y(\mod_ro_32_1.fabric[20] ),
    .A(\mod_ro_32_1.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[1].inv  (.Y(\mod_ro_32_1.fabric[2] ),
    .A(\mod_ro_32_1.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[20].inv  (.Y(\mod_ro_32_1.fabric[21] ),
    .A(\mod_ro_32_1.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[21].inv  (.Y(\mod_ro_32_1.fabric[22] ),
    .A(\mod_ro_32_1.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[22].inv  (.Y(\mod_ro_32_1.fabric[23] ),
    .A(\mod_ro_32_1.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[23].inv  (.Y(\mod_ro_32_1.fabric[24] ),
    .A(\mod_ro_32_1.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[24].inv  (.Y(\mod_ro_32_1.fabric[25] ),
    .A(\mod_ro_32_1.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[25].inv  (.Y(\mod_ro_32_1.fabric[26] ),
    .A(\mod_ro_32_1.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[26].inv  (.Y(\mod_ro_32_1.fabric[27] ),
    .A(\mod_ro_32_1.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[27].inv  (.Y(\mod_ro_32_1.fabric[28] ),
    .A(\mod_ro_32_1.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[28].inv  (.Y(\mod_ro_32_1.fabric[29] ),
    .A(\mod_ro_32_1.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[29].inv  (.Y(\mod_ro_32_1.fabric[30] ),
    .A(\mod_ro_32_1.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[2].inv  (.Y(\mod_ro_32_1.fabric[3] ),
    .A(\mod_ro_32_1.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[30].inv  (.Y(\mod_ro_32_1.fabric[31] ),
    .A(\mod_ro_32_1.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[31].inv  (.Y(\mod_ro_32_1.fabric[32] ),
    .A(\mod_ro_32_1.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[3].inv  (.Y(\mod_ro_32_1.fabric[4] ),
    .A(\mod_ro_32_1.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[4].inv  (.Y(\mod_ro_32_1.fabric[5] ),
    .A(\mod_ro_32_1.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[5].inv  (.Y(\mod_ro_32_1.fabric[6] ),
    .A(\mod_ro_32_1.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[6].inv  (.Y(\mod_ro_32_1.fabric[7] ),
    .A(\mod_ro_32_1.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[7].inv  (.Y(\mod_ro_32_1.fabric[8] ),
    .A(\mod_ro_32_1.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[8].inv  (.Y(\mod_ro_32_1.fabric[9] ),
    .A(\mod_ro_32_1.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_1.osc_gen[9].inv  (.Y(\mod_ro_32_1.fabric[10] ),
    .A(\mod_ro_32_1.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_2.feedback  (.Y(\mod_ro_32_2.fabric[0] ),
    .A(\mod_ro_32_2.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[0].inv  (.Y(\mod_ro_32_2.fabric[1] ),
    .A(\mod_ro_32_2.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[10].inv  (.Y(\mod_ro_32_2.fabric[11] ),
    .A(\mod_ro_32_2.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[11].inv  (.Y(\mod_ro_32_2.fabric[12] ),
    .A(\mod_ro_32_2.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[12].inv  (.Y(\mod_ro_32_2.fabric[13] ),
    .A(\mod_ro_32_2.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[13].inv  (.Y(\mod_ro_32_2.fabric[14] ),
    .A(\mod_ro_32_2.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[14].inv  (.Y(\mod_ro_32_2.fabric[15] ),
    .A(\mod_ro_32_2.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[15].inv  (.Y(\mod_ro_32_2.fabric[16] ),
    .A(\mod_ro_32_2.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[16].inv  (.Y(\mod_ro_32_2.fabric[17] ),
    .A(\mod_ro_32_2.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[17].inv  (.Y(\mod_ro_32_2.fabric[18] ),
    .A(\mod_ro_32_2.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[18].inv  (.Y(\mod_ro_32_2.fabric[19] ),
    .A(\mod_ro_32_2.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[19].inv  (.Y(\mod_ro_32_2.fabric[20] ),
    .A(\mod_ro_32_2.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[1].inv  (.Y(\mod_ro_32_2.fabric[2] ),
    .A(\mod_ro_32_2.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[20].inv  (.Y(\mod_ro_32_2.fabric[21] ),
    .A(\mod_ro_32_2.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[21].inv  (.Y(\mod_ro_32_2.fabric[22] ),
    .A(\mod_ro_32_2.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[22].inv  (.Y(\mod_ro_32_2.fabric[23] ),
    .A(\mod_ro_32_2.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[23].inv  (.Y(\mod_ro_32_2.fabric[24] ),
    .A(\mod_ro_32_2.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[24].inv  (.Y(\mod_ro_32_2.fabric[25] ),
    .A(\mod_ro_32_2.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[25].inv  (.Y(\mod_ro_32_2.fabric[26] ),
    .A(\mod_ro_32_2.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[26].inv  (.Y(\mod_ro_32_2.fabric[27] ),
    .A(\mod_ro_32_2.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[27].inv  (.Y(\mod_ro_32_2.fabric[28] ),
    .A(\mod_ro_32_2.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[28].inv  (.Y(\mod_ro_32_2.fabric[29] ),
    .A(\mod_ro_32_2.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[29].inv  (.Y(\mod_ro_32_2.fabric[30] ),
    .A(\mod_ro_32_2.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[2].inv  (.Y(\mod_ro_32_2.fabric[3] ),
    .A(\mod_ro_32_2.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[30].inv  (.Y(\mod_ro_32_2.fabric[31] ),
    .A(\mod_ro_32_2.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[31].inv  (.Y(\mod_ro_32_2.fabric[32] ),
    .A(\mod_ro_32_2.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[3].inv  (.Y(\mod_ro_32_2.fabric[4] ),
    .A(\mod_ro_32_2.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[4].inv  (.Y(\mod_ro_32_2.fabric[5] ),
    .A(\mod_ro_32_2.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[5].inv  (.Y(\mod_ro_32_2.fabric[6] ),
    .A(\mod_ro_32_2.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[6].inv  (.Y(\mod_ro_32_2.fabric[7] ),
    .A(\mod_ro_32_2.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[7].inv  (.Y(\mod_ro_32_2.fabric[8] ),
    .A(\mod_ro_32_2.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[8].inv  (.Y(\mod_ro_32_2.fabric[9] ),
    .A(\mod_ro_32_2.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_2.osc_gen[9].inv  (.Y(\mod_ro_32_2.fabric[10] ),
    .A(\mod_ro_32_2.fabric[9] ));
 sg13g2_inv_1 \mod_ro_32_raw.feedback  (.Y(\mod_ro_32_raw.fabric[0] ),
    .A(\mod_ro_32_raw.fabric[32] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[0].inv  (.Y(\mod_ro_32_raw.fabric[1] ),
    .A(\mod_ro_32_raw.fabric[0] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[10].inv  (.Y(\mod_ro_32_raw.fabric[11] ),
    .A(\mod_ro_32_raw.fabric[10] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[11].inv  (.Y(\mod_ro_32_raw.fabric[12] ),
    .A(\mod_ro_32_raw.fabric[11] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[12].inv  (.Y(\mod_ro_32_raw.fabric[13] ),
    .A(\mod_ro_32_raw.fabric[12] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[13].inv  (.Y(\mod_ro_32_raw.fabric[14] ),
    .A(\mod_ro_32_raw.fabric[13] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[14].inv  (.Y(\mod_ro_32_raw.fabric[15] ),
    .A(\mod_ro_32_raw.fabric[14] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[15].inv  (.Y(\mod_ro_32_raw.fabric[16] ),
    .A(\mod_ro_32_raw.fabric[15] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[16].inv  (.Y(\mod_ro_32_raw.fabric[17] ),
    .A(\mod_ro_32_raw.fabric[16] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[17].inv  (.Y(\mod_ro_32_raw.fabric[18] ),
    .A(\mod_ro_32_raw.fabric[17] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[18].inv  (.Y(\mod_ro_32_raw.fabric[19] ),
    .A(\mod_ro_32_raw.fabric[18] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[19].inv  (.Y(\mod_ro_32_raw.fabric[20] ),
    .A(\mod_ro_32_raw.fabric[19] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[1].inv  (.Y(\mod_ro_32_raw.fabric[2] ),
    .A(\mod_ro_32_raw.fabric[1] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[20].inv  (.Y(\mod_ro_32_raw.fabric[21] ),
    .A(\mod_ro_32_raw.fabric[20] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[21].inv  (.Y(\mod_ro_32_raw.fabric[22] ),
    .A(\mod_ro_32_raw.fabric[21] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[22].inv  (.Y(\mod_ro_32_raw.fabric[23] ),
    .A(\mod_ro_32_raw.fabric[22] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[23].inv  (.Y(\mod_ro_32_raw.fabric[24] ),
    .A(\mod_ro_32_raw.fabric[23] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[24].inv  (.Y(\mod_ro_32_raw.fabric[25] ),
    .A(\mod_ro_32_raw.fabric[24] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[25].inv  (.Y(\mod_ro_32_raw.fabric[26] ),
    .A(\mod_ro_32_raw.fabric[25] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[26].inv  (.Y(\mod_ro_32_raw.fabric[27] ),
    .A(\mod_ro_32_raw.fabric[26] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[27].inv  (.Y(\mod_ro_32_raw.fabric[28] ),
    .A(\mod_ro_32_raw.fabric[27] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[28].inv  (.Y(\mod_ro_32_raw.fabric[29] ),
    .A(\mod_ro_32_raw.fabric[28] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[29].inv  (.Y(\mod_ro_32_raw.fabric[30] ),
    .A(\mod_ro_32_raw.fabric[29] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[2].inv  (.Y(\mod_ro_32_raw.fabric[3] ),
    .A(\mod_ro_32_raw.fabric[2] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[30].inv  (.Y(\mod_ro_32_raw.fabric[31] ),
    .A(\mod_ro_32_raw.fabric[30] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[31].inv  (.Y(\mod_ro_32_raw.fabric[32] ),
    .A(\mod_ro_32_raw.fabric[31] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[3].inv  (.Y(\mod_ro_32_raw.fabric[4] ),
    .A(\mod_ro_32_raw.fabric[3] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[4].inv  (.Y(\mod_ro_32_raw.fabric[5] ),
    .A(\mod_ro_32_raw.fabric[4] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[5].inv  (.Y(\mod_ro_32_raw.fabric[6] ),
    .A(\mod_ro_32_raw.fabric[5] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[6].inv  (.Y(\mod_ro_32_raw.fabric[7] ),
    .A(\mod_ro_32_raw.fabric[6] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[7].inv  (.Y(\mod_ro_32_raw.fabric[8] ),
    .A(\mod_ro_32_raw.fabric[7] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[8].inv  (.Y(\mod_ro_32_raw.fabric[9] ),
    .A(\mod_ro_32_raw.fabric[8] ));
 sg13g2_inv_1 \mod_ro_32_raw.osc_gen[9].inv  (.Y(\mod_ro_32_raw.fabric[10] ),
    .A(\mod_ro_32_raw.fabric[9] ));
 sg13g2_inv_1 \mod_ro_64.feedback  (.Y(\mod_ro_64.fabric[0] ),
    .A(\mod_ro_64.fabric[64] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[0].inv  (.Y(\mod_ro_64.fabric[1] ),
    .A(\mod_ro_64.fabric[0] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[10].inv  (.Y(\mod_ro_64.fabric[11] ),
    .A(\mod_ro_64.fabric[10] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[11].inv  (.Y(\mod_ro_64.fabric[12] ),
    .A(\mod_ro_64.fabric[11] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[12].inv  (.Y(\mod_ro_64.fabric[13] ),
    .A(\mod_ro_64.fabric[12] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[13].inv  (.Y(\mod_ro_64.fabric[14] ),
    .A(\mod_ro_64.fabric[13] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[14].inv  (.Y(\mod_ro_64.fabric[15] ),
    .A(\mod_ro_64.fabric[14] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[15].inv  (.Y(\mod_ro_64.fabric[16] ),
    .A(\mod_ro_64.fabric[15] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[16].inv  (.Y(\mod_ro_64.fabric[17] ),
    .A(\mod_ro_64.fabric[16] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[17].inv  (.Y(\mod_ro_64.fabric[18] ),
    .A(\mod_ro_64.fabric[17] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[18].inv  (.Y(\mod_ro_64.fabric[19] ),
    .A(\mod_ro_64.fabric[18] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[19].inv  (.Y(\mod_ro_64.fabric[20] ),
    .A(\mod_ro_64.fabric[19] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[1].inv  (.Y(\mod_ro_64.fabric[2] ),
    .A(\mod_ro_64.fabric[1] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[20].inv  (.Y(\mod_ro_64.fabric[21] ),
    .A(\mod_ro_64.fabric[20] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[21].inv  (.Y(\mod_ro_64.fabric[22] ),
    .A(\mod_ro_64.fabric[21] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[22].inv  (.Y(\mod_ro_64.fabric[23] ),
    .A(\mod_ro_64.fabric[22] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[23].inv  (.Y(\mod_ro_64.fabric[24] ),
    .A(\mod_ro_64.fabric[23] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[24].inv  (.Y(\mod_ro_64.fabric[25] ),
    .A(\mod_ro_64.fabric[24] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[25].inv  (.Y(\mod_ro_64.fabric[26] ),
    .A(\mod_ro_64.fabric[25] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[26].inv  (.Y(\mod_ro_64.fabric[27] ),
    .A(\mod_ro_64.fabric[26] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[27].inv  (.Y(\mod_ro_64.fabric[28] ),
    .A(\mod_ro_64.fabric[27] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[28].inv  (.Y(\mod_ro_64.fabric[29] ),
    .A(\mod_ro_64.fabric[28] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[29].inv  (.Y(\mod_ro_64.fabric[30] ),
    .A(\mod_ro_64.fabric[29] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[2].inv  (.Y(\mod_ro_64.fabric[3] ),
    .A(\mod_ro_64.fabric[2] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[30].inv  (.Y(\mod_ro_64.fabric[31] ),
    .A(\mod_ro_64.fabric[30] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[31].inv  (.Y(\mod_ro_64.fabric[32] ),
    .A(\mod_ro_64.fabric[31] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[32].inv  (.Y(\mod_ro_64.fabric[33] ),
    .A(\mod_ro_64.fabric[32] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[33].inv  (.Y(\mod_ro_64.fabric[34] ),
    .A(\mod_ro_64.fabric[33] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[34].inv  (.Y(\mod_ro_64.fabric[35] ),
    .A(\mod_ro_64.fabric[34] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[35].inv  (.Y(\mod_ro_64.fabric[36] ),
    .A(\mod_ro_64.fabric[35] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[36].inv  (.Y(\mod_ro_64.fabric[37] ),
    .A(\mod_ro_64.fabric[36] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[37].inv  (.Y(\mod_ro_64.fabric[38] ),
    .A(\mod_ro_64.fabric[37] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[38].inv  (.Y(\mod_ro_64.fabric[39] ),
    .A(\mod_ro_64.fabric[38] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[39].inv  (.Y(\mod_ro_64.fabric[40] ),
    .A(\mod_ro_64.fabric[39] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[3].inv  (.Y(\mod_ro_64.fabric[4] ),
    .A(\mod_ro_64.fabric[3] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[40].inv  (.Y(\mod_ro_64.fabric[41] ),
    .A(\mod_ro_64.fabric[40] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[41].inv  (.Y(\mod_ro_64.fabric[42] ),
    .A(\mod_ro_64.fabric[41] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[42].inv  (.Y(\mod_ro_64.fabric[43] ),
    .A(\mod_ro_64.fabric[42] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[43].inv  (.Y(\mod_ro_64.fabric[44] ),
    .A(\mod_ro_64.fabric[43] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[44].inv  (.Y(\mod_ro_64.fabric[45] ),
    .A(\mod_ro_64.fabric[44] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[45].inv  (.Y(\mod_ro_64.fabric[46] ),
    .A(\mod_ro_64.fabric[45] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[46].inv  (.Y(\mod_ro_64.fabric[47] ),
    .A(\mod_ro_64.fabric[46] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[47].inv  (.Y(\mod_ro_64.fabric[48] ),
    .A(\mod_ro_64.fabric[47] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[48].inv  (.Y(\mod_ro_64.fabric[49] ),
    .A(\mod_ro_64.fabric[48] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[49].inv  (.Y(\mod_ro_64.fabric[50] ),
    .A(\mod_ro_64.fabric[49] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[4].inv  (.Y(\mod_ro_64.fabric[5] ),
    .A(\mod_ro_64.fabric[4] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[50].inv  (.Y(\mod_ro_64.fabric[51] ),
    .A(\mod_ro_64.fabric[50] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[51].inv  (.Y(\mod_ro_64.fabric[52] ),
    .A(\mod_ro_64.fabric[51] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[52].inv  (.Y(\mod_ro_64.fabric[53] ),
    .A(\mod_ro_64.fabric[52] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[53].inv  (.Y(\mod_ro_64.fabric[54] ),
    .A(\mod_ro_64.fabric[53] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[54].inv  (.Y(\mod_ro_64.fabric[55] ),
    .A(\mod_ro_64.fabric[54] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[55].inv  (.Y(\mod_ro_64.fabric[56] ),
    .A(\mod_ro_64.fabric[55] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[56].inv  (.Y(\mod_ro_64.fabric[57] ),
    .A(\mod_ro_64.fabric[56] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[57].inv  (.Y(\mod_ro_64.fabric[58] ),
    .A(\mod_ro_64.fabric[57] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[58].inv  (.Y(\mod_ro_64.fabric[59] ),
    .A(\mod_ro_64.fabric[58] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[59].inv  (.Y(\mod_ro_64.fabric[60] ),
    .A(\mod_ro_64.fabric[59] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[5].inv  (.Y(\mod_ro_64.fabric[6] ),
    .A(\mod_ro_64.fabric[5] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[60].inv  (.Y(\mod_ro_64.fabric[61] ),
    .A(\mod_ro_64.fabric[60] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[61].inv  (.Y(\mod_ro_64.fabric[62] ),
    .A(\mod_ro_64.fabric[61] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[62].inv  (.Y(\mod_ro_64.fabric[63] ),
    .A(\mod_ro_64.fabric[62] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[63].inv  (.Y(\mod_ro_64.fabric[64] ),
    .A(\mod_ro_64.fabric[63] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[6].inv  (.Y(\mod_ro_64.fabric[7] ),
    .A(\mod_ro_64.fabric[6] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[7].inv  (.Y(\mod_ro_64.fabric[8] ),
    .A(\mod_ro_64.fabric[7] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[8].inv  (.Y(\mod_ro_64.fabric[9] ),
    .A(\mod_ro_64.fabric[8] ));
 sg13g2_inv_1 \mod_ro_64.osc_gen[9].inv  (.Y(\mod_ro_64.fabric[10] ),
    .A(\mod_ro_64.fabric[9] ));
 sg13g2_buf_8 fanout13 (.A(_029_),
    .X(net13));
 sg13g2_buf_8 fanout14 (.A(net15),
    .X(net14));
 sg13g2_buf_8 fanout15 (.A(\dpll.n_count[5] ),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(net52),
    .X(net16));
 sg13g2_buf_8 fanout17 (.A(rst_n),
    .X(net17));
 sg13g2_buf_1 fanout18 (.A(rst_n),
    .X(net18));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(uio_in[3]),
    .X(net4));
 sg13g2_tielo tt_um_wedgetail_tester_5 (.L_LO(net5));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_0_clk_regs (.A(clk_regs),
    .X(clknet_0_clk_regs));
 sg13g2_buf_8 clkbuf_2_0__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_0__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_2_1__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_1__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_2_2__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_2__leaf_clk_regs));
 sg13g2_buf_8 clkbuf_2_3__f_clk_regs (.A(clknet_0_clk_regs),
    .X(clknet_2_3__leaf_clk_regs));
 sg13g2_inv_1 clkload0 (.A(clknet_2_1__leaf_clk_regs));
 sg13g2_buf_1 clkload1 (.A(clknet_2_2__leaf_clk_regs));
 sg13g2_inv_1 clkload2 (.A(clknet_2_3__leaf_clk_regs));
 sg13g2_dlygate4sd3_1 hold1 (.A(\dpll.id_out ),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold2 (.A(_001_),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold3 (.A(\dpll.id_increment_done ),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold4 (.A(_011_),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold5 (.A(\dpll.id_decrement_done ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold6 (.A(_010_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold7 (.A(\dpll.k_count_borrow ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold8 (.A(_071_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold9 (.A(_020_),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold10 (.A(\dpll.n_count[1] ),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold11 (.A(_099_),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold12 (.A(_002_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold13 (.A(\dpll.k_count_carry ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold14 (.A(_076_),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold15 (.A(_021_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold16 (.A(\dpll.n_count[2] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold17 (.A(_003_),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold18 (.A(\dpll.id_decrement ),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold19 (.A(\dpll.id_increment ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold20 (.A(\dpll.k_count[4] ),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold21 (.A(_016_),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold22 (.A(\dpll.k_count[7] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold23 (.A(_019_),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold24 (.A(\dpll.k_count[6] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold25 (.A(_018_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold26 (.A(\dpll.k_count[5] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold27 (.A(_017_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold28 (.A(\dpll.k_count[0] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold29 (.A(_012_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold30 (.A(\dpll.k_count[1] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold31 (.A(_013_),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold32 (.A(\dpll.n_count[4] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold33 (.A(_107_),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold34 (.A(_006_),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold35 (.A(\dpll.clk_fout ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold36 (.A(_007_),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold37 (.A(\dpll.clk8x_fout ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold38 (.A(\dpll.k_count[2] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold39 (.A(\dpll.k_count[3] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold40 (.A(\dpll.n_count[0] ),
    .X(net91));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_fill_2 FILLER_8_357 ();
 sg13g2_fill_1 FILLER_8_359 ();
 sg13g2_decap_8 FILLER_8_363 ();
 sg13g2_decap_8 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_377 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_decap_8 FILLER_8_391 ();
 sg13g2_decap_8 FILLER_8_398 ();
 sg13g2_decap_4 FILLER_8_405 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_decap_8 FILLER_9_372 ();
 sg13g2_decap_8 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_393 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_fill_2 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_77 ();
 sg13g2_decap_8 FILLER_10_84 ();
 sg13g2_decap_8 FILLER_10_91 ();
 sg13g2_decap_8 FILLER_10_98 ();
 sg13g2_decap_8 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_8 FILLER_10_119 ();
 sg13g2_decap_8 FILLER_10_126 ();
 sg13g2_decap_8 FILLER_10_133 ();
 sg13g2_decap_8 FILLER_10_140 ();
 sg13g2_decap_8 FILLER_10_147 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_8 FILLER_10_161 ();
 sg13g2_decap_8 FILLER_10_168 ();
 sg13g2_decap_8 FILLER_10_175 ();
 sg13g2_decap_8 FILLER_10_182 ();
 sg13g2_decap_8 FILLER_10_189 ();
 sg13g2_decap_8 FILLER_10_196 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_decap_8 FILLER_10_210 ();
 sg13g2_decap_8 FILLER_10_217 ();
 sg13g2_decap_8 FILLER_10_224 ();
 sg13g2_decap_8 FILLER_10_231 ();
 sg13g2_decap_8 FILLER_10_238 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_8 FILLER_10_259 ();
 sg13g2_decap_8 FILLER_10_266 ();
 sg13g2_decap_8 FILLER_10_273 ();
 sg13g2_decap_8 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_287 ();
 sg13g2_decap_8 FILLER_10_294 ();
 sg13g2_decap_8 FILLER_10_301 ();
 sg13g2_decap_8 FILLER_10_308 ();
 sg13g2_decap_4 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_344 ();
 sg13g2_decap_8 FILLER_10_351 ();
 sg13g2_decap_8 FILLER_10_370 ();
 sg13g2_decap_8 FILLER_10_377 ();
 sg13g2_decap_8 FILLER_10_384 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_4 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_fill_2 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_328 ();
 sg13g2_decap_8 FILLER_11_335 ();
 sg13g2_decap_8 FILLER_11_342 ();
 sg13g2_decap_8 FILLER_11_349 ();
 sg13g2_fill_2 FILLER_11_356 ();
 sg13g2_decap_8 FILLER_11_370 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_fill_2 FILLER_11_391 ();
 sg13g2_fill_1 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_8 FILLER_12_56 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_8 FILLER_12_70 ();
 sg13g2_decap_8 FILLER_12_77 ();
 sg13g2_decap_8 FILLER_12_84 ();
 sg13g2_decap_8 FILLER_12_91 ();
 sg13g2_decap_8 FILLER_12_98 ();
 sg13g2_decap_8 FILLER_12_105 ();
 sg13g2_decap_8 FILLER_12_112 ();
 sg13g2_decap_8 FILLER_12_119 ();
 sg13g2_decap_8 FILLER_12_126 ();
 sg13g2_decap_8 FILLER_12_133 ();
 sg13g2_decap_8 FILLER_12_140 ();
 sg13g2_decap_8 FILLER_12_147 ();
 sg13g2_decap_8 FILLER_12_154 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_decap_8 FILLER_12_168 ();
 sg13g2_decap_8 FILLER_12_175 ();
 sg13g2_decap_8 FILLER_12_182 ();
 sg13g2_decap_8 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_196 ();
 sg13g2_decap_8 FILLER_12_203 ();
 sg13g2_decap_8 FILLER_12_210 ();
 sg13g2_decap_8 FILLER_12_217 ();
 sg13g2_decap_8 FILLER_12_224 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_decap_8 FILLER_12_245 ();
 sg13g2_decap_8 FILLER_12_252 ();
 sg13g2_decap_8 FILLER_12_259 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_273 ();
 sg13g2_decap_8 FILLER_12_280 ();
 sg13g2_decap_8 FILLER_12_287 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_308 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_fill_2 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_325 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_fill_2 FILLER_13_353 ();
 sg13g2_fill_1 FILLER_13_355 ();
 sg13g2_fill_2 FILLER_13_362 ();
 sg13g2_fill_1 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_4 FILLER_13_389 ();
 sg13g2_decap_4 FILLER_13_405 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_4 FILLER_14_308 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_328 ();
 sg13g2_decap_4 FILLER_14_335 ();
 sg13g2_fill_1 FILLER_14_360 ();
 sg13g2_fill_1 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_377 ();
 sg13g2_decap_4 FILLER_14_384 ();
 sg13g2_fill_2 FILLER_14_388 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_decap_8 FILLER_15_49 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_8 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_98 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_8 FILLER_15_126 ();
 sg13g2_decap_8 FILLER_15_133 ();
 sg13g2_decap_8 FILLER_15_140 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_8 FILLER_15_154 ();
 sg13g2_decap_8 FILLER_15_161 ();
 sg13g2_decap_8 FILLER_15_168 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_8 FILLER_15_182 ();
 sg13g2_decap_8 FILLER_15_189 ();
 sg13g2_decap_8 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_15_203 ();
 sg13g2_decap_8 FILLER_15_210 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_decap_8 FILLER_15_238 ();
 sg13g2_decap_8 FILLER_15_245 ();
 sg13g2_decap_8 FILLER_15_252 ();
 sg13g2_decap_8 FILLER_15_259 ();
 sg13g2_decap_8 FILLER_15_266 ();
 sg13g2_decap_8 FILLER_15_273 ();
 sg13g2_decap_8 FILLER_15_280 ();
 sg13g2_decap_8 FILLER_15_287 ();
 sg13g2_decap_8 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_301 ();
 sg13g2_decap_4 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_329 ();
 sg13g2_fill_1 FILLER_15_336 ();
 sg13g2_decap_8 FILLER_15_352 ();
 sg13g2_decap_4 FILLER_15_359 ();
 sg13g2_fill_1 FILLER_15_363 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_4 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_402 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_fill_2 FILLER_16_308 ();
 sg13g2_fill_1 FILLER_16_310 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_4 FILLER_16_333 ();
 sg13g2_fill_1 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_353 ();
 sg13g2_decap_4 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_380 ();
 sg13g2_fill_2 FILLER_16_387 ();
 sg13g2_fill_1 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_402 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_2 FILLER_17_286 ();
 sg13g2_decap_8 FILLER_17_306 ();
 sg13g2_fill_2 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_327 ();
 sg13g2_decap_8 FILLER_17_334 ();
 sg13g2_fill_2 FILLER_17_341 ();
 sg13g2_fill_2 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_366 ();
 sg13g2_fill_2 FILLER_17_373 ();
 sg13g2_fill_1 FILLER_17_375 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_4 FILLER_18_266 ();
 sg13g2_decap_4 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_313 ();
 sg13g2_fill_2 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_fill_1 FILLER_18_355 ();
 sg13g2_fill_2 FILLER_18_374 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_decap_8 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_393 ();
 sg13g2_decap_8 FILLER_18_400 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_281 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_4 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_299 ();
 sg13g2_decap_8 FILLER_19_316 ();
 sg13g2_decap_8 FILLER_19_323 ();
 sg13g2_fill_2 FILLER_19_330 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_4 FILLER_19_361 ();
 sg13g2_fill_1 FILLER_19_365 ();
 sg13g2_decap_8 FILLER_19_387 ();
 sg13g2_decap_8 FILLER_19_394 ();
 sg13g2_decap_8 FILLER_19_401 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_49 ();
 sg13g2_decap_8 FILLER_20_56 ();
 sg13g2_decap_8 FILLER_20_63 ();
 sg13g2_decap_8 FILLER_20_70 ();
 sg13g2_decap_8 FILLER_20_77 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_decap_8 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_decap_8 FILLER_20_126 ();
 sg13g2_decap_8 FILLER_20_133 ();
 sg13g2_decap_8 FILLER_20_140 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_8 FILLER_20_182 ();
 sg13g2_decap_8 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_8 FILLER_20_210 ();
 sg13g2_decap_8 FILLER_20_217 ();
 sg13g2_decap_8 FILLER_20_224 ();
 sg13g2_decap_8 FILLER_20_231 ();
 sg13g2_decap_8 FILLER_20_238 ();
 sg13g2_decap_8 FILLER_20_245 ();
 sg13g2_decap_8 FILLER_20_252 ();
 sg13g2_decap_8 FILLER_20_259 ();
 sg13g2_fill_2 FILLER_20_266 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_1 FILLER_20_288 ();
 sg13g2_decap_8 FILLER_20_292 ();
 sg13g2_decap_8 FILLER_20_299 ();
 sg13g2_fill_2 FILLER_20_306 ();
 sg13g2_decap_4 FILLER_20_323 ();
 sg13g2_fill_2 FILLER_20_327 ();
 sg13g2_decap_4 FILLER_20_332 ();
 sg13g2_fill_2 FILLER_20_336 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_4 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_371 ();
 sg13g2_decap_4 FILLER_20_376 ();
 sg13g2_decap_8 FILLER_20_398 ();
 sg13g2_decap_4 FILLER_20_405 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_4 FILLER_21_315 ();
 sg13g2_fill_1 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_4 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_decap_4 FILLER_21_383 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_decap_4 FILLER_21_404 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_8 FILLER_22_35 ();
 sg13g2_decap_8 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_63 ();
 sg13g2_decap_8 FILLER_22_70 ();
 sg13g2_decap_8 FILLER_22_77 ();
 sg13g2_decap_8 FILLER_22_84 ();
 sg13g2_decap_8 FILLER_22_91 ();
 sg13g2_decap_8 FILLER_22_98 ();
 sg13g2_decap_8 FILLER_22_105 ();
 sg13g2_decap_8 FILLER_22_112 ();
 sg13g2_decap_8 FILLER_22_119 ();
 sg13g2_decap_8 FILLER_22_126 ();
 sg13g2_decap_8 FILLER_22_133 ();
 sg13g2_decap_8 FILLER_22_140 ();
 sg13g2_decap_8 FILLER_22_147 ();
 sg13g2_decap_8 FILLER_22_154 ();
 sg13g2_decap_8 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_168 ();
 sg13g2_decap_8 FILLER_22_175 ();
 sg13g2_decap_8 FILLER_22_182 ();
 sg13g2_decap_8 FILLER_22_189 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_217 ();
 sg13g2_decap_8 FILLER_22_224 ();
 sg13g2_decap_8 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_238 ();
 sg13g2_decap_8 FILLER_22_245 ();
 sg13g2_decap_8 FILLER_22_252 ();
 sg13g2_decap_8 FILLER_22_259 ();
 sg13g2_decap_8 FILLER_22_266 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_fill_2 FILLER_22_287 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_308 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_4 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_fill_1 FILLER_22_389 ();
 sg13g2_decap_4 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_4 FILLER_23_287 ();
 sg13g2_fill_2 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_311 ();
 sg13g2_fill_1 FILLER_23_318 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_8 FILLER_23_341 ();
 sg13g2_decap_8 FILLER_23_348 ();
 sg13g2_decap_8 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_362 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_4 FILLER_23_385 ();
 sg13g2_decap_4 FILLER_23_404 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_8 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_42 ();
 sg13g2_decap_8 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_56 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_decap_8 FILLER_24_70 ();
 sg13g2_decap_8 FILLER_24_77 ();
 sg13g2_decap_8 FILLER_24_84 ();
 sg13g2_decap_8 FILLER_24_91 ();
 sg13g2_decap_8 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_105 ();
 sg13g2_decap_8 FILLER_24_112 ();
 sg13g2_decap_8 FILLER_24_119 ();
 sg13g2_decap_8 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_133 ();
 sg13g2_decap_8 FILLER_24_140 ();
 sg13g2_decap_8 FILLER_24_147 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_decap_8 FILLER_24_161 ();
 sg13g2_decap_4 FILLER_24_168 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_fill_2 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_decap_4 FILLER_24_218 ();
 sg13g2_fill_2 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_decap_8 FILLER_24_240 ();
 sg13g2_decap_8 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_254 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_268 ();
 sg13g2_decap_8 FILLER_24_275 ();
 sg13g2_decap_8 FILLER_24_282 ();
 sg13g2_decap_4 FILLER_24_289 ();
 sg13g2_fill_2 FILLER_24_293 ();
 sg13g2_decap_8 FILLER_24_310 ();
 sg13g2_decap_4 FILLER_24_317 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_decap_4 FILLER_24_337 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_387 ();
 sg13g2_decap_4 FILLER_24_404 ();
 sg13g2_fill_1 FILLER_24_408 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_fill_2 FILLER_25_168 ();
 sg13g2_fill_2 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_311 ();
 sg13g2_decap_8 FILLER_25_318 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_4 FILLER_25_350 ();
 sg13g2_decap_4 FILLER_25_366 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_380 ();
 sg13g2_fill_2 FILLER_25_387 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_fill_1 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_4 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_155 ();
 sg13g2_decap_8 FILLER_26_162 ();
 sg13g2_decap_8 FILLER_26_169 ();
 sg13g2_fill_1 FILLER_26_176 ();
 sg13g2_decap_8 FILLER_26_190 ();
 sg13g2_decap_8 FILLER_26_197 ();
 sg13g2_decap_4 FILLER_26_204 ();
 sg13g2_fill_1 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_226 ();
 sg13g2_fill_1 FILLER_26_228 ();
 sg13g2_fill_1 FILLER_26_234 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_281 ();
 sg13g2_decap_8 FILLER_26_288 ();
 sg13g2_decap_8 FILLER_26_313 ();
 sg13g2_decap_4 FILLER_26_320 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_345 ();
 sg13g2_decap_4 FILLER_26_352 ();
 sg13g2_fill_1 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_366 ();
 sg13g2_decap_4 FILLER_26_382 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_4 FILLER_27_140 ();
 sg13g2_fill_2 FILLER_27_144 ();
 sg13g2_fill_2 FILLER_27_174 ();
 sg13g2_fill_1 FILLER_27_176 ();
 sg13g2_fill_2 FILLER_27_185 ();
 sg13g2_fill_1 FILLER_27_187 ();
 sg13g2_decap_4 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_27_202 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_fill_1 FILLER_27_217 ();
 sg13g2_fill_2 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_233 ();
 sg13g2_decap_4 FILLER_27_242 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_fill_2 FILLER_27_259 ();
 sg13g2_fill_1 FILLER_27_266 ();
 sg13g2_decap_4 FILLER_27_295 ();
 sg13g2_fill_2 FILLER_27_320 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_fill_2 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_fill_1 FILLER_27_356 ();
 sg13g2_decap_4 FILLER_27_369 ();
 sg13g2_fill_2 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_4 FILLER_27_403 ();
 sg13g2_fill_2 FILLER_27_407 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_fill_2 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_163 ();
 sg13g2_fill_2 FILLER_28_204 ();
 sg13g2_decap_4 FILLER_28_224 ();
 sg13g2_fill_2 FILLER_28_228 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_fill_1 FILLER_28_244 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_303 ();
 sg13g2_fill_1 FILLER_28_316 ();
 sg13g2_decap_4 FILLER_28_335 ();
 sg13g2_fill_2 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_4 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_370 ();
 sg13g2_decap_4 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_4 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_decap_8 FILLER_29_63 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_decap_8 FILLER_29_126 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_4 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_209 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_fill_2 FILLER_29_223 ();
 sg13g2_fill_1 FILLER_29_225 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_251 ();
 sg13g2_fill_2 FILLER_29_258 ();
 sg13g2_fill_1 FILLER_29_260 ();
 sg13g2_decap_4 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_321 ();
 sg13g2_decap_4 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_332 ();
 sg13g2_decap_8 FILLER_29_352 ();
 sg13g2_fill_2 FILLER_29_359 ();
 sg13g2_fill_1 FILLER_29_361 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_387 ();
 sg13g2_decap_8 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_fill_2 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_160 ();
 sg13g2_decap_4 FILLER_30_167 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_decap_4 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_231 ();
 sg13g2_fill_2 FILLER_30_269 ();
 sg13g2_fill_1 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_fill_2 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_4 FILLER_30_336 ();
 sg13g2_fill_1 FILLER_30_340 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_decap_4 FILLER_30_358 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_4 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_402 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_fill_2 FILLER_31_154 ();
 sg13g2_fill_1 FILLER_31_192 ();
 sg13g2_fill_2 FILLER_31_203 ();
 sg13g2_fill_2 FILLER_31_210 ();
 sg13g2_fill_1 FILLER_31_212 ();
 sg13g2_fill_1 FILLER_31_219 ();
 sg13g2_fill_2 FILLER_31_246 ();
 sg13g2_fill_1 FILLER_31_248 ();
 sg13g2_fill_2 FILLER_31_277 ();
 sg13g2_fill_1 FILLER_31_279 ();
 sg13g2_fill_2 FILLER_31_285 ();
 sg13g2_fill_1 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_fill_2 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_324 ();
 sg13g2_decap_4 FILLER_31_346 ();
 sg13g2_fill_1 FILLER_31_353 ();
 sg13g2_fill_1 FILLER_31_357 ();
 sg13g2_decap_4 FILLER_31_376 ();
 sg13g2_fill_1 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_fill_2 FILLER_31_406 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_42 ();
 sg13g2_decap_8 FILLER_32_49 ();
 sg13g2_decap_8 FILLER_32_56 ();
 sg13g2_decap_8 FILLER_32_63 ();
 sg13g2_decap_8 FILLER_32_70 ();
 sg13g2_decap_8 FILLER_32_77 ();
 sg13g2_decap_8 FILLER_32_84 ();
 sg13g2_decap_8 FILLER_32_91 ();
 sg13g2_decap_8 FILLER_32_98 ();
 sg13g2_decap_8 FILLER_32_105 ();
 sg13g2_decap_8 FILLER_32_112 ();
 sg13g2_decap_8 FILLER_32_119 ();
 sg13g2_decap_8 FILLER_32_126 ();
 sg13g2_decap_8 FILLER_32_133 ();
 sg13g2_decap_8 FILLER_32_140 ();
 sg13g2_decap_8 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_154 ();
 sg13g2_fill_2 FILLER_32_161 ();
 sg13g2_fill_1 FILLER_32_163 ();
 sg13g2_decap_8 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_fill_2 FILLER_32_208 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_267 ();
 sg13g2_fill_2 FILLER_32_273 ();
 sg13g2_fill_1 FILLER_32_275 ();
 sg13g2_decap_8 FILLER_32_317 ();
 sg13g2_decap_8 FILLER_32_324 ();
 sg13g2_fill_2 FILLER_32_331 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_decap_8 FILLER_32_364 ();
 sg13g2_fill_2 FILLER_32_371 ();
 sg13g2_fill_2 FILLER_32_379 ();
 sg13g2_decap_4 FILLER_32_387 ();
 sg13g2_fill_1 FILLER_32_391 ();
 sg13g2_decap_4 FILLER_32_404 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_4 FILLER_33_161 ();
 sg13g2_fill_1 FILLER_33_165 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_fill_2 FILLER_33_213 ();
 sg13g2_fill_1 FILLER_33_215 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_fill_2 FILLER_33_329 ();
 sg13g2_decap_4 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_355 ();
 sg13g2_decap_8 FILLER_33_362 ();
 sg13g2_fill_2 FILLER_33_369 ();
 sg13g2_fill_1 FILLER_33_371 ();
 sg13g2_fill_2 FILLER_33_390 ();
 sg13g2_decap_4 FILLER_33_404 ();
 sg13g2_fill_1 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_105 ();
 sg13g2_decap_8 FILLER_34_112 ();
 sg13g2_decap_8 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_126 ();
 sg13g2_fill_1 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_156 ();
 sg13g2_decap_8 FILLER_34_163 ();
 sg13g2_fill_2 FILLER_34_170 ();
 sg13g2_decap_8 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_192 ();
 sg13g2_fill_2 FILLER_34_206 ();
 sg13g2_fill_2 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_decap_4 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_325 ();
 sg13g2_fill_2 FILLER_34_333 ();
 sg13g2_fill_1 FILLER_34_335 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_fill_2 FILLER_34_356 ();
 sg13g2_fill_1 FILLER_34_358 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_4 FILLER_34_403 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_fill_1 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_142 ();
 sg13g2_fill_1 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_157 ();
 sg13g2_decap_8 FILLER_35_164 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_fill_1 FILLER_35_227 ();
 sg13g2_decap_8 FILLER_35_236 ();
 sg13g2_decap_8 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_2 FILLER_35_257 ();
 sg13g2_fill_1 FILLER_35_259 ();
 sg13g2_decap_4 FILLER_35_310 ();
 sg13g2_fill_2 FILLER_35_314 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_decap_4 FILLER_35_338 ();
 sg13g2_fill_1 FILLER_35_342 ();
 sg13g2_decap_8 FILLER_35_353 ();
 sg13g2_decap_4 FILLER_35_360 ();
 sg13g2_fill_1 FILLER_35_364 ();
 sg13g2_fill_2 FILLER_35_374 ();
 sg13g2_fill_1 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_119 ();
 sg13g2_fill_1 FILLER_36_121 ();
 sg13g2_fill_1 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_135 ();
 sg13g2_fill_2 FILLER_36_142 ();
 sg13g2_decap_4 FILLER_36_156 ();
 sg13g2_fill_1 FILLER_36_160 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_fill_2 FILLER_36_189 ();
 sg13g2_fill_1 FILLER_36_191 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_decap_4 FILLER_36_234 ();
 sg13g2_fill_1 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_296 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_330 ();
 sg13g2_fill_2 FILLER_36_337 ();
 sg13g2_fill_2 FILLER_36_345 ();
 sg13g2_fill_1 FILLER_36_347 ();
 sg13g2_decap_4 FILLER_36_366 ();
 sg13g2_fill_1 FILLER_36_370 ();
 sg13g2_fill_1 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_381 ();
 sg13g2_decap_4 FILLER_36_388 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_146 ();
 sg13g2_decap_8 FILLER_37_153 ();
 sg13g2_decap_4 FILLER_37_160 ();
 sg13g2_fill_1 FILLER_37_164 ();
 sg13g2_decap_4 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_209 ();
 sg13g2_fill_2 FILLER_37_221 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_decap_8 FILLER_37_345 ();
 sg13g2_decap_8 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_380 ();
 sg13g2_fill_1 FILLER_37_382 ();
 sg13g2_fill_2 FILLER_37_386 ();
 sg13g2_fill_1 FILLER_37_391 ();
 sg13g2_decap_4 FILLER_37_404 ();
 sg13g2_fill_1 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_4 FILLER_38_60 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_decap_4 FILLER_38_76 ();
 sg13g2_decap_4 FILLER_38_84 ();
 sg13g2_decap_4 FILLER_38_92 ();
 sg13g2_decap_4 FILLER_38_100 ();
 sg13g2_decap_4 FILLER_38_108 ();
 sg13g2_decap_4 FILLER_38_116 ();
 sg13g2_decap_4 FILLER_38_124 ();
 sg13g2_fill_1 FILLER_38_132 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_decap_4 FILLER_38_148 ();
 sg13g2_decap_4 FILLER_38_156 ();
 sg13g2_decap_4 FILLER_38_164 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_fill_2 FILLER_38_180 ();
 sg13g2_fill_1 FILLER_38_182 ();
 sg13g2_fill_1 FILLER_38_191 ();
 sg13g2_decap_4 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_204 ();
 sg13g2_fill_2 FILLER_38_220 ();
 sg13g2_fill_1 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_292 ();
 sg13g2_decap_4 FILLER_38_327 ();
 sg13g2_fill_2 FILLER_38_331 ();
 sg13g2_fill_1 FILLER_38_351 ();
 sg13g2_fill_1 FILLER_38_367 ();
 sg13g2_decap_4 FILLER_38_387 ();
 sg13g2_fill_1 FILLER_38_391 ();
 sg13g2_decap_4 FILLER_38_404 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net5;
 assign uio_oe[1] = net6;
 assign uio_oe[2] = net7;
 assign uio_oe[3] = net8;
 assign uio_oe[4] = net9;
 assign uio_oe[5] = net10;
 assign uio_oe[6] = net11;
 assign uio_oe[7] = net12;
 assign uio_out[0] = net19;
 assign uio_out[1] = net20;
 assign uio_out[2] = net21;
 assign uio_out[3] = net22;
 assign uio_out[4] = net23;
 assign uio_out[5] = net24;
 assign uio_out[6] = net25;
 assign uio_out[7] = net26;
 assign uo_out[5] = net27;
 assign uo_out[6] = net28;
 assign uo_out[7] = net29;
endmodule
