module tt_um_posit_mac_stream (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire \u_mac.u_adder.sign_b ;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;

 sg13g2_inv_1 _1093_ (.Y(_0367_),
    .A(net3));
 sg13g2_inv_1 _1094_ (.Y(_0378_),
    .A(net11));
 sg13g2_inv_1 _1095_ (.Y(_0389_),
    .A(net17));
 sg13g2_inv_4 _1096_ (.A(\u_mac.u_adder.sign_b ),
    .Y(_0400_));
 sg13g2_inv_1 _1097_ (.Y(_0411_),
    .A(net35));
 sg13g2_inv_1 _1098_ (.Y(_0422_),
    .A(net41));
 sg13g2_inv_1 _1099_ (.Y(_0433_),
    .A(net42));
 sg13g2_inv_1 _1100_ (.Y(_0444_),
    .A(net34));
 sg13g2_inv_1 _1101_ (.Y(_0455_),
    .A(net36));
 sg13g2_inv_2 _1102_ (.Y(_0466_),
    .A(net39));
 sg13g2_nor3_1 _1103_ (.A(net4),
    .B(net3),
    .C(net5),
    .Y(_0477_));
 sg13g2_or4_1 _1104_ (.A(net4),
    .B(net3),
    .C(net6),
    .D(net5),
    .X(_0488_));
 sg13g2_or2_1 _1105_ (.X(_0499_),
    .B(net7),
    .A(net8));
 sg13g2_nor3_2 _1106_ (.A(net9),
    .B(_0488_),
    .C(_0499_),
    .Y(_0510_));
 sg13g2_or3_1 _1107_ (.A(net9),
    .B(_0488_),
    .C(_0499_),
    .X(_0521_));
 sg13g2_nor3_1 _1108_ (.A(net12),
    .B(net11),
    .C(net13),
    .Y(_0532_));
 sg13g2_or4_1 _1109_ (.A(net12),
    .B(net11),
    .C(net14),
    .D(net13),
    .X(_0543_));
 sg13g2_or3_1 _1110_ (.A(net16),
    .B(net15),
    .C(_0543_),
    .X(_0554_));
 sg13g2_nor2_2 _1111_ (.A(net17),
    .B(_0554_),
    .Y(_0565_));
 sg13g2_nand2b_2 _1112_ (.Y(_0576_),
    .B(_0389_),
    .A_N(_0554_));
 sg13g2_nor2_2 _1113_ (.A(_0510_),
    .B(_0565_),
    .Y(_0587_));
 sg13g2_nand2_1 _1114_ (.Y(_0598_),
    .A(_0521_),
    .B(_0576_));
 sg13g2_a22oi_1 _1115_ (.Y(_0609_),
    .B1(_0565_),
    .B2(net104),
    .A2(_0510_),
    .A1(net105));
 sg13g2_nand2_1 _1116_ (.Y(_0620_),
    .A(net98),
    .B(_0609_));
 sg13g2_nand2_2 _1117_ (.Y(_0631_),
    .A(net1),
    .B(_0620_));
 sg13g2_o21ai_1 _1118_ (.B1(net105),
    .Y(_0642_),
    .A1(_0488_),
    .A2(_0499_));
 sg13g2_xor2_1 _1119_ (.B(_0642_),
    .A(net9),
    .X(_0653_));
 sg13g2_nand3_1 _1120_ (.B(net102),
    .C(_0554_),
    .A(_0389_),
    .Y(_0664_));
 sg13g2_a21o_1 _1121_ (.A2(_0554_),
    .A1(net102),
    .B1(_0389_),
    .X(_0675_));
 sg13g2_a21oi_2 _1122_ (.B1(net17),
    .Y(_0686_),
    .A2(_0554_),
    .A1(net103));
 sg13g2_a21o_2 _1123_ (.A2(_0554_),
    .A1(net103),
    .B1(net17),
    .X(_0697_));
 sg13g2_and3_2 _1124_ (.X(_0708_),
    .A(net17),
    .B(net102),
    .C(_0554_));
 sg13g2_nand3_1 _1125_ (.B(net103),
    .C(_0554_),
    .A(net17),
    .Y(_0719_));
 sg13g2_nand2_2 _1126_ (.Y(_0730_),
    .A(_0697_),
    .B(_0719_));
 sg13g2_and4_1 _1127_ (.A(_0521_),
    .B(_0576_),
    .C(net101),
    .D(_0730_),
    .X(_0741_));
 sg13g2_inv_1 _1128_ (.Y(_0752_),
    .A(_0741_));
 sg13g2_nand2_1 _1129_ (.Y(_0763_),
    .A(net105),
    .B(_0488_));
 sg13g2_xor2_1 _1130_ (.B(_0763_),
    .A(net7),
    .X(_0774_));
 sg13g2_xnor2_1 _1131_ (.Y(_0785_),
    .A(net100),
    .B(_0774_));
 sg13g2_inv_1 _1132_ (.Y(_0796_),
    .A(_0785_));
 sg13g2_nor2b_1 _1133_ (.A(_0477_),
    .B_N(net105),
    .Y(_0807_));
 sg13g2_xnor2_1 _1134_ (.Y(_0818_),
    .A(net6),
    .B(_0807_));
 sg13g2_xnor2_1 _1135_ (.Y(_0829_),
    .A(net100),
    .B(_0818_));
 sg13g2_and2_1 _1136_ (.A(_0785_),
    .B(_0829_),
    .X(_0840_));
 sg13g2_o21ai_1 _1137_ (.B1(net105),
    .Y(_0851_),
    .A1(net7),
    .A2(_0488_));
 sg13g2_xnor2_1 _1138_ (.Y(_0862_),
    .A(net8),
    .B(_0851_));
 sg13g2_xor2_1 _1139_ (.B(_0862_),
    .A(net100),
    .X(_0873_));
 sg13g2_xnor2_1 _1140_ (.Y(_0884_),
    .A(net100),
    .B(_0862_));
 sg13g2_nand2_2 _1141_ (.Y(_0895_),
    .A(_0840_),
    .B(_0873_));
 sg13g2_o21ai_1 _1142_ (.B1(net105),
    .Y(_0906_),
    .A1(net4),
    .A2(net3));
 sg13g2_xnor2_1 _1143_ (.Y(_0917_),
    .A(net5),
    .B(_0906_));
 sg13g2_inv_2 _1144_ (.Y(_0928_),
    .A(_0917_));
 sg13g2_nand2_1 _1145_ (.Y(_0939_),
    .A(net101),
    .B(_0895_));
 sg13g2_o21ai_1 _1146_ (.B1(_0939_),
    .Y(_0950_),
    .A1(_0895_),
    .A2(_0928_));
 sg13g2_nand2_1 _1147_ (.Y(_0961_),
    .A(net102),
    .B(_0543_));
 sg13g2_xor2_1 _1148_ (.B(_0961_),
    .A(net15),
    .X(_0972_));
 sg13g2_nand3_1 _1149_ (.B(_0719_),
    .C(_0972_),
    .A(_0697_),
    .Y(_0983_));
 sg13g2_a21o_1 _1150_ (.A2(_0719_),
    .A1(_0697_),
    .B1(_0972_),
    .X(_0994_));
 sg13g2_nand2_1 _1151_ (.Y(_1005_),
    .A(_0983_),
    .B(_0994_));
 sg13g2_nand2b_1 _1152_ (.Y(_1016_),
    .B(net102),
    .A_N(_0532_));
 sg13g2_xnor2_1 _1153_ (.Y(_1027_),
    .A(net14),
    .B(_1016_));
 sg13g2_or3_1 _1154_ (.A(_0686_),
    .B(_0708_),
    .C(_1027_),
    .X(_1038_));
 sg13g2_o21ai_1 _1155_ (.B1(_1027_),
    .Y(_1049_),
    .A1(_0686_),
    .A2(_0708_));
 sg13g2_and2_1 _1156_ (.A(_1038_),
    .B(_1049_),
    .X(_1060_));
 sg13g2_nand2_1 _1157_ (.Y(_1071_),
    .A(_1038_),
    .B(_1049_));
 sg13g2_nand4_1 _1158_ (.B(_0994_),
    .C(_1038_),
    .A(_0983_),
    .Y(_1082_),
    .D(_1049_));
 sg13g2_o21ai_1 _1159_ (.B1(net102),
    .Y(_0008_),
    .A1(net15),
    .A2(_0543_));
 sg13g2_xor2_1 _1160_ (.B(_0008_),
    .A(net16),
    .X(_0019_));
 sg13g2_xnor2_1 _1161_ (.Y(_0030_),
    .A(_0730_),
    .B(_0019_));
 sg13g2_xor2_1 _1162_ (.B(_0019_),
    .A(_0730_),
    .X(_0041_));
 sg13g2_nand2b_1 _1163_ (.Y(_0052_),
    .B(_0030_),
    .A_N(_1082_));
 sg13g2_o21ai_1 _1164_ (.B1(net102),
    .Y(_0063_),
    .A1(net12),
    .A2(net11));
 sg13g2_xnor2_1 _1165_ (.Y(_0074_),
    .A(net13),
    .B(_0063_));
 sg13g2_inv_2 _1166_ (.Y(_0084_),
    .A(_0074_));
 sg13g2_nand2_1 _1167_ (.Y(_0094_),
    .A(_0730_),
    .B(_0052_));
 sg13g2_o21ai_1 _1168_ (.B1(_0094_),
    .Y(_0104_),
    .A1(_0052_),
    .A2(_0084_));
 sg13g2_and2_1 _1169_ (.A(_0950_),
    .B(_0104_),
    .X(_0114_));
 sg13g2_xnor2_1 _1170_ (.Y(_0124_),
    .A(net100),
    .B(_0928_));
 sg13g2_nand2_1 _1171_ (.Y(_0134_),
    .A(net3),
    .B(net10));
 sg13g2_xor2_1 _1172_ (.B(_0134_),
    .A(net4),
    .X(_0140_));
 sg13g2_xnor2_1 _1173_ (.Y(_0141_),
    .A(net100),
    .B(_0140_));
 sg13g2_nand2_2 _1174_ (.Y(_0142_),
    .A(_0124_),
    .B(_0141_));
 sg13g2_nand3b_1 _1175_ (.B(net4),
    .C(_0367_),
    .Y(_0143_),
    .A_N(net101));
 sg13g2_nand3_1 _1176_ (.B(net101),
    .C(_0140_),
    .A(net3),
    .Y(_0144_));
 sg13g2_nand3_1 _1177_ (.B(_0143_),
    .C(_0144_),
    .A(_0124_),
    .Y(_0145_));
 sg13g2_a21oi_2 _1178_ (.B1(_0796_),
    .Y(_0146_),
    .A2(_0145_),
    .A1(_0829_));
 sg13g2_a21o_2 _1179_ (.A2(_0145_),
    .A1(_0829_),
    .B1(_0796_),
    .X(_0147_));
 sg13g2_a21oi_1 _1180_ (.A1(_0840_),
    .A2(_0142_),
    .Y(_0148_),
    .B1(_0884_));
 sg13g2_nand2_2 _1181_ (.Y(_0149_),
    .A(_0146_),
    .B(_0148_));
 sg13g2_nand2_2 _1182_ (.Y(_0150_),
    .A(_0873_),
    .B(_0147_));
 sg13g2_nand4_1 _1183_ (.B(_0873_),
    .C(_0142_),
    .A(_0840_),
    .Y(_0151_),
    .D(_0147_));
 sg13g2_and2_1 _1184_ (.A(_0149_),
    .B(_0151_),
    .X(_0152_));
 sg13g2_xor2_1 _1185_ (.B(_0152_),
    .A(net100),
    .X(_0153_));
 sg13g2_nand2_1 _1186_ (.Y(_0154_),
    .A(net11),
    .B(net102));
 sg13g2_xor2_1 _1187_ (.B(_0154_),
    .A(net12),
    .X(_0155_));
 sg13g2_xnor2_1 _1188_ (.Y(_0156_),
    .A(net12),
    .B(_0154_));
 sg13g2_nand3_1 _1189_ (.B(_0719_),
    .C(_0156_),
    .A(_0697_),
    .Y(_0157_));
 sg13g2_o21ai_1 _1190_ (.B1(_0155_),
    .Y(_0158_),
    .A1(_0686_),
    .A2(_0708_));
 sg13g2_o21ai_1 _1191_ (.B1(_0074_),
    .Y(_0159_),
    .A1(_0686_),
    .A2(_0708_));
 sg13g2_nand3_1 _1192_ (.B(_0719_),
    .C(_0084_),
    .A(_0697_),
    .Y(_0160_));
 sg13g2_nand3_1 _1193_ (.B(_0719_),
    .C(_0074_),
    .A(_0697_),
    .Y(_0161_));
 sg13g2_o21ai_1 _1194_ (.B1(_0084_),
    .Y(_0162_),
    .A1(_0686_),
    .A2(_0708_));
 sg13g2_a22oi_1 _1195_ (.Y(_0163_),
    .B1(_0161_),
    .B2(_0162_),
    .A2(_0158_),
    .A1(_0157_));
 sg13g2_o21ai_1 _1196_ (.B1(_0030_),
    .Y(_0164_),
    .A1(_1082_),
    .A2(_0163_));
 sg13g2_nand4_1 _1197_ (.B(_0697_),
    .C(_0719_),
    .A(_0378_),
    .Y(_0165_),
    .D(_0156_));
 sg13g2_nand4_1 _1198_ (.B(_0664_),
    .C(_0675_),
    .A(net11),
    .Y(_0166_),
    .D(_0155_));
 sg13g2_nand4_1 _1199_ (.B(_0160_),
    .C(_0165_),
    .A(_0159_),
    .Y(_0167_),
    .D(_0166_));
 sg13g2_a21oi_1 _1200_ (.A1(_1060_),
    .A2(_0167_),
    .Y(_0168_),
    .B1(_1005_));
 sg13g2_a21o_2 _1201_ (.A2(_0167_),
    .A1(_1060_),
    .B1(_1005_),
    .X(_0169_));
 sg13g2_nand2_1 _1202_ (.Y(_0170_),
    .A(_0019_),
    .B(_0169_));
 sg13g2_o21ai_1 _1203_ (.B1(_0170_),
    .Y(_0171_),
    .A1(_0730_),
    .A2(_0169_));
 sg13g2_xnor2_1 _1204_ (.Y(_0172_),
    .A(_0164_),
    .B(_0171_));
 sg13g2_nor2_1 _1205_ (.A(_0153_),
    .B(_0172_),
    .Y(_0173_));
 sg13g2_inv_1 _1206_ (.Y(_0174_),
    .A(_0173_));
 sg13g2_nor2_1 _1207_ (.A(_0862_),
    .B(_0146_),
    .Y(_0175_));
 sg13g2_nor2_1 _1208_ (.A(_0510_),
    .B(_0175_),
    .Y(_0176_));
 sg13g2_o21ai_1 _1209_ (.B1(_0176_),
    .Y(_0177_),
    .A1(net100),
    .A2(_0147_));
 sg13g2_nand2b_1 _1210_ (.Y(_0178_),
    .B(_0576_),
    .A_N(_0171_));
 sg13g2_nor2_1 _1211_ (.A(_0177_),
    .B(_0178_),
    .Y(_0179_));
 sg13g2_nand2b_1 _1212_ (.Y(_0180_),
    .B(_0168_),
    .A_N(_0164_));
 sg13g2_a21o_2 _1213_ (.A2(_0169_),
    .A1(_1082_),
    .B1(_0041_),
    .X(_0181_));
 sg13g2_nand2_2 _1214_ (.Y(_0182_),
    .A(_0030_),
    .B(_0169_));
 sg13g2_nor3_1 _1215_ (.A(_0041_),
    .B(_0156_),
    .C(_0168_),
    .Y(_0183_));
 sg13g2_a21oi_1 _1216_ (.A1(_0084_),
    .A2(_0182_),
    .Y(_0184_),
    .B1(_0183_));
 sg13g2_nor3_1 _1217_ (.A(_1071_),
    .B(_0164_),
    .C(_0169_),
    .Y(_0185_));
 sg13g2_nor2_1 _1218_ (.A(_0181_),
    .B(_0185_),
    .Y(_0186_));
 sg13g2_nor2b_1 _1219_ (.A(_0052_),
    .B_N(_0163_),
    .Y(_0187_));
 sg13g2_nor3_1 _1220_ (.A(_0181_),
    .B(_0185_),
    .C(_0187_),
    .Y(_0188_));
 sg13g2_nor4_1 _1221_ (.A(_0378_),
    .B(_1060_),
    .C(_0180_),
    .D(_0187_),
    .Y(_0189_));
 sg13g2_a21oi_1 _1222_ (.A1(_0181_),
    .A2(_0184_),
    .Y(_0190_),
    .B1(_0189_));
 sg13g2_a21o_2 _1223_ (.A2(_0184_),
    .A1(_0181_),
    .B1(_0189_),
    .X(_0191_));
 sg13g2_o21ai_1 _1224_ (.B1(_0140_),
    .Y(_0192_),
    .A1(_0884_),
    .A2(_0146_));
 sg13g2_nor2_1 _1225_ (.A(_0895_),
    .B(_0142_),
    .Y(_0193_));
 sg13g2_or2_1 _1226_ (.X(_0194_),
    .B(_0142_),
    .A(_0895_));
 sg13g2_nand3_1 _1227_ (.B(_0873_),
    .C(_0147_),
    .A(_0367_),
    .Y(_0195_));
 sg13g2_nand3_1 _1228_ (.B(_0194_),
    .C(_0195_),
    .A(_0192_),
    .Y(_0196_));
 sg13g2_o21ai_1 _1229_ (.B1(_0873_),
    .Y(_0197_),
    .A1(_0840_),
    .A2(_0146_));
 sg13g2_nand2_1 _1230_ (.Y(_0198_),
    .A(_0895_),
    .B(_0149_));
 sg13g2_nor2_1 _1231_ (.A(_0193_),
    .B(_0197_),
    .Y(_0199_));
 sg13g2_a21oi_1 _1232_ (.A1(_0146_),
    .A2(_0193_),
    .Y(_0200_),
    .B1(_0197_));
 sg13g2_and4_1 _1233_ (.A(_0192_),
    .B(_0194_),
    .C(_0195_),
    .D(_0197_),
    .X(_0201_));
 sg13g2_inv_1 _1234_ (.Y(_0202_),
    .A(_0201_));
 sg13g2_nand2_1 _1235_ (.Y(_0203_),
    .A(_0191_),
    .B(_0201_));
 sg13g2_a21oi_1 _1236_ (.A1(_0030_),
    .A2(_0169_),
    .Y(_0204_),
    .B1(_0156_));
 sg13g2_nor3_1 _1237_ (.A(net11),
    .B(_0041_),
    .C(_0168_),
    .Y(_0205_));
 sg13g2_nor3_1 _1238_ (.A(_0187_),
    .B(_0204_),
    .C(_0205_),
    .Y(_0206_));
 sg13g2_nand2b_2 _1239_ (.Y(_0207_),
    .B(_0206_),
    .A_N(_0186_));
 sg13g2_and3_1 _1240_ (.X(_0208_),
    .A(_0873_),
    .B(_0140_),
    .C(_0147_));
 sg13g2_a21oi_1 _1241_ (.A1(_0928_),
    .A2(_0150_),
    .Y(_0209_),
    .B1(_0208_));
 sg13g2_a221oi_1 _1242_ (.B2(_0149_),
    .C1(_0208_),
    .B1(_0151_),
    .A1(_0928_),
    .Y(_0210_),
    .A2(_0150_));
 sg13g2_and3_1 _1243_ (.X(_0211_),
    .A(net3),
    .B(_0149_),
    .C(_0150_));
 sg13g2_nor2_1 _1244_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_nor2_2 _1245_ (.A(_0198_),
    .B(_0212_),
    .Y(_0213_));
 sg13g2_o21ai_1 _1246_ (.B1(_0197_),
    .Y(_0214_),
    .A1(_0210_),
    .A2(_0211_));
 sg13g2_or2_1 _1247_ (.X(_0215_),
    .B(_0207_),
    .A(_0202_));
 sg13g2_nand2_2 _1248_ (.Y(_0216_),
    .A(_0191_),
    .B(_0213_));
 sg13g2_xor2_1 _1249_ (.B(_0216_),
    .A(_0215_),
    .X(_0217_));
 sg13g2_nor3_1 _1250_ (.A(_0367_),
    .B(_0149_),
    .C(_0193_),
    .Y(_0218_));
 sg13g2_a21o_2 _1251_ (.A2(_0209_),
    .A1(_0197_),
    .B1(_0218_),
    .X(_0219_));
 sg13g2_nand3_1 _1252_ (.B(_0164_),
    .C(_0169_),
    .A(_0030_),
    .Y(_0220_));
 sg13g2_nand2_1 _1253_ (.Y(_0221_),
    .A(_0180_),
    .B(_0220_));
 sg13g2_a221oi_1 _1254_ (.B2(_0180_),
    .C1(_0183_),
    .B1(_0220_),
    .A1(_0084_),
    .Y(_0222_),
    .A2(_0182_));
 sg13g2_and3_1 _1255_ (.X(_0223_),
    .A(net11),
    .B(_0164_),
    .C(_0182_));
 sg13g2_nor2_1 _1256_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sg13g2_nor2b_2 _1257_ (.A(_0224_),
    .B_N(_0181_),
    .Y(_0225_));
 sg13g2_and2_1 _1258_ (.A(_0219_),
    .B(_0225_),
    .X(_0226_));
 sg13g2_nand2_1 _1259_ (.Y(_0227_),
    .A(_0217_),
    .B(_0226_));
 sg13g2_o21ai_1 _1260_ (.B1(_0198_),
    .Y(_0228_),
    .A1(_0152_),
    .A2(_0196_));
 sg13g2_mux2_1 _1261_ (.A0(_0928_),
    .A1(_0818_),
    .S(_0150_),
    .X(_0229_));
 sg13g2_nand2b_2 _1262_ (.Y(_0230_),
    .B(_0229_),
    .A_N(_0200_));
 sg13g2_and2_1 _1263_ (.A(_0228_),
    .B(_0230_),
    .X(_0231_));
 sg13g2_nand2_1 _1264_ (.Y(_0232_),
    .A(_0228_),
    .B(_0230_));
 sg13g2_a21oi_1 _1265_ (.A1(_0206_),
    .A2(_0221_),
    .Y(_0233_),
    .B1(_0181_));
 sg13g2_mux2_1 _1266_ (.A0(_0074_),
    .A1(_1027_),
    .S(_0182_),
    .X(_0234_));
 sg13g2_nor2_1 _1267_ (.A(_0186_),
    .B(_0234_),
    .Y(_0235_));
 sg13g2_nor2_2 _1268_ (.A(_0233_),
    .B(_0235_),
    .Y(_0236_));
 sg13g2_nand2_2 _1269_ (.Y(_0237_),
    .A(_0231_),
    .B(_0236_));
 sg13g2_nand2_2 _1270_ (.Y(_0238_),
    .A(_0213_),
    .B(_0225_));
 sg13g2_nand2_1 _1271_ (.Y(_0239_),
    .A(_0213_),
    .B(_0236_));
 sg13g2_nand2_1 _1272_ (.Y(_0240_),
    .A(_0225_),
    .B(_0231_));
 sg13g2_or2_1 _1273_ (.X(_0241_),
    .B(_0238_),
    .A(_0237_));
 sg13g2_nand2_2 _1274_ (.Y(_0242_),
    .A(_0191_),
    .B(_0219_));
 sg13g2_nand2b_1 _1275_ (.Y(_0243_),
    .B(_0219_),
    .A_N(_0207_));
 sg13g2_or2_1 _1276_ (.X(_0244_),
    .B(_0242_),
    .A(_0215_));
 sg13g2_xnor2_1 _1277_ (.Y(_0245_),
    .A(_0203_),
    .B(_0243_));
 sg13g2_nor3_1 _1278_ (.A(_0215_),
    .B(_0216_),
    .C(_0245_),
    .Y(_0246_));
 sg13g2_xor2_1 _1279_ (.B(_0240_),
    .A(_0239_),
    .X(_0247_));
 sg13g2_o21ai_1 _1280_ (.B1(_0245_),
    .Y(_0248_),
    .A1(_0215_),
    .A2(_0216_));
 sg13g2_nand2b_1 _1281_ (.Y(_0249_),
    .B(_0248_),
    .A_N(_0246_));
 sg13g2_a21o_1 _1282_ (.A2(_0248_),
    .A1(_0247_),
    .B1(_0246_),
    .X(_0250_));
 sg13g2_o21ai_1 _1283_ (.B1(_0199_),
    .Y(_0251_),
    .A1(_0210_),
    .A2(_0211_));
 sg13g2_nand2_1 _1284_ (.Y(_0252_),
    .A(_0774_),
    .B(_0150_));
 sg13g2_nand3_1 _1285_ (.B(_0873_),
    .C(_0147_),
    .A(_0818_),
    .Y(_0253_));
 sg13g2_nand3_1 _1286_ (.B(_0252_),
    .C(_0253_),
    .A(_0197_),
    .Y(_0254_));
 sg13g2_nand2_2 _1287_ (.Y(_0255_),
    .A(_0251_),
    .B(_0254_));
 sg13g2_nand2_1 _1288_ (.Y(_0256_),
    .A(_0225_),
    .B(_0255_));
 sg13g2_o21ai_1 _1289_ (.B1(_0188_),
    .Y(_0257_),
    .A1(_0222_),
    .A2(_0223_));
 sg13g2_o21ai_1 _1290_ (.B1(_0181_),
    .Y(_0258_),
    .A1(_1027_),
    .A2(_0182_));
 sg13g2_a21o_2 _1291_ (.A2(_0182_),
    .A1(_0972_),
    .B1(_0258_),
    .X(_0259_));
 sg13g2_nand2_2 _1292_ (.Y(_0260_),
    .A(_0257_),
    .B(_0259_));
 sg13g2_a21oi_1 _1293_ (.A1(_0257_),
    .A2(_0259_),
    .Y(_0261_),
    .B1(_0202_));
 sg13g2_nor3_1 _1294_ (.A(_0202_),
    .B(_0233_),
    .C(_0235_),
    .Y(_0262_));
 sg13g2_a21oi_1 _1295_ (.A1(_0257_),
    .A2(_0259_),
    .Y(_0263_),
    .B1(_0214_));
 sg13g2_nand2_1 _1296_ (.Y(_0264_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_xnor2_1 _1297_ (.Y(_0265_),
    .A(_0262_),
    .B(_0263_));
 sg13g2_xnor2_1 _1298_ (.Y(_0266_),
    .A(_0256_),
    .B(_0265_));
 sg13g2_nand3_1 _1299_ (.B(_0228_),
    .C(_0230_),
    .A(_0191_),
    .Y(_0267_));
 sg13g2_nor2_1 _1300_ (.A(_0207_),
    .B(_0232_),
    .Y(_0268_));
 sg13g2_nand3b_1 _1301_ (.B(_0228_),
    .C(_0230_),
    .Y(_0269_),
    .A_N(_0207_));
 sg13g2_or2_1 _1302_ (.X(_0270_),
    .B(_0269_),
    .A(_0242_));
 sg13g2_xor2_1 _1303_ (.B(_0269_),
    .A(_0242_),
    .X(_0271_));
 sg13g2_nor2b_1 _1304_ (.A(_0244_),
    .B_N(_0271_),
    .Y(_0272_));
 sg13g2_xnor2_1 _1305_ (.Y(_0273_),
    .A(_0244_),
    .B(_0271_));
 sg13g2_nor2b_1 _1306_ (.A(_0266_),
    .B_N(_0273_),
    .Y(_0274_));
 sg13g2_xnor2_1 _1307_ (.Y(_0275_),
    .A(_0266_),
    .B(_0273_));
 sg13g2_nand2_1 _1308_ (.Y(_0276_),
    .A(_0250_),
    .B(_0275_));
 sg13g2_xnor2_1 _1309_ (.Y(_0277_),
    .A(_0250_),
    .B(_0275_));
 sg13g2_xor2_1 _1310_ (.B(_0277_),
    .A(_0241_),
    .X(_0278_));
 sg13g2_xnor2_1 _1311_ (.Y(_0279_),
    .A(_0247_),
    .B(_0249_));
 sg13g2_nand2_1 _1312_ (.Y(_0280_),
    .A(_0278_),
    .B(_0279_));
 sg13g2_o21ai_1 _1313_ (.B1(_0276_),
    .Y(_0281_),
    .A1(_0241_),
    .A2(_0277_));
 sg13g2_o21ai_1 _1314_ (.B1(_0264_),
    .Y(_0282_),
    .A1(_0256_),
    .A2(_0265_));
 sg13g2_nor2_1 _1315_ (.A(_0272_),
    .B(_0274_),
    .Y(_0283_));
 sg13g2_nor2_1 _1316_ (.A(_0565_),
    .B(_0214_),
    .Y(_0284_));
 sg13g2_a21oi_1 _1317_ (.A1(_0251_),
    .A2(_0254_),
    .Y(_0285_),
    .B1(_0190_));
 sg13g2_a21oi_1 _1318_ (.A1(_0251_),
    .A2(_0254_),
    .Y(_0286_),
    .B1(_0207_));
 sg13g2_xnor2_1 _1319_ (.Y(_0287_),
    .A(_0267_),
    .B(_0286_));
 sg13g2_xnor2_1 _1320_ (.Y(_0288_),
    .A(_0284_),
    .B(_0287_));
 sg13g2_nor2_1 _1321_ (.A(_0270_),
    .B(_0288_),
    .Y(_0289_));
 sg13g2_xor2_1 _1322_ (.B(_0288_),
    .A(_0270_),
    .X(_0290_));
 sg13g2_nand2_1 _1323_ (.Y(_0291_),
    .A(_0521_),
    .B(_0225_));
 sg13g2_nand2_1 _1324_ (.Y(_0292_),
    .A(_0219_),
    .B(_0260_));
 sg13g2_and2_1 _1325_ (.A(_0219_),
    .B(_0236_),
    .X(_0293_));
 sg13g2_nand2_1 _1326_ (.Y(_0294_),
    .A(_0261_),
    .B(_0293_));
 sg13g2_xnor2_1 _1327_ (.Y(_0295_),
    .A(_0261_),
    .B(_0293_));
 sg13g2_xor2_1 _1328_ (.B(_0295_),
    .A(_0291_),
    .X(_0296_));
 sg13g2_xnor2_1 _1329_ (.Y(_0297_),
    .A(_0290_),
    .B(_0296_));
 sg13g2_nor2_1 _1330_ (.A(_0283_),
    .B(_0297_),
    .Y(_0298_));
 sg13g2_xor2_1 _1331_ (.B(_0297_),
    .A(_0283_),
    .X(_0299_));
 sg13g2_xnor2_1 _1332_ (.Y(_0300_),
    .A(_0282_),
    .B(_0299_));
 sg13g2_nor2b_2 _1333_ (.A(_0300_),
    .B_N(_0281_),
    .Y(_0301_));
 sg13g2_xor2_1 _1334_ (.B(_0300_),
    .A(_0281_),
    .X(_0302_));
 sg13g2_nor3_1 _1335_ (.A(_0227_),
    .B(_0280_),
    .C(_0302_),
    .Y(_0303_));
 sg13g2_o21ai_1 _1336_ (.B1(_0302_),
    .Y(_0304_),
    .A1(_0227_),
    .A2(_0280_));
 sg13g2_nand2b_1 _1337_ (.Y(_0305_),
    .B(_0304_),
    .A_N(_0303_));
 sg13g2_xnor2_1 _1338_ (.Y(_0306_),
    .A(_0217_),
    .B(_0226_));
 sg13g2_inv_1 _1339_ (.Y(_0307_),
    .A(_0306_));
 sg13g2_nand2_1 _1340_ (.Y(_0308_),
    .A(_0201_),
    .B(_0225_));
 sg13g2_nor2_1 _1341_ (.A(_0215_),
    .B(_0238_),
    .Y(_0309_));
 sg13g2_nand2_1 _1342_ (.Y(_0310_),
    .A(_0307_),
    .B(_0309_));
 sg13g2_and4_1 _1343_ (.A(_0278_),
    .B(_0279_),
    .C(_0307_),
    .D(_0309_),
    .X(_0311_));
 sg13g2_a21oi_2 _1344_ (.B1(_0303_),
    .Y(_0312_),
    .A2(_0311_),
    .A1(_0304_));
 sg13g2_a21oi_2 _1345_ (.B1(_0298_),
    .Y(_0313_),
    .A2(_0299_),
    .A1(_0282_));
 sg13g2_o21ai_1 _1346_ (.B1(_0294_),
    .Y(_0314_),
    .A1(_0291_),
    .A2(_0295_));
 sg13g2_a21oi_1 _1347_ (.A1(_0290_),
    .A2(_0296_),
    .Y(_0315_),
    .B1(_0289_));
 sg13g2_nand2_1 _1348_ (.Y(_0316_),
    .A(_0231_),
    .B(_0260_));
 sg13g2_or2_1 _1349_ (.X(_0317_),
    .B(_0292_),
    .A(_0237_));
 sg13g2_xnor2_1 _1350_ (.Y(_0318_),
    .A(_0237_),
    .B(_0292_));
 sg13g2_a22oi_1 _1351_ (.Y(_0319_),
    .B1(_0287_),
    .B2(_0284_),
    .A2(_0285_),
    .A1(_0268_));
 sg13g2_nand2_1 _1352_ (.Y(_0320_),
    .A(_0576_),
    .B(_0201_));
 sg13g2_nor2_1 _1353_ (.A(_0510_),
    .B(_0207_),
    .Y(_0321_));
 sg13g2_nand2_1 _1354_ (.Y(_0322_),
    .A(_0285_),
    .B(_0321_));
 sg13g2_xnor2_1 _1355_ (.Y(_0323_),
    .A(_0285_),
    .B(_0321_));
 sg13g2_xnor2_1 _1356_ (.Y(_0324_),
    .A(_0320_),
    .B(_0323_));
 sg13g2_or2_1 _1357_ (.X(_0325_),
    .B(_0324_),
    .A(_0319_));
 sg13g2_and2_1 _1358_ (.A(_0319_),
    .B(_0324_),
    .X(_0326_));
 sg13g2_xor2_1 _1359_ (.B(_0324_),
    .A(_0319_),
    .X(_0327_));
 sg13g2_xnor2_1 _1360_ (.Y(_0328_),
    .A(_0318_),
    .B(_0327_));
 sg13g2_nor2b_1 _1361_ (.A(_0315_),
    .B_N(_0328_),
    .Y(_0329_));
 sg13g2_xnor2_1 _1362_ (.Y(_0330_),
    .A(_0315_),
    .B(_0328_));
 sg13g2_xnor2_1 _1363_ (.Y(_0331_),
    .A(_0314_),
    .B(_0330_));
 sg13g2_nor2_1 _1364_ (.A(_0313_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_or2_1 _1365_ (.X(_0333_),
    .B(_0331_),
    .A(_0313_));
 sg13g2_a21oi_1 _1366_ (.A1(_0314_),
    .A2(_0330_),
    .Y(_0334_),
    .B1(_0329_));
 sg13g2_o21ai_1 _1367_ (.B1(_0325_),
    .Y(_0335_),
    .A1(_0318_),
    .A2(_0326_));
 sg13g2_nand2_2 _1368_ (.Y(_0336_),
    .A(_0255_),
    .B(_0260_));
 sg13g2_nand2_1 _1369_ (.Y(_0337_),
    .A(_0236_),
    .B(_0255_));
 sg13g2_or2_1 _1370_ (.X(_0338_),
    .B(_0336_),
    .A(_0237_));
 sg13g2_inv_1 _1371_ (.Y(_0339_),
    .A(_0338_));
 sg13g2_xnor2_1 _1372_ (.Y(_0340_),
    .A(_0316_),
    .B(_0337_));
 sg13g2_o21ai_1 _1373_ (.B1(_0322_),
    .Y(_0341_),
    .A1(_0320_),
    .A2(_0323_));
 sg13g2_a22oi_1 _1374_ (.Y(_0342_),
    .B1(_0219_),
    .B2(_0576_),
    .A2(_0191_),
    .A1(_0521_));
 sg13g2_a21oi_1 _1375_ (.A1(_0191_),
    .A2(_0219_),
    .Y(_0343_),
    .B1(_0342_));
 sg13g2_nand2_1 _1376_ (.Y(_0344_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_xnor2_1 _1377_ (.Y(_0345_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_xor2_1 _1378_ (.B(_0345_),
    .A(_0340_),
    .X(_0346_));
 sg13g2_and2_1 _1379_ (.A(_0335_),
    .B(_0346_),
    .X(_0347_));
 sg13g2_nand2_1 _1380_ (.Y(_0348_),
    .A(_0335_),
    .B(_0346_));
 sg13g2_xnor2_1 _1381_ (.Y(_0349_),
    .A(_0335_),
    .B(_0346_));
 sg13g2_nor2_1 _1382_ (.A(_0317_),
    .B(_0349_),
    .Y(_0350_));
 sg13g2_xnor2_1 _1383_ (.Y(_0351_),
    .A(_0317_),
    .B(_0349_));
 sg13g2_or2_1 _1384_ (.X(_0352_),
    .B(_0351_),
    .A(_0334_));
 sg13g2_xor2_1 _1385_ (.B(_0351_),
    .A(_0334_),
    .X(_0353_));
 sg13g2_and2_1 _1386_ (.A(_0332_),
    .B(_0353_),
    .X(_0354_));
 sg13g2_xnor2_1 _1387_ (.Y(_0355_),
    .A(_0332_),
    .B(_0353_));
 sg13g2_nand2_1 _1388_ (.Y(_0356_),
    .A(_0313_),
    .B(_0331_));
 sg13g2_xor2_1 _1389_ (.B(_0331_),
    .A(_0313_),
    .X(_0357_));
 sg13g2_nand2_1 _1390_ (.Y(_0358_),
    .A(_0301_),
    .B(_0357_));
 sg13g2_xnor2_1 _1391_ (.Y(_0359_),
    .A(_0301_),
    .B(_0357_));
 sg13g2_or2_1 _1392_ (.X(_0360_),
    .B(_0359_),
    .A(_0355_));
 sg13g2_nor2_1 _1393_ (.A(_0312_),
    .B(_0360_),
    .Y(_0361_));
 sg13g2_and4_1 _1394_ (.A(_0301_),
    .B(_0333_),
    .C(_0353_),
    .D(_0356_),
    .X(_0362_));
 sg13g2_o21ai_1 _1395_ (.B1(_0348_),
    .Y(_0363_),
    .A1(_0317_),
    .A2(_0349_));
 sg13g2_o21ai_1 _1396_ (.B1(_0344_),
    .Y(_0364_),
    .A1(_0340_),
    .A2(_0345_));
 sg13g2_nor2_1 _1397_ (.A(_0232_),
    .B(_0242_),
    .Y(_0365_));
 sg13g2_o21ai_1 _1398_ (.B1(_0242_),
    .Y(_0366_),
    .A1(_0565_),
    .A2(_0232_));
 sg13g2_nand2b_1 _1399_ (.Y(_0368_),
    .B(_0366_),
    .A_N(_0365_));
 sg13g2_nand2_1 _1400_ (.Y(_0369_),
    .A(_0521_),
    .B(_0236_));
 sg13g2_or2_1 _1401_ (.X(_0370_),
    .B(_0369_),
    .A(_0336_));
 sg13g2_xnor2_1 _1402_ (.Y(_0371_),
    .A(_0336_),
    .B(_0369_));
 sg13g2_nor2_1 _1403_ (.A(_0368_),
    .B(_0371_),
    .Y(_0372_));
 sg13g2_xor2_1 _1404_ (.B(_0371_),
    .A(_0368_),
    .X(_0373_));
 sg13g2_and2_1 _1405_ (.A(_0364_),
    .B(_0373_),
    .X(_0374_));
 sg13g2_or2_1 _1406_ (.X(_0375_),
    .B(_0373_),
    .A(_0364_));
 sg13g2_xor2_1 _1407_ (.B(_0373_),
    .A(_0364_),
    .X(_0376_));
 sg13g2_xnor2_1 _1408_ (.Y(_0377_),
    .A(_0338_),
    .B(_0376_));
 sg13g2_and2_1 _1409_ (.A(_0363_),
    .B(_0377_),
    .X(_0379_));
 sg13g2_nand2_1 _1410_ (.Y(_0380_),
    .A(_0363_),
    .B(_0377_));
 sg13g2_a22oi_1 _1411_ (.Y(_0381_),
    .B1(_0260_),
    .B2(_0521_),
    .A2(_0255_),
    .A1(_0576_));
 sg13g2_a21oi_1 _1412_ (.A1(_0255_),
    .A2(_0260_),
    .Y(_0382_),
    .B1(_0381_));
 sg13g2_nor2_1 _1413_ (.A(_0365_),
    .B(_0372_),
    .Y(_0383_));
 sg13g2_xnor2_1 _1414_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_nor3_1 _1415_ (.A(_0336_),
    .B(_0369_),
    .C(_0383_),
    .Y(_0385_));
 sg13g2_xnor2_1 _1416_ (.Y(_0386_),
    .A(_0370_),
    .B(_0384_));
 sg13g2_a21oi_1 _1417_ (.A1(_0339_),
    .A2(_0375_),
    .Y(_0387_),
    .B1(_0374_));
 sg13g2_nor2b_1 _1418_ (.A(_0387_),
    .B_N(_0386_),
    .Y(_0388_));
 sg13g2_xor2_1 _1419_ (.B(_0387_),
    .A(_0386_),
    .X(_0390_));
 sg13g2_nor2_1 _1420_ (.A(_0380_),
    .B(_0390_),
    .Y(_0391_));
 sg13g2_nand2_1 _1421_ (.Y(_0392_),
    .A(_0380_),
    .B(_0390_));
 sg13g2_nor3_1 _1422_ (.A(_0347_),
    .B(_0350_),
    .C(_0377_),
    .Y(_0393_));
 sg13g2_or2_1 _1423_ (.X(_0394_),
    .B(_0393_),
    .A(_0379_));
 sg13g2_nor2_1 _1424_ (.A(_0352_),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_nor4_1 _1425_ (.A(_0352_),
    .B(_0379_),
    .C(_0390_),
    .D(_0393_),
    .Y(_0396_));
 sg13g2_nor4_1 _1426_ (.A(_0354_),
    .B(_0362_),
    .C(_0391_),
    .D(_0396_),
    .Y(_0397_));
 sg13g2_o21ai_1 _1427_ (.B1(_0397_),
    .Y(_0398_),
    .A1(_0312_),
    .A2(_0360_));
 sg13g2_nand2_1 _1428_ (.Y(_0399_),
    .A(_0352_),
    .B(_0394_));
 sg13g2_or2_1 _1429_ (.X(_0401_),
    .B(_0399_),
    .A(_0391_));
 sg13g2_and3_1 _1430_ (.X(_0402_),
    .A(_0392_),
    .B(_0398_),
    .C(_0401_));
 sg13g2_o21ai_1 _1431_ (.B1(_0336_),
    .Y(_0403_),
    .A1(_0381_),
    .A2(_0383_));
 sg13g2_nor2_1 _1432_ (.A(net98),
    .B(_0403_),
    .Y(_0404_));
 sg13g2_nor2_1 _1433_ (.A(_0385_),
    .B(_0404_),
    .Y(_0405_));
 sg13g2_nor2b_1 _1434_ (.A(_0405_),
    .B_N(_0388_),
    .Y(_0406_));
 sg13g2_xnor2_1 _1435_ (.Y(_0407_),
    .A(_0388_),
    .B(_0405_));
 sg13g2_nand4_1 _1436_ (.B(_0398_),
    .C(_0401_),
    .A(_0392_),
    .Y(_0408_),
    .D(_0407_));
 sg13g2_nor2_1 _1437_ (.A(_0403_),
    .B(_0406_),
    .Y(_0409_));
 sg13g2_nand2_1 _1438_ (.Y(_0410_),
    .A(_0408_),
    .B(_0409_));
 sg13g2_xor2_1 _1439_ (.B(_0178_),
    .A(_0177_),
    .X(_0412_));
 sg13g2_inv_1 _1440_ (.Y(_0413_),
    .A(_0412_));
 sg13g2_a21oi_1 _1441_ (.A1(_0408_),
    .A2(_0409_),
    .Y(_0414_),
    .B1(_0413_));
 sg13g2_xor2_1 _1442_ (.B(_0172_),
    .A(_0153_),
    .X(_0415_));
 sg13g2_o21ai_1 _1443_ (.B1(_0415_),
    .Y(_0416_),
    .A1(_0179_),
    .A2(_0414_));
 sg13g2_xor2_1 _1444_ (.B(_0104_),
    .A(_0950_),
    .X(_0417_));
 sg13g2_xnor2_1 _1445_ (.Y(_0418_),
    .A(_0950_),
    .B(_0104_));
 sg13g2_a21oi_1 _1446_ (.A1(_0174_),
    .A2(_0416_),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_nor2_1 _1447_ (.A(_0114_),
    .B(_0419_),
    .Y(_0420_));
 sg13g2_a22oi_1 _1448_ (.Y(_0421_),
    .B1(_0730_),
    .B2(_0576_),
    .A2(net101),
    .A1(_0521_));
 sg13g2_nor2_1 _1449_ (.A(_0741_),
    .B(_0421_),
    .Y(_0423_));
 sg13g2_nor4_1 _1450_ (.A(_0741_),
    .B(_0114_),
    .C(_0419_),
    .D(_0421_),
    .Y(_0424_));
 sg13g2_or4_1 _1451_ (.A(_0741_),
    .B(_0114_),
    .C(_0419_),
    .D(_0421_),
    .X(_0425_));
 sg13g2_nand2_2 _1452_ (.Y(_0426_),
    .A(_0752_),
    .B(_0425_));
 sg13g2_inv_2 _1453_ (.Y(_0427_),
    .A(_0426_));
 sg13g2_nor3_1 _1454_ (.A(_0752_),
    .B(_0114_),
    .C(_0419_),
    .Y(_0428_));
 sg13g2_xnor2_1 _1455_ (.Y(_0429_),
    .A(_0420_),
    .B(_0423_));
 sg13g2_xnor2_1 _1456_ (.Y(_0430_),
    .A(net92),
    .B(_0413_));
 sg13g2_inv_1 _1457_ (.Y(_0431_),
    .A(_0430_));
 sg13g2_or3_1 _1458_ (.A(_0179_),
    .B(_0414_),
    .C(_0415_),
    .X(_0432_));
 sg13g2_and2_1 _1459_ (.A(_0416_),
    .B(_0432_),
    .X(_0434_));
 sg13g2_or2_1 _1460_ (.X(_0435_),
    .B(_0434_),
    .A(_0430_));
 sg13g2_and3_1 _1461_ (.X(_0436_),
    .A(_0174_),
    .B(_0416_),
    .C(_0417_));
 sg13g2_a21oi_1 _1462_ (.A1(_0174_),
    .A2(_0416_),
    .Y(_0437_),
    .B1(_0417_));
 sg13g2_nor2_1 _1463_ (.A(_0436_),
    .B(_0437_),
    .Y(_0438_));
 sg13g2_nor4_1 _1464_ (.A(_0430_),
    .B(_0434_),
    .C(_0436_),
    .D(_0437_),
    .Y(_0439_));
 sg13g2_o21ai_1 _1465_ (.B1(_0435_),
    .Y(_0440_),
    .A1(_0741_),
    .A2(_0424_));
 sg13g2_a21o_1 _1466_ (.A2(_0425_),
    .A1(_0752_),
    .B1(_0439_),
    .X(_0441_));
 sg13g2_a21o_2 _1467_ (.A2(_0441_),
    .A1(_0429_),
    .B1(_0428_),
    .X(_0442_));
 sg13g2_o21ai_1 _1468_ (.B1(_0430_),
    .Y(_0443_),
    .A1(_0741_),
    .A2(_0424_));
 sg13g2_xnor2_1 _1469_ (.Y(_0445_),
    .A(_0434_),
    .B(_0443_));
 sg13g2_xor2_1 _1470_ (.B(_0443_),
    .A(_0434_),
    .X(_0446_));
 sg13g2_nor2_1 _1471_ (.A(_0442_),
    .B(_0445_),
    .Y(_0447_));
 sg13g2_nand2b_2 _1472_ (.Y(_0448_),
    .B(_0446_),
    .A_N(_0442_));
 sg13g2_xnor2_1 _1473_ (.Y(_0449_),
    .A(_0438_),
    .B(_0440_));
 sg13g2_nor2_1 _1474_ (.A(_0446_),
    .B(_0449_),
    .Y(_0450_));
 sg13g2_a221oi_1 _1475_ (.B2(_0441_),
    .C1(_0431_),
    .B1(_0429_),
    .A1(_0741_),
    .Y(_0451_),
    .A2(_0420_));
 sg13g2_nor2b_1 _1476_ (.A(_0450_),
    .B_N(_0451_),
    .Y(_0452_));
 sg13g2_o21ai_1 _1477_ (.B1(_0451_),
    .Y(_0453_),
    .A1(_0446_),
    .A2(_0449_));
 sg13g2_nand2_1 _1478_ (.Y(_0454_),
    .A(_0426_),
    .B(_0453_));
 sg13g2_nor4_2 _1479_ (.A(_0427_),
    .B(_0430_),
    .C(_0442_),
    .Y(_0456_),
    .D(_0445_));
 sg13g2_nor2b_2 _1480_ (.A(_0442_),
    .B_N(_0449_),
    .Y(_0457_));
 sg13g2_nor2_2 _1481_ (.A(_0456_),
    .B(_0457_),
    .Y(_0458_));
 sg13g2_or2_1 _1482_ (.X(_0459_),
    .B(_0457_),
    .A(_0456_));
 sg13g2_a21oi_2 _1483_ (.B1(_0447_),
    .Y(_0460_),
    .A2(_0453_),
    .A1(_0426_));
 sg13g2_nor2_2 _1484_ (.A(_0456_),
    .B(_0460_),
    .Y(_0461_));
 sg13g2_or2_1 _1485_ (.X(_0462_),
    .B(_0460_),
    .A(_0456_));
 sg13g2_o21ai_1 _1486_ (.B1(_0426_),
    .Y(_0463_),
    .A1(_0456_),
    .A2(_0460_));
 sg13g2_nand2_1 _1487_ (.Y(_0464_),
    .A(_0453_),
    .B(_0461_));
 sg13g2_a21o_1 _1488_ (.A2(_0464_),
    .A1(_0463_),
    .B1(_0458_),
    .X(_0465_));
 sg13g2_inv_1 _1489_ (.Y(_0467_),
    .A(_0465_));
 sg13g2_xnor2_1 _1490_ (.Y(_0468_),
    .A(_0426_),
    .B(_0453_));
 sg13g2_inv_1 _1491_ (.Y(_0469_),
    .A(net89));
 sg13g2_o21ai_1 _1492_ (.B1(_0358_),
    .Y(_0470_),
    .A1(_0312_),
    .A2(_0359_));
 sg13g2_xor2_1 _1493_ (.B(_0470_),
    .A(_0355_),
    .X(_0471_));
 sg13g2_a21oi_1 _1494_ (.A1(_0408_),
    .A2(_0409_),
    .Y(_0472_),
    .B1(_0471_));
 sg13g2_xnor2_1 _1495_ (.Y(_0473_),
    .A(_0312_),
    .B(_0359_));
 sg13g2_or2_1 _1496_ (.X(_0474_),
    .B(_0473_),
    .A(net90));
 sg13g2_nor2b_1 _1497_ (.A(_0472_),
    .B_N(_0474_),
    .Y(_0475_));
 sg13g2_nand2b_1 _1498_ (.Y(_0476_),
    .B(_0474_),
    .A_N(_0472_));
 sg13g2_nand2_1 _1499_ (.Y(_0478_),
    .A(_0468_),
    .B(_0475_));
 sg13g2_xor2_1 _1500_ (.B(_0311_),
    .A(_0305_),
    .X(_0479_));
 sg13g2_mux2_1 _1501_ (.A0(_0479_),
    .A1(_0473_),
    .S(net90),
    .X(_0480_));
 sg13g2_inv_1 _1502_ (.Y(_0481_),
    .A(_0480_));
 sg13g2_mux2_1 _1503_ (.A0(_0481_),
    .A1(_0476_),
    .S(net89),
    .X(_0482_));
 sg13g2_o21ai_1 _1504_ (.B1(_0478_),
    .Y(_0483_),
    .A1(_0468_),
    .A2(_0481_));
 sg13g2_nand2b_1 _1505_ (.Y(_0484_),
    .B(_0399_),
    .A_N(_0395_));
 sg13g2_nor3_1 _1506_ (.A(_0354_),
    .B(_0361_),
    .C(_0362_),
    .Y(_0485_));
 sg13g2_nor2_1 _1507_ (.A(_0484_),
    .B(_0485_),
    .Y(_0486_));
 sg13g2_xor2_1 _1508_ (.B(_0485_),
    .A(_0484_),
    .X(_0487_));
 sg13g2_nand2_1 _1509_ (.Y(_0489_),
    .A(net91),
    .B(_0487_));
 sg13g2_o21ai_1 _1510_ (.B1(_0489_),
    .Y(_0490_),
    .A1(net91),
    .A2(_0471_));
 sg13g2_inv_1 _1511_ (.Y(_0491_),
    .A(_0490_));
 sg13g2_nor2b_1 _1512_ (.A(_0391_),
    .B_N(_0392_),
    .Y(_0492_));
 sg13g2_nor2_1 _1513_ (.A(_0395_),
    .B(_0486_),
    .Y(_0493_));
 sg13g2_xnor2_1 _1514_ (.Y(_0494_),
    .A(_0492_),
    .B(_0493_));
 sg13g2_mux2_1 _1515_ (.A0(_0487_),
    .A1(_0494_),
    .S(net91),
    .X(_0495_));
 sg13g2_inv_1 _1516_ (.Y(_0496_),
    .A(_0495_));
 sg13g2_mux2_1 _1517_ (.A0(_0490_),
    .A1(_0495_),
    .S(net89),
    .X(_0497_));
 sg13g2_xnor2_1 _1518_ (.Y(_0498_),
    .A(_0402_),
    .B(_0407_));
 sg13g2_nand2_1 _1519_ (.Y(_0500_),
    .A(net90),
    .B(_0498_));
 sg13g2_o21ai_1 _1520_ (.B1(_0500_),
    .Y(_0501_),
    .A1(net91),
    .A2(_0494_));
 sg13g2_inv_1 _1521_ (.Y(_0502_),
    .A(_0501_));
 sg13g2_o21ai_1 _1522_ (.B1(_0502_),
    .Y(_0503_),
    .A1(_0426_),
    .A2(_0453_));
 sg13g2_nand2_1 _1523_ (.Y(_0504_),
    .A(_0454_),
    .B(_0503_));
 sg13g2_o21ai_1 _1524_ (.B1(_0463_),
    .Y(_0505_),
    .A1(_0448_),
    .A2(_0504_));
 sg13g2_nand2_1 _1525_ (.Y(_0506_),
    .A(_0462_),
    .B(_0497_));
 sg13g2_a21oi_1 _1526_ (.A1(_0461_),
    .A2(_0482_),
    .Y(_0507_),
    .B1(_0458_));
 sg13g2_a22oi_1 _1527_ (.Y(_0508_),
    .B1(_0506_),
    .B2(_0507_),
    .A2(_0505_),
    .A1(_0458_));
 sg13g2_nand2_1 _1528_ (.Y(_0509_),
    .A(_0227_),
    .B(_0310_));
 sg13g2_nand2_1 _1529_ (.Y(_0511_),
    .A(_0279_),
    .B(_0509_));
 sg13g2_xor2_1 _1530_ (.B(_0511_),
    .A(_0278_),
    .X(_0512_));
 sg13g2_mux2_1 _1531_ (.A0(_0512_),
    .A1(_0479_),
    .S(net90),
    .X(_0513_));
 sg13g2_inv_1 _1532_ (.Y(_0514_),
    .A(_0513_));
 sg13g2_mux2_1 _1533_ (.A0(_0513_),
    .A1(_0480_),
    .S(_0468_),
    .X(_0515_));
 sg13g2_mux2_1 _1534_ (.A0(_0476_),
    .A1(_0490_),
    .S(net89),
    .X(_0516_));
 sg13g2_mux2_1 _1535_ (.A0(_0475_),
    .A1(_0491_),
    .S(net89),
    .X(_0517_));
 sg13g2_mux2_1 _1536_ (.A0(_0496_),
    .A1(_0501_),
    .S(net89),
    .X(_0518_));
 sg13g2_mux2_1 _1537_ (.A0(_0495_),
    .A1(_0502_),
    .S(net89),
    .X(_0519_));
 sg13g2_nand2_1 _1538_ (.Y(_0520_),
    .A(_0461_),
    .B(_0519_));
 sg13g2_nand2_1 _1539_ (.Y(_0522_),
    .A(_0448_),
    .B(_0452_));
 sg13g2_mux4_1 _1540_ (.S0(_0459_),
    .A0(_0453_),
    .A1(_0517_),
    .A2(_0518_),
    .A3(_0515_),
    .S1(_0461_),
    .X(_0523_));
 sg13g2_a221oi_1 _1541_ (.B2(_0507_),
    .C1(_0523_),
    .B1(_0506_),
    .A1(_0458_),
    .Y(_0524_),
    .A2(_0505_));
 sg13g2_a21oi_1 _1542_ (.A1(_0462_),
    .A2(_0519_),
    .Y(_0525_),
    .B1(_0516_));
 sg13g2_mux4_1 _1543_ (.S0(_0461_),
    .A0(_0427_),
    .A1(_0452_),
    .A2(_0519_),
    .A3(_0516_),
    .S1(_0459_),
    .X(_0526_));
 sg13g2_nor2_1 _1544_ (.A(_0427_),
    .B(_0459_),
    .Y(_0527_));
 sg13g2_nand2_1 _1545_ (.Y(_0528_),
    .A(_0426_),
    .B(_0458_));
 sg13g2_nand3_1 _1546_ (.B(_0454_),
    .C(_0503_),
    .A(_0448_),
    .Y(_0529_));
 sg13g2_o21ai_1 _1547_ (.B1(_0529_),
    .Y(_0530_),
    .A1(_0462_),
    .A2(_0497_));
 sg13g2_a21oi_1 _1548_ (.A1(_0459_),
    .A2(_0530_),
    .Y(_0531_),
    .B1(_0527_));
 sg13g2_nand3_1 _1549_ (.B(_0526_),
    .C(_0531_),
    .A(_0524_),
    .Y(_0533_));
 sg13g2_nand3_1 _1550_ (.B(_0520_),
    .C(_0522_),
    .A(_0459_),
    .Y(_0534_));
 sg13g2_nand4_1 _1551_ (.B(_0526_),
    .C(_0531_),
    .A(_0524_),
    .Y(_0535_),
    .D(_0534_));
 sg13g2_a21oi_1 _1552_ (.A1(_0459_),
    .A2(_0505_),
    .Y(_0536_),
    .B1(_0527_));
 sg13g2_nand2b_1 _1553_ (.Y(_0537_),
    .B(_0536_),
    .A_N(_0535_));
 sg13g2_o21ai_1 _1554_ (.B1(_0426_),
    .Y(_0538_),
    .A1(_0467_),
    .A2(_0537_));
 sg13g2_xor2_1 _1555_ (.B(net104),
    .A(net105),
    .X(_0539_));
 sg13g2_xnor2_1 _1556_ (.Y(_0540_),
    .A(net105),
    .B(net104));
 sg13g2_nand2_1 _1557_ (.Y(_0541_),
    .A(_0465_),
    .B(_0528_));
 sg13g2_mux2_1 _1558_ (.A0(_0465_),
    .A1(_0541_),
    .S(_0537_),
    .X(_0542_));
 sg13g2_xor2_1 _1559_ (.B(_0536_),
    .A(_0535_),
    .X(_0544_));
 sg13g2_nand2_1 _1560_ (.Y(_0545_),
    .A(_0528_),
    .B(_0534_));
 sg13g2_mux2_1 _1561_ (.A0(_0534_),
    .A1(_0545_),
    .S(_0533_),
    .X(_0546_));
 sg13g2_a21o_1 _1562_ (.A2(_0526_),
    .A1(_0524_),
    .B1(_0531_),
    .X(_0547_));
 sg13g2_nand2_1 _1563_ (.Y(_0548_),
    .A(_0533_),
    .B(_0547_));
 sg13g2_xor2_1 _1564_ (.B(_0509_),
    .A(_0279_),
    .X(_0549_));
 sg13g2_nand2_1 _1565_ (.Y(_0550_),
    .A(net90),
    .B(_0549_));
 sg13g2_xor2_1 _1566_ (.B(_0309_),
    .A(_0306_),
    .X(_0551_));
 sg13g2_inv_1 _1567_ (.Y(_0552_),
    .A(_0551_));
 sg13g2_o21ai_1 _1568_ (.B1(_0550_),
    .Y(_0553_),
    .A1(net90),
    .A2(_0551_));
 sg13g2_o21ai_1 _1569_ (.B1(_0308_),
    .Y(_0555_),
    .A1(_0207_),
    .A2(_0214_));
 sg13g2_o21ai_1 _1570_ (.B1(_0555_),
    .Y(_0556_),
    .A1(_0215_),
    .A2(_0238_));
 sg13g2_nor2_1 _1571_ (.A(net92),
    .B(_0556_),
    .Y(_0557_));
 sg13g2_a21oi_1 _1572_ (.A1(net92),
    .A2(_0552_),
    .Y(_0558_),
    .B1(_0557_));
 sg13g2_nand2b_1 _1573_ (.Y(_0559_),
    .B(_0558_),
    .A_N(_0553_));
 sg13g2_mux2_1 _1574_ (.A0(_0238_),
    .A1(_0556_),
    .S(net92),
    .X(_0560_));
 sg13g2_or2_1 _1575_ (.X(_0561_),
    .B(_0549_),
    .A(net90));
 sg13g2_nand2_1 _1576_ (.Y(_0562_),
    .A(net90),
    .B(_0512_));
 sg13g2_and2_1 _1577_ (.A(net89),
    .B(_0514_),
    .X(_0563_));
 sg13g2_xor2_1 _1578_ (.B(_0460_),
    .A(_0457_),
    .X(_0564_));
 sg13g2_a21oi_1 _1579_ (.A1(_0483_),
    .A2(_0515_),
    .Y(_0566_),
    .B1(_0564_));
 sg13g2_nor3_1 _1580_ (.A(_0456_),
    .B(_0460_),
    .C(_0560_),
    .Y(_0567_));
 sg13g2_o21ai_1 _1581_ (.B1(_0469_),
    .Y(_0568_),
    .A1(_0553_),
    .A2(_0567_));
 sg13g2_a221oi_1 _1582_ (.B2(_0562_),
    .C1(_0563_),
    .B1(_0561_),
    .A1(_0461_),
    .Y(_0569_),
    .A2(_0559_));
 sg13g2_a21oi_1 _1583_ (.A1(_0568_),
    .A2(_0569_),
    .Y(_0570_),
    .B1(_0458_));
 sg13g2_a21oi_1 _1584_ (.A1(_0462_),
    .A2(_0504_),
    .Y(_0571_),
    .B1(_0497_));
 sg13g2_a21oi_1 _1585_ (.A1(_0525_),
    .A2(_0571_),
    .Y(_0572_),
    .B1(_0459_));
 sg13g2_or4_1 _1586_ (.A(_0508_),
    .B(_0566_),
    .C(_0570_),
    .D(_0572_),
    .X(_0573_));
 sg13g2_xnor2_1 _1587_ (.Y(_0574_),
    .A(_0508_),
    .B(_0523_));
 sg13g2_and2_1 _1588_ (.A(_0573_),
    .B(_0574_),
    .X(_0575_));
 sg13g2_nand2_1 _1589_ (.Y(_0577_),
    .A(_0573_),
    .B(_0574_));
 sg13g2_xor2_1 _1590_ (.B(_0526_),
    .A(_0524_),
    .X(_0578_));
 sg13g2_inv_2 _1591_ (.Y(_0579_),
    .A(_0578_));
 sg13g2_a221oi_1 _1592_ (.B2(_0574_),
    .C1(_0578_),
    .B1(_0573_),
    .A1(_0533_),
    .Y(_0580_),
    .A2(_0547_));
 sg13g2_and2_1 _1593_ (.A(_0546_),
    .B(_0580_),
    .X(_0581_));
 sg13g2_nand2_1 _1594_ (.Y(_0582_),
    .A(_0546_),
    .B(_0580_));
 sg13g2_and3_1 _1595_ (.X(_0583_),
    .A(_0544_),
    .B(_0546_),
    .C(_0580_));
 sg13g2_nor2_1 _1596_ (.A(_0540_),
    .B(_0580_),
    .Y(_0584_));
 sg13g2_nand2_1 _1597_ (.Y(_0585_),
    .A(_0539_),
    .B(_0582_));
 sg13g2_o21ai_1 _1598_ (.B1(_0542_),
    .Y(_0586_),
    .A1(_0540_),
    .A2(_0583_));
 sg13g2_a21oi_1 _1599_ (.A1(_0542_),
    .A2(_0583_),
    .Y(_0588_),
    .B1(_0540_));
 sg13g2_xnor2_1 _1600_ (.Y(_0589_),
    .A(_0538_),
    .B(_0588_));
 sg13g2_nor2_2 _1601_ (.A(net97),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_o21ai_1 _1602_ (.B1(_0609_),
    .Y(_0591_),
    .A1(net97),
    .A2(_0540_));
 sg13g2_inv_1 _1603_ (.Y(_0592_),
    .A(_0591_));
 sg13g2_or3_1 _1604_ (.A(_0540_),
    .B(_0542_),
    .C(_0583_),
    .X(_0593_));
 sg13g2_and3_2 _1605_ (.X(_0594_),
    .A(net99),
    .B(_0586_),
    .C(_0593_));
 sg13g2_o21ai_1 _1606_ (.B1(net99),
    .Y(_0595_),
    .A1(_0544_),
    .A2(_0585_));
 sg13g2_a21oi_1 _1607_ (.A1(_0544_),
    .A2(_0585_),
    .Y(_0596_),
    .B1(_0595_));
 sg13g2_xnor2_1 _1608_ (.Y(_0597_),
    .A(_0546_),
    .B(_0584_));
 sg13g2_and2_1 _1609_ (.A(net99),
    .B(_0597_),
    .X(_0599_));
 sg13g2_a21oi_1 _1610_ (.A1(_0544_),
    .A2(_0581_),
    .Y(_0600_),
    .B1(net97));
 sg13g2_nor2_1 _1611_ (.A(_0594_),
    .B(_0600_),
    .Y(_0601_));
 sg13g2_o21ai_1 _1612_ (.B1(_0591_),
    .Y(_0602_),
    .A1(_0594_),
    .A2(_0600_));
 sg13g2_xor2_1 _1613_ (.B(_0602_),
    .A(_0590_),
    .X(_0603_));
 sg13g2_nor2_2 _1614_ (.A(net97),
    .B(_0546_),
    .Y(_0604_));
 sg13g2_xor2_1 _1615_ (.B(_0604_),
    .A(net88),
    .X(_0605_));
 sg13g2_a21oi_1 _1616_ (.A1(_0577_),
    .A2(_0579_),
    .Y(_0606_),
    .B1(_0540_));
 sg13g2_xnor2_1 _1617_ (.Y(_0607_),
    .A(_0548_),
    .B(_0606_));
 sg13g2_nor2_1 _1618_ (.A(net98),
    .B(_0548_),
    .Y(_0608_));
 sg13g2_xnor2_1 _1619_ (.Y(_0610_),
    .A(net88),
    .B(_0608_));
 sg13g2_nand2_2 _1620_ (.Y(_0611_),
    .A(net99),
    .B(_0575_));
 sg13g2_o21ai_1 _1621_ (.B1(_0579_),
    .Y(_0612_),
    .A1(_0540_),
    .A2(_0577_));
 sg13g2_nand3_1 _1622_ (.B(_0575_),
    .C(_0578_),
    .A(_0539_),
    .Y(_0613_));
 sg13g2_nor2_2 _1623_ (.A(net98),
    .B(_0579_),
    .Y(_0614_));
 sg13g2_nand3b_1 _1624_ (.B(_0611_),
    .C(_0614_),
    .Y(_0615_),
    .A_N(net88));
 sg13g2_nand4_1 _1625_ (.B(_0575_),
    .C(_0579_),
    .A(net99),
    .Y(_0616_),
    .D(net88));
 sg13g2_nand3b_1 _1626_ (.B(_0615_),
    .C(_0616_),
    .Y(_0617_),
    .A_N(_0610_));
 sg13g2_nand3_1 _1627_ (.B(_0582_),
    .C(_0591_),
    .A(net99),
    .Y(_0618_));
 sg13g2_xor2_1 _1628_ (.B(_0618_),
    .A(_0596_),
    .X(_0619_));
 sg13g2_xor2_1 _1629_ (.B(_0619_),
    .A(_0603_),
    .X(_0621_));
 sg13g2_a21oi_2 _1630_ (.B1(_0621_),
    .Y(_0622_),
    .A2(_0617_),
    .A1(_0605_));
 sg13g2_a21o_2 _1631_ (.A2(_0617_),
    .A1(_0605_),
    .B1(_0621_),
    .X(_0623_));
 sg13g2_o21ai_1 _1632_ (.B1(_0594_),
    .Y(_0624_),
    .A1(_0592_),
    .A2(_0600_));
 sg13g2_xor2_1 _1633_ (.B(_0624_),
    .A(_0590_),
    .X(_0625_));
 sg13g2_inv_1 _1634_ (.Y(_0626_),
    .A(net86));
 sg13g2_nand2_2 _1635_ (.Y(_0627_),
    .A(_0623_),
    .B(net87));
 sg13g2_xnor2_1 _1636_ (.Y(_0628_),
    .A(net88),
    .B(_0614_));
 sg13g2_nor2b_1 _1637_ (.A(_0621_),
    .B_N(_0605_),
    .Y(_0629_));
 sg13g2_o21ai_1 _1638_ (.B1(_0629_),
    .Y(_0630_),
    .A1(_0610_),
    .A2(_0628_));
 sg13g2_nand3b_1 _1639_ (.B(_0623_),
    .C(net86),
    .Y(_0632_),
    .A_N(_0630_));
 sg13g2_nand3_1 _1640_ (.B(net86),
    .C(_0630_),
    .A(_0622_),
    .Y(_0633_));
 sg13g2_and2_1 _1641_ (.A(_0632_),
    .B(_0633_),
    .X(_0634_));
 sg13g2_xnor2_1 _1642_ (.Y(_0635_),
    .A(net88),
    .B(_0634_));
 sg13g2_nor3_1 _1643_ (.A(uo_out[2]),
    .B(uo_out[1]),
    .C(uo_out[0]),
    .Y(_0636_));
 sg13g2_and2_1 _1644_ (.A(_0411_),
    .B(_0636_),
    .X(_0637_));
 sg13g2_nand2_2 _1645_ (.Y(_0638_),
    .A(_0455_),
    .B(_0637_));
 sg13g2_nor2_1 _1646_ (.A(uo_out[5]),
    .B(_0638_),
    .Y(_0639_));
 sg13g2_nor2_1 _1647_ (.A(_0400_),
    .B(_0639_),
    .Y(_0640_));
 sg13g2_xnor2_1 _1648_ (.Y(_0641_),
    .A(uo_out[6]),
    .B(_0640_));
 sg13g2_inv_2 _1649_ (.Y(_0643_),
    .A(_0641_));
 sg13g2_nor2_1 _1650_ (.A(_0400_),
    .B(_0637_),
    .Y(_0644_));
 sg13g2_xnor2_1 _1651_ (.Y(_0645_),
    .A(uo_out[4]),
    .B(_0644_));
 sg13g2_xnor2_1 _1652_ (.Y(_0646_),
    .A(_0641_),
    .B(_0645_));
 sg13g2_nor2_1 _1653_ (.A(_0400_),
    .B(_0636_),
    .Y(_0647_));
 sg13g2_xnor2_1 _1654_ (.Y(_0648_),
    .A(uo_out[3]),
    .B(_0647_));
 sg13g2_xnor2_1 _1655_ (.Y(_0649_),
    .A(_0641_),
    .B(_0648_));
 sg13g2_nand2_1 _1656_ (.Y(_0650_),
    .A(_0646_),
    .B(_0649_));
 sg13g2_o21ai_1 _1657_ (.B1(\u_mac.u_adder.sign_b ),
    .Y(_0651_),
    .A1(uo_out[1]),
    .A2(uo_out[0]));
 sg13g2_xnor2_1 _1658_ (.Y(_0652_),
    .A(_0422_),
    .B(_0651_));
 sg13g2_xnor2_1 _1659_ (.Y(_0654_),
    .A(uo_out[2]),
    .B(_0651_));
 sg13g2_xnor2_1 _1660_ (.Y(_0655_),
    .A(_0641_),
    .B(_0652_));
 sg13g2_nand2_1 _1661_ (.Y(_0656_),
    .A(\u_mac.u_adder.sign_b ),
    .B(uo_out[0]));
 sg13g2_xor2_1 _1662_ (.B(_0656_),
    .A(uo_out[1]),
    .X(_0657_));
 sg13g2_xnor2_1 _1663_ (.Y(_0658_),
    .A(_0641_),
    .B(_0657_));
 sg13g2_and2_1 _1664_ (.A(_0655_),
    .B(_0658_),
    .X(_0659_));
 sg13g2_o21ai_1 _1665_ (.B1(uo_out[5]),
    .Y(_0660_),
    .A1(_0400_),
    .A2(_0638_));
 sg13g2_xnor2_1 _1666_ (.Y(_0661_),
    .A(_0466_),
    .B(_0660_));
 sg13g2_o21ai_1 _1667_ (.B1(_0661_),
    .Y(_0662_),
    .A1(_0650_),
    .A2(_0659_));
 sg13g2_nand3_1 _1668_ (.B(_0641_),
    .C(_0657_),
    .A(uo_out[0]),
    .Y(_0663_));
 sg13g2_nand3_1 _1669_ (.B(_0433_),
    .C(_0643_),
    .A(uo_out[1]),
    .Y(_0665_));
 sg13g2_nand3_1 _1670_ (.B(_0663_),
    .C(_0665_),
    .A(_0655_),
    .Y(_0666_));
 sg13g2_nand2_1 _1671_ (.Y(_0667_),
    .A(_0649_),
    .B(_0666_));
 sg13g2_nand2_1 _1672_ (.Y(_0668_),
    .A(_0646_),
    .B(_0667_));
 sg13g2_nand2_1 _1673_ (.Y(_0669_),
    .A(_0661_),
    .B(_0668_));
 sg13g2_nor2_1 _1674_ (.A(_0662_),
    .B(_0668_),
    .Y(_0670_));
 sg13g2_xor2_1 _1675_ (.B(net93),
    .A(_0662_),
    .X(_0671_));
 sg13g2_xnor2_1 _1676_ (.Y(_0672_),
    .A(_0643_),
    .B(_0671_));
 sg13g2_inv_1 _1677_ (.Y(_0673_),
    .A(_0672_));
 sg13g2_nand2_1 _1678_ (.Y(_0674_),
    .A(_0635_),
    .B(_0672_));
 sg13g2_xnor2_1 _1679_ (.Y(_0676_),
    .A(_0635_),
    .B(_0672_));
 sg13g2_xnor2_1 _1680_ (.Y(_0677_),
    .A(_0635_),
    .B(_0673_));
 sg13g2_nor2_1 _1681_ (.A(net88),
    .B(_0627_),
    .Y(_0678_));
 sg13g2_nor2b_2 _1682_ (.A(_0601_),
    .B_N(_0603_),
    .Y(_0679_));
 sg13g2_inv_1 _1683_ (.Y(_0680_),
    .A(_0679_));
 sg13g2_a21oi_2 _1684_ (.B1(_0678_),
    .Y(_0681_),
    .A2(_0679_),
    .A1(_0627_));
 sg13g2_nor3_2 _1685_ (.A(uo_out[5]),
    .B(uo_out[6]),
    .C(_0638_),
    .Y(_0682_));
 sg13g2_nand2_2 _1686_ (.Y(_0683_),
    .A(_0466_),
    .B(_0639_));
 sg13g2_nand2_1 _1687_ (.Y(_0684_),
    .A(_0641_),
    .B(_0683_));
 sg13g2_nand2_1 _1688_ (.Y(_0685_),
    .A(net93),
    .B(_0684_));
 sg13g2_o21ai_1 _1689_ (.B1(_0685_),
    .Y(_0687_),
    .A1(_0643_),
    .A2(net93));
 sg13g2_inv_2 _1690_ (.Y(_0688_),
    .A(_0687_));
 sg13g2_nor2_1 _1691_ (.A(_0681_),
    .B(_0688_),
    .Y(_0689_));
 sg13g2_nand2b_1 _1692_ (.Y(_0690_),
    .B(_0687_),
    .A_N(_0681_));
 sg13g2_nor2_2 _1693_ (.A(_0621_),
    .B(_0626_),
    .Y(_0691_));
 sg13g2_inv_2 _1694_ (.Y(_0692_),
    .A(_0691_));
 sg13g2_o21ai_1 _1695_ (.B1(_0614_),
    .Y(_0693_),
    .A1(_0622_),
    .A2(_0626_));
 sg13g2_nand4_1 _1696_ (.B(_0575_),
    .C(_0623_),
    .A(net99),
    .Y(_0694_),
    .D(net87));
 sg13g2_and2_1 _1697_ (.A(_0693_),
    .B(_0694_),
    .X(_0695_));
 sg13g2_a21oi_1 _1698_ (.A1(_0634_),
    .A2(_0695_),
    .Y(_0696_),
    .B1(_0691_));
 sg13g2_a21o_2 _1699_ (.A2(_0695_),
    .A1(_0634_),
    .B1(_0691_),
    .X(_0698_));
 sg13g2_nand3_1 _1700_ (.B(_0649_),
    .C(_0661_),
    .A(_0646_),
    .Y(_0699_));
 sg13g2_o21ai_1 _1701_ (.B1(_0699_),
    .Y(_0700_),
    .A1(_0662_),
    .A2(_0668_));
 sg13g2_inv_1 _1702_ (.Y(_0701_),
    .A(_0700_));
 sg13g2_nand2_1 _1703_ (.Y(_0702_),
    .A(_0657_),
    .B(net93));
 sg13g2_o21ai_1 _1704_ (.B1(_0702_),
    .Y(_0703_),
    .A1(uo_out[0]),
    .A2(net93));
 sg13g2_inv_1 _1705_ (.Y(_0704_),
    .A(_0703_));
 sg13g2_nor2_2 _1706_ (.A(_0700_),
    .B(_0703_),
    .Y(_0705_));
 sg13g2_inv_1 _1707_ (.Y(_0706_),
    .A(_0705_));
 sg13g2_nand2_1 _1708_ (.Y(_0707_),
    .A(_0698_),
    .B(_0705_));
 sg13g2_mux2_1 _1709_ (.A0(_0614_),
    .A1(_0608_),
    .S(_0627_),
    .X(_0709_));
 sg13g2_a21oi_1 _1710_ (.A1(_0623_),
    .A2(net86),
    .Y(_0710_),
    .B1(_0611_));
 sg13g2_mux2_1 _1711_ (.A0(_0709_),
    .A1(_0710_),
    .S(_0634_),
    .X(_0711_));
 sg13g2_and2_1 _1712_ (.A(_0692_),
    .B(_0711_),
    .X(_0712_));
 sg13g2_nand2_1 _1713_ (.Y(_0713_),
    .A(_0654_),
    .B(net93));
 sg13g2_o21ai_1 _1714_ (.B1(_0713_),
    .Y(_0714_),
    .A1(_0657_),
    .A2(net94));
 sg13g2_nand2_1 _1715_ (.Y(_0715_),
    .A(_0671_),
    .B(_0714_));
 sg13g2_nand3_1 _1716_ (.B(_0662_),
    .C(net93),
    .A(uo_out[0]),
    .Y(_0716_));
 sg13g2_nand2_1 _1717_ (.Y(_0717_),
    .A(_0715_),
    .B(_0716_));
 sg13g2_a21oi_1 _1718_ (.A1(_0715_),
    .A2(_0716_),
    .Y(_0718_),
    .B1(_0700_));
 sg13g2_inv_1 _1719_ (.Y(_0720_),
    .A(_0718_));
 sg13g2_a21o_1 _1720_ (.A2(_0711_),
    .A1(_0692_),
    .B1(_0720_),
    .X(_0721_));
 sg13g2_nand3_1 _1721_ (.B(_0623_),
    .C(net87),
    .A(_0604_),
    .Y(_0722_));
 sg13g2_a21o_1 _1722_ (.A2(net86),
    .A1(_0623_),
    .B1(_0619_),
    .X(_0723_));
 sg13g2_a22oi_1 _1723_ (.Y(_0724_),
    .B1(_0722_),
    .B2(_0723_),
    .A2(_0633_),
    .A1(_0632_));
 sg13g2_and4_1 _1724_ (.A(_0605_),
    .B(_0622_),
    .C(net86),
    .D(_0630_),
    .X(_0725_));
 sg13g2_nand2b_1 _1725_ (.Y(_0726_),
    .B(_0605_),
    .A_N(_0633_));
 sg13g2_nor2_1 _1726_ (.A(_0692_),
    .B(_0725_),
    .Y(_0727_));
 sg13g2_a221oi_1 _1727_ (.B2(_0691_),
    .C1(_0724_),
    .B1(_0726_),
    .A1(_0634_),
    .Y(_0728_),
    .A2(_0709_));
 sg13g2_or3_1 _1728_ (.A(_0605_),
    .B(_0611_),
    .C(_0633_),
    .X(_0729_));
 sg13g2_a21oi_2 _1729_ (.B1(_0728_),
    .Y(_0731_),
    .A2(_0729_),
    .A1(_0691_));
 sg13g2_a21o_1 _1730_ (.A2(_0729_),
    .A1(_0691_),
    .B1(_0728_),
    .X(_0732_));
 sg13g2_a21oi_2 _1731_ (.B1(_0701_),
    .Y(_0733_),
    .A2(_0670_),
    .A1(_0649_));
 sg13g2_a21o_1 _1732_ (.A2(_0699_),
    .A1(uo_out[0]),
    .B1(_0701_),
    .X(_0734_));
 sg13g2_o21ai_1 _1733_ (.B1(_0734_),
    .Y(_0735_),
    .A1(_0714_),
    .A2(_0733_));
 sg13g2_inv_1 _1734_ (.Y(_0736_),
    .A(_0735_));
 sg13g2_nor2_1 _1735_ (.A(_0698_),
    .B(_0705_),
    .Y(_0737_));
 sg13g2_a221oi_1 _1736_ (.B2(_0735_),
    .C1(_0737_),
    .B1(_0731_),
    .A1(_0707_),
    .Y(_0738_),
    .A2(_0721_));
 sg13g2_a21oi_1 _1737_ (.A1(_0648_),
    .A2(net94),
    .Y(_0739_),
    .B1(_0700_));
 sg13g2_o21ai_1 _1738_ (.B1(_0739_),
    .Y(_0740_),
    .A1(_0654_),
    .A2(net94));
 sg13g2_nand3_1 _1739_ (.B(_0704_),
    .C(_0733_),
    .A(_0671_),
    .Y(_0742_));
 sg13g2_nand2_2 _1740_ (.Y(_0743_),
    .A(_0740_),
    .B(_0742_));
 sg13g2_inv_1 _1741_ (.Y(_0744_),
    .A(_0743_));
 sg13g2_a221oi_1 _1742_ (.B2(_0694_),
    .C1(_0725_),
    .B1(_0693_),
    .A1(_0632_),
    .Y(_0745_),
    .A2(_0633_));
 sg13g2_nor2_1 _1743_ (.A(_0692_),
    .B(_0745_),
    .Y(_0746_));
 sg13g2_nand3_1 _1744_ (.B(_0623_),
    .C(net86),
    .A(_0608_),
    .Y(_0747_));
 sg13g2_o21ai_1 _1745_ (.B1(_0604_),
    .Y(_0748_),
    .A1(_0622_),
    .A2(_0626_));
 sg13g2_nand4_1 _1746_ (.B(_0633_),
    .C(_0747_),
    .A(_0632_),
    .Y(_0749_),
    .D(_0748_));
 sg13g2_nor2b_2 _1747_ (.A(_0746_),
    .B_N(_0749_),
    .Y(_0750_));
 sg13g2_o21ai_1 _1748_ (.B1(_0749_),
    .Y(_0751_),
    .A1(_0692_),
    .A2(_0745_));
 sg13g2_nand2_1 _1749_ (.Y(_0753_),
    .A(_0743_),
    .B(_0751_));
 sg13g2_o21ai_1 _1750_ (.B1(_0753_),
    .Y(_0754_),
    .A1(_0731_),
    .A2(_0735_));
 sg13g2_and2_1 _1751_ (.A(_0717_),
    .B(_0733_),
    .X(_0755_));
 sg13g2_nand2_1 _1752_ (.Y(_0756_),
    .A(_0645_),
    .B(net93));
 sg13g2_nor2b_1 _1753_ (.A(net94),
    .B_N(_0648_),
    .Y(_0757_));
 sg13g2_nor2_1 _1754_ (.A(_0700_),
    .B(_0757_),
    .Y(_0758_));
 sg13g2_a22oi_1 _1755_ (.Y(_0759_),
    .B1(_0756_),
    .B2(_0758_),
    .A2(_0733_),
    .A1(_0717_));
 sg13g2_a21o_2 _1756_ (.A2(_0758_),
    .A1(_0756_),
    .B1(_0755_),
    .X(_0760_));
 sg13g2_nand4_1 _1757_ (.B(_0633_),
    .C(_0722_),
    .A(_0632_),
    .Y(_0761_),
    .D(_0723_));
 sg13g2_and2_1 _1758_ (.A(_0692_),
    .B(_0761_),
    .X(_0762_));
 sg13g2_a21oi_2 _1759_ (.B1(_0762_),
    .Y(_0764_),
    .A2(_0727_),
    .A1(_0711_));
 sg13g2_a21o_1 _1760_ (.A2(_0727_),
    .A1(_0711_),
    .B1(_0762_),
    .X(_0765_));
 sg13g2_a22oi_1 _1761_ (.Y(_0766_),
    .B1(_0759_),
    .B2(_0765_),
    .A2(_0750_),
    .A1(_0744_));
 sg13g2_o21ai_1 _1762_ (.B1(_0766_),
    .Y(_0767_),
    .A1(_0738_),
    .A2(_0754_));
 sg13g2_a22oi_1 _1763_ (.Y(_0768_),
    .B1(_0760_),
    .B2(_0764_),
    .A2(_0683_),
    .A1(net97));
 sg13g2_nand3_1 _1764_ (.B(_0629_),
    .C(_0632_),
    .A(net86),
    .Y(_0769_));
 sg13g2_mux2_1 _1765_ (.A0(net88),
    .A1(_0680_),
    .S(_0769_),
    .X(_0770_));
 sg13g2_mux2_1 _1766_ (.A0(_0652_),
    .A1(_0643_),
    .S(_0699_),
    .X(_0771_));
 sg13g2_nor2_1 _1767_ (.A(_0770_),
    .B(_0771_),
    .Y(_0772_));
 sg13g2_xnor2_1 _1768_ (.Y(_0773_),
    .A(_0770_),
    .B(_0771_));
 sg13g2_inv_1 _1769_ (.Y(_0775_),
    .A(_0773_));
 sg13g2_or2_1 _1770_ (.X(_0776_),
    .B(_0684_),
    .A(_0679_));
 sg13g2_nand2_1 _1771_ (.Y(_0777_),
    .A(_0679_),
    .B(_0684_));
 sg13g2_and2_1 _1772_ (.A(_0776_),
    .B(_0777_),
    .X(_0778_));
 sg13g2_nand3_1 _1773_ (.B(_0773_),
    .C(_0778_),
    .A(_0676_),
    .Y(_0779_));
 sg13g2_nor2_1 _1774_ (.A(net97),
    .B(_0683_),
    .Y(_0780_));
 sg13g2_nand2_2 _1775_ (.Y(_0781_),
    .A(_0681_),
    .B(_0688_));
 sg13g2_inv_1 _1776_ (.Y(_0782_),
    .A(_0781_));
 sg13g2_nand2_2 _1777_ (.Y(_0783_),
    .A(_0690_),
    .B(_0781_));
 sg13g2_nand2b_1 _1778_ (.Y(_0784_),
    .B(_0781_),
    .A_N(_0779_));
 sg13g2_or3_1 _1779_ (.A(_0779_),
    .B(_0780_),
    .C(net85),
    .X(_0786_));
 sg13g2_a21oi_1 _1780_ (.A1(_0767_),
    .A2(_0768_),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_a21o_2 _1781_ (.A2(_0768_),
    .A1(_0767_),
    .B1(_0786_),
    .X(_0788_));
 sg13g2_nand4_1 _1782_ (.B(_0673_),
    .C(_0773_),
    .A(_0635_),
    .Y(_0789_),
    .D(_0778_));
 sg13g2_nand3b_1 _1783_ (.B(_0771_),
    .C(_0777_),
    .Y(_0790_),
    .A_N(_0770_));
 sg13g2_and4_1 _1784_ (.A(_0776_),
    .B(_0784_),
    .C(_0789_),
    .D(_0790_),
    .X(_0791_));
 sg13g2_nand4_1 _1785_ (.B(_0784_),
    .C(_0789_),
    .A(_0776_),
    .Y(_0792_),
    .D(_0790_));
 sg13g2_nand2_2 _1786_ (.Y(_0793_),
    .A(_0788_),
    .B(_0792_));
 sg13g2_a21oi_1 _1787_ (.A1(_0788_),
    .A2(_0792_),
    .Y(_0794_),
    .B1(_0689_));
 sg13g2_o21ai_1 _1788_ (.B1(_0690_),
    .Y(_0795_),
    .A1(_0787_),
    .A2(_0791_));
 sg13g2_nor3_1 _1789_ (.A(_0782_),
    .B(_0787_),
    .C(_0791_),
    .Y(_0797_));
 sg13g2_nand3_1 _1790_ (.B(_0788_),
    .C(_0792_),
    .A(_0781_),
    .Y(_0798_));
 sg13g2_a21oi_2 _1791_ (.B1(_0677_),
    .Y(_0799_),
    .A2(_0798_),
    .A1(_0795_));
 sg13g2_o21ai_1 _1792_ (.B1(_0676_),
    .Y(_0800_),
    .A1(_0794_),
    .A2(_0797_));
 sg13g2_nor3_2 _1793_ (.A(_0676_),
    .B(_0794_),
    .C(_0797_),
    .Y(_0801_));
 sg13g2_nand3_1 _1794_ (.B(_0795_),
    .C(_0798_),
    .A(_0677_),
    .Y(_0802_));
 sg13g2_nor2_2 _1795_ (.A(_0799_),
    .B(_0801_),
    .Y(_0803_));
 sg13g2_mux2_1 _1796_ (.A0(_0682_),
    .A1(net97),
    .S(net83),
    .X(_0804_));
 sg13g2_nor2_1 _1797_ (.A(net85),
    .B(_0804_),
    .Y(_0805_));
 sg13g2_nor4_1 _1798_ (.A(_0677_),
    .B(_0689_),
    .C(_0782_),
    .D(_0804_),
    .Y(_0806_));
 sg13g2_nand3b_1 _1799_ (.B(_0788_),
    .C(_0792_),
    .Y(_0808_),
    .A_N(_0635_));
 sg13g2_o21ai_1 _1800_ (.B1(_0673_),
    .Y(_0809_),
    .A1(_0787_),
    .A2(_0791_));
 sg13g2_and2_1 _1801_ (.A(_0808_),
    .B(_0809_),
    .X(_0810_));
 sg13g2_and3_1 _1802_ (.X(_0811_),
    .A(_0674_),
    .B(_0808_),
    .C(_0809_));
 sg13g2_nand3_1 _1803_ (.B(_0808_),
    .C(_0809_),
    .A(_0674_),
    .Y(_0812_));
 sg13g2_o21ai_1 _1804_ (.B1(_0773_),
    .Y(_0813_),
    .A1(_0799_),
    .A2(_0811_));
 sg13g2_nand3_1 _1805_ (.B(_0800_),
    .C(_0812_),
    .A(_0775_),
    .Y(_0814_));
 sg13g2_o21ai_1 _1806_ (.B1(_0775_),
    .Y(_0815_),
    .A1(_0799_),
    .A2(_0811_));
 sg13g2_nand3_1 _1807_ (.B(_0800_),
    .C(_0812_),
    .A(_0773_),
    .Y(_0816_));
 sg13g2_nand2_2 _1808_ (.Y(_0817_),
    .A(_0813_),
    .B(_0814_));
 sg13g2_mux2_1 _1809_ (.A0(_0770_),
    .A1(_0771_),
    .S(net84),
    .X(_0819_));
 sg13g2_or2_1 _1810_ (.X(_0820_),
    .B(_0819_),
    .A(_0772_));
 sg13g2_a21o_2 _1811_ (.A2(_0820_),
    .A1(_0813_),
    .B1(_0778_),
    .X(_0821_));
 sg13g2_and2_1 _1812_ (.A(net79),
    .B(_0821_),
    .X(_0822_));
 sg13g2_nand2_1 _1813_ (.Y(_0823_),
    .A(_0806_),
    .B(net78));
 sg13g2_mux4_1 _1814_ (.S0(net83),
    .A0(_0759_),
    .A1(_0764_),
    .A2(_0682_),
    .A3(net97),
    .S1(_0783_),
    .X(_0824_));
 sg13g2_nor2_2 _1815_ (.A(_0803_),
    .B(_0824_),
    .Y(_0825_));
 sg13g2_nand2_1 _1816_ (.Y(_0826_),
    .A(net79),
    .B(_0825_));
 sg13g2_and2_1 _1817_ (.A(net78),
    .B(_0825_),
    .X(_0827_));
 sg13g2_inv_1 _1818_ (.Y(_0828_),
    .A(_0827_));
 sg13g2_nand2_1 _1819_ (.Y(_0830_),
    .A(_0760_),
    .B(net84));
 sg13g2_o21ai_1 _1820_ (.B1(_0830_),
    .Y(_0831_),
    .A1(_0764_),
    .A2(_0793_));
 sg13g2_and2_1 _1821_ (.A(_0827_),
    .B(_0831_),
    .X(_0832_));
 sg13g2_nor2_1 _1822_ (.A(_0828_),
    .B(_0831_),
    .Y(_0833_));
 sg13g2_inv_1 _1823_ (.Y(_0834_),
    .A(_0833_));
 sg13g2_nand2_1 _1824_ (.Y(_0835_),
    .A(_0828_),
    .B(_0831_));
 sg13g2_nor2b_1 _1825_ (.A(_0833_),
    .B_N(_0835_),
    .Y(_0836_));
 sg13g2_inv_1 _1826_ (.Y(_0837_),
    .A(_0836_));
 sg13g2_mux4_1 _1827_ (.S0(net81),
    .A0(_0743_),
    .A1(_0750_),
    .A2(_0760_),
    .A3(_0765_),
    .S1(_0783_),
    .X(_0838_));
 sg13g2_mux2_1 _1828_ (.A0(_0838_),
    .A1(_0805_),
    .S(_0803_),
    .X(_0839_));
 sg13g2_nand2_1 _1829_ (.Y(_0841_),
    .A(net79),
    .B(_0839_));
 sg13g2_nand2_1 _1830_ (.Y(_0842_),
    .A(net78),
    .B(_0839_));
 sg13g2_nand2_1 _1831_ (.Y(_0843_),
    .A(_0743_),
    .B(net82));
 sg13g2_o21ai_1 _1832_ (.B1(_0843_),
    .Y(_0844_),
    .A1(_0751_),
    .A2(net83));
 sg13g2_a21oi_1 _1833_ (.A1(_0822_),
    .A2(_0839_),
    .Y(_0845_),
    .B1(_0844_));
 sg13g2_nand3_1 _1834_ (.B(_0839_),
    .C(_0844_),
    .A(_0822_),
    .Y(_0846_));
 sg13g2_nand3_1 _1835_ (.B(_0802_),
    .C(_0824_),
    .A(_0800_),
    .Y(_0847_));
 sg13g2_mux4_1 _1836_ (.S0(net85),
    .A0(_0735_),
    .A1(_0744_),
    .A2(_0732_),
    .A3(_0751_),
    .S1(net82),
    .X(_0848_));
 sg13g2_mux4_1 _1837_ (.S0(net85),
    .A0(_0736_),
    .A1(_0743_),
    .A2(_0731_),
    .A3(_0750_),
    .S1(net81),
    .X(_0849_));
 sg13g2_o21ai_1 _1838_ (.B1(_0848_),
    .Y(_0850_),
    .A1(_0799_),
    .A2(_0801_));
 sg13g2_and2_1 _1839_ (.A(_0847_),
    .B(_0850_),
    .X(_0852_));
 sg13g2_nand4_1 _1840_ (.B(_0816_),
    .C(_0847_),
    .A(_0815_),
    .Y(_0853_),
    .D(_0850_));
 sg13g2_nand2_1 _1841_ (.Y(_0854_),
    .A(net78),
    .B(_0852_));
 sg13g2_nand2_1 _1842_ (.Y(_0855_),
    .A(_0735_),
    .B(net81));
 sg13g2_o21ai_1 _1843_ (.B1(_0855_),
    .Y(_0856_),
    .A1(_0731_),
    .A2(net81));
 sg13g2_nand2_1 _1844_ (.Y(_0857_),
    .A(_0854_),
    .B(_0856_));
 sg13g2_nor2_1 _1845_ (.A(_0854_),
    .B(_0856_),
    .Y(_0858_));
 sg13g2_nand3b_1 _1846_ (.B(_0802_),
    .C(_0800_),
    .Y(_0859_),
    .A_N(_0838_));
 sg13g2_mux2_1 _1847_ (.A0(_0705_),
    .A1(_0696_),
    .S(net81),
    .X(_0860_));
 sg13g2_mux4_1 _1848_ (.S0(_0783_),
    .A0(_0706_),
    .A1(_0735_),
    .A2(_0698_),
    .A3(_0732_),
    .S1(net82),
    .X(_0861_));
 sg13g2_o21ai_1 _1849_ (.B1(_0861_),
    .Y(_0863_),
    .A1(_0799_),
    .A2(_0801_));
 sg13g2_and2_1 _1850_ (.A(_0859_),
    .B(_0863_),
    .X(_0864_));
 sg13g2_nand4_1 _1851_ (.B(_0816_),
    .C(_0859_),
    .A(_0815_),
    .Y(_0865_),
    .D(_0863_));
 sg13g2_nand3_1 _1852_ (.B(_0813_),
    .C(_0814_),
    .A(_0806_),
    .Y(_0866_));
 sg13g2_nand2_1 _1853_ (.Y(_0867_),
    .A(_0865_),
    .B(_0866_));
 sg13g2_nand2_1 _1854_ (.Y(_0868_),
    .A(_0821_),
    .B(_0867_));
 sg13g2_nor2_1 _1855_ (.A(_0696_),
    .B(net81),
    .Y(_0869_));
 sg13g2_a21oi_1 _1856_ (.A1(_0706_),
    .A2(net81),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_a21oi_1 _1857_ (.A1(_0821_),
    .A2(_0867_),
    .Y(_0871_),
    .B1(_0870_));
 sg13g2_nand3_1 _1858_ (.B(_0867_),
    .C(_0870_),
    .A(_0821_),
    .Y(_0872_));
 sg13g2_mux2_1 _1859_ (.A0(_0718_),
    .A1(_0712_),
    .S(net81),
    .X(_0874_));
 sg13g2_mux2_1 _1860_ (.A0(_0874_),
    .A1(_0860_),
    .S(net85),
    .X(_0875_));
 sg13g2_mux2_1 _1861_ (.A0(_0875_),
    .A1(_0849_),
    .S(_0803_),
    .X(_0876_));
 sg13g2_mux2_1 _1862_ (.A0(_0825_),
    .A1(_0876_),
    .S(net79),
    .X(_0877_));
 sg13g2_nor2_1 _1863_ (.A(_0712_),
    .B(net82),
    .Y(_0878_));
 sg13g2_a21oi_2 _1864_ (.B1(_0878_),
    .Y(_0879_),
    .A2(net82),
    .A1(_0720_));
 sg13g2_nand2_1 _1865_ (.Y(_0880_),
    .A(_0877_),
    .B(_0879_));
 sg13g2_o21ai_1 _1866_ (.B1(_0872_),
    .Y(_0881_),
    .A1(_0871_),
    .A2(_0880_));
 sg13g2_a21oi_1 _1867_ (.A1(_0857_),
    .A2(_0881_),
    .Y(_0882_),
    .B1(_0858_));
 sg13g2_o21ai_1 _1868_ (.B1(_0846_),
    .Y(_0883_),
    .A1(_0845_),
    .A2(_0882_));
 sg13g2_a21oi_1 _1869_ (.A1(_0837_),
    .A2(_0883_),
    .Y(_0885_),
    .B1(_0832_));
 sg13g2_xnor2_1 _1870_ (.Y(_0886_),
    .A(_0400_),
    .B(_0591_));
 sg13g2_xnor2_1 _1871_ (.Y(_0887_),
    .A(\u_mac.u_adder.sign_b ),
    .B(_0591_));
 sg13g2_nor2_1 _1872_ (.A(_0587_),
    .B(net84),
    .Y(_0888_));
 sg13g2_a21oi_1 _1873_ (.A1(_0823_),
    .A2(_0885_),
    .Y(_0889_),
    .B1(_0886_));
 sg13g2_a221oi_1 _1874_ (.B2(net78),
    .C1(_0888_),
    .B1(_0806_),
    .A1(_0682_),
    .Y(_0890_),
    .A2(net84));
 sg13g2_and2_1 _1875_ (.A(_0842_),
    .B(_0844_),
    .X(_0891_));
 sg13g2_nand2b_1 _1876_ (.Y(_0892_),
    .B(_0846_),
    .A_N(_0845_));
 sg13g2_inv_1 _1877_ (.Y(_0893_),
    .A(_0892_));
 sg13g2_a21oi_1 _1878_ (.A1(net78),
    .A2(_0852_),
    .Y(_0894_),
    .B1(_0856_));
 sg13g2_inv_1 _1879_ (.Y(_0896_),
    .A(_0894_));
 sg13g2_and2_1 _1880_ (.A(_0868_),
    .B(_0870_),
    .X(_0897_));
 sg13g2_nor2b_1 _1881_ (.A(_0871_),
    .B_N(_0872_),
    .Y(_0898_));
 sg13g2_nand2b_1 _1882_ (.Y(_0899_),
    .B(_0879_),
    .A_N(_0877_));
 sg13g2_a21oi_1 _1883_ (.A1(_0821_),
    .A2(_0864_),
    .Y(_0900_),
    .B1(net80));
 sg13g2_or4_1 _1884_ (.A(net85),
    .B(_0803_),
    .C(_0804_),
    .D(_0821_),
    .X(_0901_));
 sg13g2_nand2_1 _1885_ (.Y(_0902_),
    .A(net85),
    .B(_0874_));
 sg13g2_nand3_1 _1886_ (.B(_0803_),
    .C(_0874_),
    .A(net85),
    .Y(_0903_));
 sg13g2_and2_1 _1887_ (.A(net80),
    .B(_0903_),
    .X(_0904_));
 sg13g2_a21oi_2 _1888_ (.B1(_0900_),
    .Y(_0905_),
    .A2(_0904_),
    .A1(_0901_));
 sg13g2_nand2b_1 _1889_ (.Y(_0907_),
    .B(_0876_),
    .A_N(net79));
 sg13g2_a21oi_2 _1890_ (.B1(net78),
    .Y(_0908_),
    .A2(_0907_),
    .A1(_0826_));
 sg13g2_a21oi_1 _1891_ (.A1(_0865_),
    .A2(_0866_),
    .Y(_0909_),
    .B1(_0821_));
 sg13g2_nor2_1 _1892_ (.A(net79),
    .B(_0903_),
    .Y(_0910_));
 sg13g2_nor2_1 _1893_ (.A(_0909_),
    .B(_0910_),
    .Y(_0911_));
 sg13g2_nand2_1 _1894_ (.Y(_0912_),
    .A(_0803_),
    .B(_0875_));
 sg13g2_a22oi_1 _1895_ (.Y(_0913_),
    .B1(_0853_),
    .B2(_0912_),
    .A2(_0821_),
    .A1(net80));
 sg13g2_nor3_1 _1896_ (.A(_0909_),
    .B(_0910_),
    .C(_0913_),
    .Y(_0914_));
 sg13g2_or3_1 _1897_ (.A(_0909_),
    .B(_0910_),
    .C(_0913_),
    .X(_0915_));
 sg13g2_mux2_1 _1898_ (.A0(_0902_),
    .A1(_0861_),
    .S(_0803_),
    .X(_0916_));
 sg13g2_a21oi_2 _1899_ (.B1(net78),
    .Y(_0918_),
    .A2(_0916_),
    .A1(_0841_));
 sg13g2_nand2b_1 _1900_ (.Y(_0919_),
    .B(_0914_),
    .A_N(_0918_));
 sg13g2_nor2_1 _1901_ (.A(_0908_),
    .B(_0919_),
    .Y(_0920_));
 sg13g2_nand2_1 _1902_ (.Y(_0921_),
    .A(_0886_),
    .B(_0919_));
 sg13g2_xnor2_1 _1903_ (.Y(_0922_),
    .A(_0908_),
    .B(_0921_));
 sg13g2_nor2_1 _1904_ (.A(_0887_),
    .B(_0914_),
    .Y(_0923_));
 sg13g2_xnor2_1 _1905_ (.Y(_0924_),
    .A(_0918_),
    .B(_0923_));
 sg13g2_xor2_1 _1906_ (.B(_0923_),
    .A(_0918_),
    .X(_0925_));
 sg13g2_nor2_1 _1907_ (.A(_0887_),
    .B(_0920_),
    .Y(_0926_));
 sg13g2_xor2_1 _1908_ (.B(_0926_),
    .A(_0905_),
    .X(_0927_));
 sg13g2_xnor2_1 _1909_ (.Y(_0929_),
    .A(_0905_),
    .B(_0926_));
 sg13g2_nor4_2 _1910_ (.A(_0905_),
    .B(_0908_),
    .C(_0915_),
    .Y(_0930_),
    .D(_0918_));
 sg13g2_nand2_1 _1911_ (.Y(_0931_),
    .A(net80),
    .B(_0912_));
 sg13g2_o21ai_1 _1912_ (.B1(_0931_),
    .Y(_0932_),
    .A1(net80),
    .A2(_0852_));
 sg13g2_nor2_1 _1913_ (.A(net79),
    .B(_0839_),
    .Y(_0933_));
 sg13g2_a21oi_1 _1914_ (.A1(net79),
    .A2(_0916_),
    .Y(_0934_),
    .B1(_0933_));
 sg13g2_inv_2 _1915_ (.Y(_0935_),
    .A(_0934_));
 sg13g2_and3_1 _1916_ (.X(_0936_),
    .A(_0930_),
    .B(_0932_),
    .C(_0935_));
 sg13g2_xnor2_1 _1917_ (.Y(_0937_),
    .A(_0877_),
    .B(_0879_));
 sg13g2_nand4_1 _1918_ (.B(_0932_),
    .C(_0935_),
    .A(_0930_),
    .Y(_0938_),
    .D(_0937_));
 sg13g2_nand2_1 _1919_ (.Y(_0940_),
    .A(_0899_),
    .B(_0938_));
 sg13g2_a21oi_1 _1920_ (.A1(_0899_),
    .A2(_0938_),
    .Y(_0941_),
    .B1(_0898_));
 sg13g2_or2_1 _1921_ (.X(_0942_),
    .B(_0941_),
    .A(_0897_));
 sg13g2_xnor2_1 _1922_ (.Y(_0943_),
    .A(_0854_),
    .B(_0856_));
 sg13g2_o21ai_1 _1923_ (.B1(_0943_),
    .Y(_0944_),
    .A1(_0897_),
    .A2(_0941_));
 sg13g2_nand2_1 _1924_ (.Y(_0945_),
    .A(_0896_),
    .B(_0944_));
 sg13g2_a21oi_1 _1925_ (.A1(_0896_),
    .A2(_0944_),
    .Y(_0946_),
    .B1(_0893_));
 sg13g2_nor2_1 _1926_ (.A(_0891_),
    .B(_0946_),
    .Y(_0947_));
 sg13g2_o21ai_1 _1927_ (.B1(_0834_),
    .Y(_0948_),
    .A1(_0891_),
    .A2(_0946_));
 sg13g2_a21oi_1 _1928_ (.A1(_0828_),
    .A2(_0831_),
    .Y(_0949_),
    .B1(_0887_));
 sg13g2_nand2_1 _1929_ (.Y(_0951_),
    .A(_0835_),
    .B(_0948_));
 sg13g2_nor3_1 _1930_ (.A(_0887_),
    .B(_0890_),
    .C(_0951_),
    .Y(_0952_));
 sg13g2_or2_1 _1931_ (.X(_0953_),
    .B(_0952_),
    .A(_0889_));
 sg13g2_mux2_1 _1932_ (.A0(_0880_),
    .A1(_0940_),
    .S(_0886_),
    .X(_0954_));
 sg13g2_xnor2_1 _1933_ (.Y(_0955_),
    .A(_0898_),
    .B(_0954_));
 sg13g2_inv_1 _1934_ (.Y(_0956_),
    .A(_0955_));
 sg13g2_nor2_1 _1935_ (.A(_0887_),
    .B(_0936_),
    .Y(_0957_));
 sg13g2_xnor2_1 _1936_ (.Y(_0958_),
    .A(_0937_),
    .B(_0957_));
 sg13g2_inv_1 _1937_ (.Y(_0959_),
    .A(_0958_));
 sg13g2_nor2_1 _1938_ (.A(_0955_),
    .B(_0958_),
    .Y(_0960_));
 sg13g2_a21oi_1 _1939_ (.A1(_0930_),
    .A2(_0932_),
    .Y(_0962_),
    .B1(_0887_));
 sg13g2_xnor2_1 _1940_ (.Y(_0963_),
    .A(_0935_),
    .B(_0962_));
 sg13g2_nor2_1 _1941_ (.A(_0887_),
    .B(_0930_),
    .Y(_0964_));
 sg13g2_xnor2_1 _1942_ (.Y(_0965_),
    .A(_0932_),
    .B(_0964_));
 sg13g2_or2_1 _1943_ (.X(_0966_),
    .B(_0965_),
    .A(_0963_));
 sg13g2_or3_1 _1944_ (.A(_0955_),
    .B(_0958_),
    .C(_0966_),
    .X(_0967_));
 sg13g2_nor2_1 _1945_ (.A(_0885_),
    .B(_0886_),
    .Y(_0968_));
 sg13g2_a21oi_1 _1946_ (.A1(_0948_),
    .A2(_0949_),
    .Y(_0969_),
    .B1(_0968_));
 sg13g2_nor2_1 _1947_ (.A(_0890_),
    .B(_0969_),
    .Y(_0970_));
 sg13g2_xor2_1 _1948_ (.B(_0969_),
    .A(_0890_),
    .X(_0971_));
 sg13g2_mux2_1 _1949_ (.A0(_0883_),
    .A1(_0947_),
    .S(_0886_),
    .X(_0973_));
 sg13g2_xnor2_1 _1950_ (.Y(_0974_),
    .A(_0836_),
    .B(_0973_));
 sg13g2_xnor2_1 _1951_ (.Y(_0975_),
    .A(_0837_),
    .B(_0973_));
 sg13g2_mux2_1 _1952_ (.A0(_0882_),
    .A1(_0945_),
    .S(_0886_),
    .X(_0976_));
 sg13g2_xnor2_1 _1953_ (.Y(_0977_),
    .A(_0893_),
    .B(_0976_));
 sg13g2_xnor2_1 _1954_ (.Y(_0978_),
    .A(_0892_),
    .B(_0976_));
 sg13g2_nor2_1 _1955_ (.A(_0881_),
    .B(_0886_),
    .Y(_0979_));
 sg13g2_a21oi_1 _1956_ (.A1(_0886_),
    .A2(_0942_),
    .Y(_0980_),
    .B1(_0979_));
 sg13g2_xnor2_1 _1957_ (.Y(_0981_),
    .A(_0943_),
    .B(_0980_));
 sg13g2_inv_2 _1958_ (.Y(_0982_),
    .A(_0981_));
 sg13g2_nand4_1 _1959_ (.B(_0975_),
    .C(_0978_),
    .A(_0971_),
    .Y(_0984_),
    .D(_0982_));
 sg13g2_nor2_1 _1960_ (.A(_0967_),
    .B(_0984_),
    .Y(_0985_));
 sg13g2_and2_1 _1961_ (.A(_0930_),
    .B(_0985_),
    .X(_0986_));
 sg13g2_nor2_1 _1962_ (.A(_0681_),
    .B(net84),
    .Y(_0987_));
 sg13g2_a21oi_2 _1963_ (.B1(_0987_),
    .Y(_0988_),
    .A2(net84),
    .A1(_0688_));
 sg13g2_inv_1 _1964_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_nand2_1 _1965_ (.Y(_0990_),
    .A(_0810_),
    .B(_0989_));
 sg13g2_nor2_1 _1966_ (.A(_0819_),
    .B(_0990_),
    .Y(_0991_));
 sg13g2_xor2_1 _1967_ (.B(_0990_),
    .A(_0819_),
    .X(_0992_));
 sg13g2_nor2_1 _1968_ (.A(_0887_),
    .B(_0911_),
    .Y(_0993_));
 sg13g2_xor2_1 _1969_ (.B(_0993_),
    .A(_0913_),
    .X(_0995_));
 sg13g2_nor2_1 _1970_ (.A(_0925_),
    .B(_0995_),
    .Y(_0996_));
 sg13g2_nor3_1 _1971_ (.A(_0922_),
    .B(_0927_),
    .C(_0996_),
    .Y(_0997_));
 sg13g2_o21ai_1 _1972_ (.B1(_0960_),
    .Y(_0998_),
    .A1(_0966_),
    .A2(_0997_));
 sg13g2_nand3_1 _1973_ (.B(_0982_),
    .C(_0998_),
    .A(_0978_),
    .Y(_0999_));
 sg13g2_nand3_1 _1974_ (.B(_0975_),
    .C(_0999_),
    .A(_0971_),
    .Y(_1000_));
 sg13g2_inv_2 _1975_ (.Y(_1001_),
    .A(_1000_));
 sg13g2_and2_1 _1976_ (.A(_0810_),
    .B(_1000_),
    .X(_1002_));
 sg13g2_a21o_1 _1977_ (.A2(_0995_),
    .A1(_0924_),
    .B1(_0922_),
    .X(_1003_));
 sg13g2_a21oi_1 _1978_ (.A1(_0929_),
    .A2(_1003_),
    .Y(_1004_),
    .B1(_0965_));
 sg13g2_o21ai_1 _1979_ (.B1(_0959_),
    .Y(_1006_),
    .A1(_0963_),
    .A2(_1004_));
 sg13g2_a21oi_1 _1980_ (.A1(_0956_),
    .A2(_1006_),
    .Y(_1007_),
    .B1(_0981_));
 sg13g2_nor2_1 _1981_ (.A(_0977_),
    .B(_1007_),
    .Y(_1008_));
 sg13g2_o21ai_1 _1982_ (.B1(_0971_),
    .Y(_1009_),
    .A1(_0974_),
    .A2(_1008_));
 sg13g2_nand2b_2 _1983_ (.Y(_1010_),
    .B(_0988_),
    .A_N(_1009_));
 sg13g2_xor2_1 _1984_ (.B(_1000_),
    .A(_0810_),
    .X(_1011_));
 sg13g2_a21oi_1 _1985_ (.A1(_1010_),
    .A2(_1011_),
    .Y(_1012_),
    .B1(_1002_));
 sg13g2_nor3_1 _1986_ (.A(_0911_),
    .B(_0922_),
    .C(_0927_),
    .Y(_1013_));
 sg13g2_a21oi_1 _1987_ (.A1(_0996_),
    .A2(_1013_),
    .Y(_1014_),
    .B1(_0967_));
 sg13g2_nor2_2 _1988_ (.A(_0984_),
    .B(_1014_),
    .Y(_1015_));
 sg13g2_or2_1 _1989_ (.X(_1017_),
    .B(_1015_),
    .A(_0819_));
 sg13g2_xnor2_1 _1990_ (.Y(_1018_),
    .A(_0819_),
    .B(_1015_));
 sg13g2_nor2_2 _1991_ (.A(net77),
    .B(_0986_),
    .Y(_1019_));
 sg13g2_or2_1 _1992_ (.X(_1020_),
    .B(_0986_),
    .A(net76));
 sg13g2_xor2_1 _1993_ (.B(_1018_),
    .A(_1012_),
    .X(_1021_));
 sg13g2_a22oi_1 _1994_ (.Y(_1022_),
    .B1(_1019_),
    .B2(_1021_),
    .A2(_0992_),
    .A1(net77));
 sg13g2_o21ai_1 _1995_ (.B1(_1017_),
    .Y(_1023_),
    .A1(_1012_),
    .A2(_1018_));
 sg13g2_a21oi_2 _1996_ (.B1(net77),
    .Y(_1024_),
    .A2(_1023_),
    .A1(_1019_));
 sg13g2_nand2_1 _1997_ (.Y(_1025_),
    .A(net77),
    .B(_0991_));
 sg13g2_nand4_1 _1998_ (.B(_0679_),
    .C(_0683_),
    .A(_0641_),
    .Y(_1026_),
    .D(_1025_));
 sg13g2_inv_2 _1999_ (.Y(_1028_),
    .A(_1026_));
 sg13g2_nand2b_1 _2000_ (.Y(_1029_),
    .B(_0985_),
    .A_N(_0930_));
 sg13g2_nor2_2 _2001_ (.A(_1024_),
    .B(_1028_),
    .Y(_1030_));
 sg13g2_nand2b_2 _2002_ (.Y(_1031_),
    .B(_1026_),
    .A_N(_1024_));
 sg13g2_xor2_1 _2003_ (.B(_1011_),
    .A(_1010_),
    .X(_1032_));
 sg13g2_xnor2_1 _2004_ (.Y(_1033_),
    .A(_0810_),
    .B(_0988_));
 sg13g2_a22oi_1 _2005_ (.Y(_1034_),
    .B1(_1033_),
    .B2(net77),
    .A2(_1032_),
    .A1(_1019_));
 sg13g2_and2_1 _2006_ (.A(_1031_),
    .B(_1034_),
    .X(_1035_));
 sg13g2_nor2b_2 _2007_ (.A(net77),
    .B_N(_0986_),
    .Y(_1036_));
 sg13g2_nand2_2 _2008_ (.Y(_1037_),
    .A(_0609_),
    .B(_0683_));
 sg13g2_nor2_2 _2009_ (.A(_1036_),
    .B(_1037_),
    .Y(_1039_));
 sg13g2_nor2_1 _2010_ (.A(_1022_),
    .B(_1031_),
    .Y(_1040_));
 sg13g2_inv_1 _2011_ (.Y(_1041_),
    .A(_1040_));
 sg13g2_xnor2_1 _2012_ (.Y(_1042_),
    .A(_1022_),
    .B(_1030_));
 sg13g2_xnor2_1 _2013_ (.Y(_1043_),
    .A(_1030_),
    .B(_1034_));
 sg13g2_inv_1 _2014_ (.Y(_1044_),
    .A(net72));
 sg13g2_nand2_1 _2015_ (.Y(_1045_),
    .A(_0989_),
    .B(_1009_));
 sg13g2_a21o_1 _2016_ (.A2(_1045_),
    .A1(_1010_),
    .B1(_1020_),
    .X(_1046_));
 sg13g2_nand2_1 _2017_ (.Y(_1047_),
    .A(net77),
    .B(_0988_));
 sg13g2_nand2_1 _2018_ (.Y(_1048_),
    .A(_1046_),
    .B(_1047_));
 sg13g2_and2_1 _2019_ (.A(_1046_),
    .B(_1047_),
    .X(_1050_));
 sg13g2_nor4_2 _2020_ (.A(_1022_),
    .B(_1024_),
    .C(_1028_),
    .Y(_1051_),
    .D(_1034_));
 sg13g2_or4_1 _2021_ (.A(_1022_),
    .B(_1024_),
    .C(_1028_),
    .D(_1034_),
    .X(_1052_));
 sg13g2_nor2_1 _2022_ (.A(_1050_),
    .B(_1051_),
    .Y(_1053_));
 sg13g2_inv_1 _2023_ (.Y(_1054_),
    .A(_1053_));
 sg13g2_nor3_2 _2024_ (.A(_1031_),
    .B(_1050_),
    .C(_1051_),
    .Y(_1055_));
 sg13g2_nand3_1 _2025_ (.B(_1048_),
    .C(_1052_),
    .A(_1030_),
    .Y(_1056_));
 sg13g2_a21oi_2 _2026_ (.B1(_1030_),
    .Y(_1057_),
    .A2(_1052_),
    .A1(_1048_));
 sg13g2_o21ai_1 _2027_ (.B1(_1031_),
    .Y(_1058_),
    .A1(_1050_),
    .A2(_1051_));
 sg13g2_nor2_2 _2028_ (.A(_1055_),
    .B(_1057_),
    .Y(_1059_));
 sg13g2_nand2_2 _2029_ (.Y(_1061_),
    .A(_1056_),
    .B(_1058_));
 sg13g2_nand2_1 _2030_ (.Y(_1062_),
    .A(net76),
    .B(_0974_));
 sg13g2_nand2_1 _2031_ (.Y(_1063_),
    .A(_0955_),
    .B(net74));
 sg13g2_o21ai_1 _2032_ (.B1(_1063_),
    .Y(_1064_),
    .A1(_0959_),
    .A2(net75));
 sg13g2_nand2b_1 _2033_ (.Y(_1065_),
    .B(_1001_),
    .A_N(_1064_));
 sg13g2_nand2_1 _2034_ (.Y(_1066_),
    .A(_0977_),
    .B(net75));
 sg13g2_o21ai_1 _2035_ (.B1(_1066_),
    .Y(_1067_),
    .A1(_0982_),
    .A2(net75));
 sg13g2_nand2b_2 _2036_ (.Y(_1068_),
    .B(_1029_),
    .A_N(_1015_));
 sg13g2_mux2_1 _2037_ (.A0(_0965_),
    .A1(_0963_),
    .S(net75),
    .X(_1069_));
 sg13g2_nand2_1 _2038_ (.Y(_1070_),
    .A(_1000_),
    .B(_1069_));
 sg13g2_nor2_1 _2039_ (.A(_0922_),
    .B(net74),
    .Y(_1072_));
 sg13g2_a21oi_1 _2040_ (.A1(_0929_),
    .A2(net74),
    .Y(_1073_),
    .B1(_1072_));
 sg13g2_nand2_1 _2041_ (.Y(_1074_),
    .A(_1001_),
    .B(_1073_));
 sg13g2_nand3_1 _2042_ (.B(_1070_),
    .C(_1074_),
    .A(_1029_),
    .Y(_1075_));
 sg13g2_a22oi_1 _2043_ (.Y(_1076_),
    .B1(_1068_),
    .B2(_1075_),
    .A2(_1067_),
    .A1(_1065_));
 sg13g2_o21ai_1 _2044_ (.B1(_1062_),
    .Y(_1077_),
    .A1(_1020_),
    .A2(_1076_));
 sg13g2_nand2b_2 _2045_ (.Y(_1078_),
    .B(_1019_),
    .A_N(_1015_));
 sg13g2_nor2_1 _2046_ (.A(_0955_),
    .B(net75),
    .Y(_1079_));
 sg13g2_a21oi_1 _2047_ (.A1(_0982_),
    .A2(net75),
    .Y(_1080_),
    .B1(_1079_));
 sg13g2_nand2_1 _2048_ (.Y(_1081_),
    .A(_1000_),
    .B(_1080_));
 sg13g2_nor2_1 _2049_ (.A(_0963_),
    .B(net75),
    .Y(_1083_));
 sg13g2_a21oi_1 _2050_ (.A1(_0959_),
    .A2(net74),
    .Y(_1084_),
    .B1(_1083_));
 sg13g2_a21oi_1 _2051_ (.A1(_1001_),
    .A2(_1084_),
    .Y(_1085_),
    .B1(_1068_));
 sg13g2_a21oi_1 _2052_ (.A1(_1081_),
    .A2(_1085_),
    .Y(_1086_),
    .B1(_1078_));
 sg13g2_a21o_2 _2053_ (.A2(_0977_),
    .A1(net76),
    .B1(_1086_),
    .X(_1087_));
 sg13g2_nand3_1 _2054_ (.B(_1058_),
    .C(_1087_),
    .A(_1056_),
    .Y(_1088_));
 sg13g2_o21ai_1 _2055_ (.B1(_1077_),
    .Y(_1089_),
    .A1(_1055_),
    .A2(_1057_));
 sg13g2_a21o_1 _2056_ (.A2(_1089_),
    .A1(_1088_),
    .B1(net72),
    .X(_1090_));
 sg13g2_nand2_1 _2057_ (.Y(_1091_),
    .A(net76),
    .B(_0955_));
 sg13g2_nand2_1 _2058_ (.Y(_1092_),
    .A(_0965_),
    .B(net74));
 sg13g2_o21ai_1 _2059_ (.B1(_1092_),
    .Y(_0009_),
    .A1(_0929_),
    .A2(net74));
 sg13g2_mux2_1 _2060_ (.A0(_1084_),
    .A1(_0009_),
    .S(_1001_),
    .X(_0010_));
 sg13g2_nor2_1 _2061_ (.A(_1068_),
    .B(_0010_),
    .Y(_0011_));
 sg13g2_o21ai_1 _2062_ (.B1(_1091_),
    .Y(_0012_),
    .A1(_1078_),
    .A2(_0011_));
 sg13g2_nand2_1 _2063_ (.Y(_0013_),
    .A(net76),
    .B(_0981_));
 sg13g2_a21o_1 _2064_ (.A2(_1064_),
    .A1(_1000_),
    .B1(_1068_),
    .X(_0014_));
 sg13g2_a21oi_1 _2065_ (.A1(_1001_),
    .A2(_1069_),
    .Y(_0015_),
    .B1(_0014_));
 sg13g2_o21ai_1 _2066_ (.B1(_0013_),
    .Y(_0016_),
    .A1(_1078_),
    .A2(_0015_));
 sg13g2_inv_1 _2067_ (.Y(_0017_),
    .A(_0016_));
 sg13g2_mux2_1 _2068_ (.A0(_0012_),
    .A1(_0016_),
    .S(_1061_),
    .X(_0018_));
 sg13g2_mux4_1 _2069_ (.S0(_1059_),
    .A0(_1077_),
    .A1(_1087_),
    .A2(_0016_),
    .A3(_0012_),
    .S1(net72),
    .X(_0020_));
 sg13g2_nand2b_1 _2070_ (.Y(_0021_),
    .B(_1015_),
    .A_N(_0010_));
 sg13g2_nand2_1 _2071_ (.Y(_0022_),
    .A(_1001_),
    .B(_1080_));
 sg13g2_a21oi_1 _2072_ (.A1(_0971_),
    .A2(_0978_),
    .Y(_0023_),
    .B1(_0975_));
 sg13g2_nor2_1 _2073_ (.A(_1015_),
    .B(_0023_),
    .Y(_0024_));
 sg13g2_a21oi_1 _2074_ (.A1(_0022_),
    .A2(_0024_),
    .Y(_0025_),
    .B1(_1020_));
 sg13g2_a21oi_1 _2075_ (.A1(_0021_),
    .A2(_0025_),
    .Y(_0026_),
    .B1(_0970_));
 sg13g2_inv_1 _2076_ (.Y(_0027_),
    .A(_0026_));
 sg13g2_o21ai_1 _2077_ (.B1(_1056_),
    .Y(_0028_),
    .A1(_1057_),
    .A2(_0027_));
 sg13g2_a21oi_1 _2078_ (.A1(net73),
    .A2(_0028_),
    .Y(_0029_),
    .B1(_1035_));
 sg13g2_mux2_1 _2079_ (.A0(_0029_),
    .A1(_0020_),
    .S(_1042_),
    .X(_0031_));
 sg13g2_a21oi_1 _2080_ (.A1(_1056_),
    .A2(_1058_),
    .Y(_0032_),
    .B1(_1087_));
 sg13g2_a21oi_1 _2081_ (.A1(_1059_),
    .A2(_0017_),
    .Y(_0033_),
    .B1(_0032_));
 sg13g2_a21o_1 _2082_ (.A2(_0017_),
    .A1(_1059_),
    .B1(_0032_),
    .X(_0034_));
 sg13g2_nor2b_1 _2083_ (.A(_1078_),
    .B_N(_1075_),
    .Y(_0035_));
 sg13g2_a21o_1 _2084_ (.A2(_0958_),
    .A1(net76),
    .B1(_0035_),
    .X(_0036_));
 sg13g2_nand3_1 _2085_ (.B(_1058_),
    .C(_0036_),
    .A(_1056_),
    .Y(_0037_));
 sg13g2_o21ai_1 _2086_ (.B1(_0012_),
    .Y(_0038_),
    .A1(_1055_),
    .A2(_1057_));
 sg13g2_nand2_1 _2087_ (.Y(_0039_),
    .A(_0037_),
    .B(_0038_));
 sg13g2_and2_1 _2088_ (.A(_0037_),
    .B(_0038_),
    .X(_0040_));
 sg13g2_mux4_1 _2089_ (.S0(net72),
    .A0(_1087_),
    .A1(_0012_),
    .A2(_0016_),
    .A3(_0036_),
    .S1(_1059_),
    .X(_0042_));
 sg13g2_o21ai_1 _2090_ (.B1(_0026_),
    .Y(_0043_),
    .A1(_1055_),
    .A2(_1057_));
 sg13g2_mux2_1 _2091_ (.A0(_1077_),
    .A1(_0027_),
    .S(_1061_),
    .X(_0044_));
 sg13g2_o21ai_1 _2092_ (.B1(_0043_),
    .Y(_0045_),
    .A1(_1061_),
    .A2(_1077_));
 sg13g2_nor2_1 _2093_ (.A(net73),
    .B(_1053_),
    .Y(_0046_));
 sg13g2_a21oi_1 _2094_ (.A1(net73),
    .A2(_0045_),
    .Y(_0047_),
    .B1(_0046_));
 sg13g2_mux4_1 _2095_ (.S0(_1042_),
    .A0(_1053_),
    .A1(_0033_),
    .A2(_0044_),
    .A3(_0039_),
    .S1(net73),
    .X(_0048_));
 sg13g2_mux4_1 _2096_ (.S0(_1042_),
    .A0(_1054_),
    .A1(_0034_),
    .A2(_0045_),
    .A3(_0040_),
    .S1(net72),
    .X(_0049_));
 sg13g2_nand2_1 _2097_ (.Y(_0050_),
    .A(_0031_),
    .B(_0048_));
 sg13g2_nor2_1 _2098_ (.A(_0020_),
    .B(_0029_),
    .Y(_0051_));
 sg13g2_nor2_1 _2099_ (.A(net73),
    .B(_0028_),
    .Y(_0053_));
 sg13g2_a21oi_1 _2100_ (.A1(_1088_),
    .A2(_1089_),
    .Y(_0054_),
    .B1(_1044_));
 sg13g2_nor2_1 _2101_ (.A(_0053_),
    .B(_0054_),
    .Y(_0055_));
 sg13g2_mux4_1 _2102_ (.S0(net72),
    .A0(_1077_),
    .A1(_0016_),
    .A2(_0027_),
    .A3(_1087_),
    .S1(_1061_),
    .X(_0056_));
 sg13g2_nor4_1 _2103_ (.A(_0042_),
    .B(_0053_),
    .C(_0054_),
    .D(_0056_),
    .Y(_0057_));
 sg13g2_nor2_1 _2104_ (.A(_0995_),
    .B(net74),
    .Y(_0058_));
 sg13g2_a21oi_1 _2105_ (.A1(_0924_),
    .A2(net74),
    .Y(_0059_),
    .B1(_0058_));
 sg13g2_nand3_1 _2106_ (.B(_1019_),
    .C(_1073_),
    .A(_1000_),
    .Y(_0060_));
 sg13g2_a22oi_1 _2107_ (.Y(_0061_),
    .B1(net72),
    .B2(_0059_),
    .A2(_0965_),
    .A1(net76));
 sg13g2_a21oi_1 _2108_ (.A1(_0060_),
    .A2(_0061_),
    .Y(_0062_),
    .B1(_1061_));
 sg13g2_o21ai_1 _2109_ (.B1(_0036_),
    .Y(_0064_),
    .A1(_1055_),
    .A2(_1057_));
 sg13g2_a21oi_1 _2110_ (.A1(_1000_),
    .A2(_0009_),
    .Y(_0065_),
    .B1(_1068_));
 sg13g2_nor2_1 _2111_ (.A(_1078_),
    .B(_0065_),
    .Y(_0066_));
 sg13g2_a21oi_1 _2112_ (.A1(net76),
    .A2(_0963_),
    .Y(_0067_),
    .B1(_0066_));
 sg13g2_nand3_1 _2113_ (.B(_0064_),
    .C(_0067_),
    .A(_1042_),
    .Y(_0068_));
 sg13g2_a21oi_1 _2114_ (.A1(_0037_),
    .A2(_0038_),
    .Y(_0069_),
    .B1(net72));
 sg13g2_nor4_1 _2115_ (.A(_0018_),
    .B(_0062_),
    .C(_0068_),
    .D(_0069_),
    .Y(_0070_));
 sg13g2_a221oi_1 _2116_ (.B2(_1090_),
    .C1(_0049_),
    .B1(_0070_),
    .A1(_0051_),
    .Y(_0071_),
    .A2(_0057_));
 sg13g2_o21ai_1 _2117_ (.B1(_0050_),
    .Y(_0072_),
    .A1(_0031_),
    .A2(_0071_));
 sg13g2_nor3_1 _2118_ (.A(_1036_),
    .B(_1037_),
    .C(_0072_),
    .Y(_0073_));
 sg13g2_nor2_2 _2119_ (.A(net38),
    .B(_0683_),
    .Y(_0075_));
 sg13g2_nor2b_1 _2120_ (.A(_0611_),
    .B_N(_0075_),
    .Y(_0076_));
 sg13g2_nor3_1 _2121_ (.A(net95),
    .B(_0073_),
    .C(_0076_),
    .Y(_0077_));
 sg13g2_a21oi_1 _2122_ (.A1(_0433_),
    .A2(net95),
    .Y(_0000_),
    .B1(_0077_));
 sg13g2_nor2_1 _2123_ (.A(_0591_),
    .B(net84),
    .Y(_0078_));
 sg13g2_a21oi_2 _2124_ (.B1(_0078_),
    .Y(_0079_),
    .A2(net84),
    .A1(_0400_));
 sg13g2_inv_2 _2125_ (.Y(_0080_),
    .A(_0079_));
 sg13g2_a21oi_1 _2126_ (.A1(net73),
    .A2(_1054_),
    .Y(_0081_),
    .B1(_1035_));
 sg13g2_mux2_1 _2127_ (.A0(_0081_),
    .A1(_0056_),
    .S(_1042_),
    .X(_0082_));
 sg13g2_nand3_1 _2128_ (.B(_0048_),
    .C(_0082_),
    .A(_0031_),
    .Y(_0083_));
 sg13g2_xor2_1 _2129_ (.B(_0082_),
    .A(_0050_),
    .X(_0085_));
 sg13g2_o21ai_1 _2130_ (.B1(_0085_),
    .Y(_0086_),
    .A1(_0072_),
    .A2(_0080_));
 sg13g2_or3_1 _2131_ (.A(_0072_),
    .B(_0080_),
    .C(_0085_),
    .X(_0087_));
 sg13g2_nand3_1 _2132_ (.B(_0086_),
    .C(_0087_),
    .A(_1039_),
    .Y(_0088_));
 sg13g2_nand4_1 _2133_ (.B(_0612_),
    .C(_0613_),
    .A(net99),
    .Y(_0089_),
    .D(_0075_));
 sg13g2_a21oi_1 _2134_ (.A1(_0088_),
    .A2(_0089_),
    .Y(_0090_),
    .B1(net95));
 sg13g2_a21o_1 _2135_ (.A2(_0631_),
    .A1(net40),
    .B1(_0090_),
    .X(_0001_));
 sg13g2_a21oi_1 _2136_ (.A1(_0072_),
    .A2(_0085_),
    .Y(_0091_),
    .B1(_0080_));
 sg13g2_a21oi_1 _2137_ (.A1(_1041_),
    .A2(_0055_),
    .Y(_0092_),
    .B1(_1036_));
 sg13g2_a21o_2 _2138_ (.A2(_0055_),
    .A1(_1041_),
    .B1(_1036_),
    .X(_0093_));
 sg13g2_nand2b_1 _2139_ (.Y(_0095_),
    .B(_0092_),
    .A_N(_0083_));
 sg13g2_xnor2_1 _2140_ (.Y(_0096_),
    .A(_0083_),
    .B(_0092_));
 sg13g2_xnor2_1 _2141_ (.Y(_0097_),
    .A(_0083_),
    .B(_0093_));
 sg13g2_o21ai_1 _2142_ (.B1(_1039_),
    .Y(_0098_),
    .A1(_0091_),
    .A2(_0096_));
 sg13g2_a21o_1 _2143_ (.A2(_0096_),
    .A1(_0091_),
    .B1(_0098_),
    .X(_0099_));
 sg13g2_nand3_1 _2144_ (.B(_0607_),
    .C(_0075_),
    .A(_0587_),
    .Y(_0100_));
 sg13g2_nor2b_1 _2145_ (.A(net96),
    .B_N(_0100_),
    .Y(_0101_));
 sg13g2_a22oi_1 _2146_ (.Y(_0002_),
    .B1(_0099_),
    .B2(_0101_),
    .A2(net96),
    .A1(_0422_));
 sg13g2_a221oi_1 _2147_ (.B2(_0047_),
    .C1(_1040_),
    .B1(_1042_),
    .A1(_1022_),
    .Y(_0102_),
    .A2(_1035_));
 sg13g2_nor3_1 _2148_ (.A(_0083_),
    .B(_0093_),
    .C(_0102_),
    .Y(_0103_));
 sg13g2_or2_1 _2149_ (.X(_0105_),
    .B(_0102_),
    .A(_1036_));
 sg13g2_a21oi_1 _2150_ (.A1(_0095_),
    .A2(_0105_),
    .Y(_0106_),
    .B1(_0103_));
 sg13g2_nand3_1 _2151_ (.B(_0085_),
    .C(_0097_),
    .A(_0072_),
    .Y(_0107_));
 sg13g2_nand2_1 _2152_ (.Y(_0108_),
    .A(_0079_),
    .B(_0107_));
 sg13g2_xnor2_1 _2153_ (.Y(_0109_),
    .A(_0106_),
    .B(_0108_));
 sg13g2_a221oi_1 _2154_ (.B2(_1039_),
    .C1(net95),
    .B1(_0109_),
    .A1(_0599_),
    .Y(_0110_),
    .A2(_0075_));
 sg13g2_a21oi_1 _2155_ (.A1(_0411_),
    .A2(net95),
    .Y(_0003_),
    .B1(_0110_));
 sg13g2_a21o_1 _2156_ (.A2(_0029_),
    .A1(_1042_),
    .B1(_1040_),
    .X(_0111_));
 sg13g2_inv_1 _2157_ (.Y(_0112_),
    .A(_0111_));
 sg13g2_nor4_1 _2158_ (.A(_0083_),
    .B(_0093_),
    .C(_0102_),
    .D(_0112_),
    .Y(_0113_));
 sg13g2_xnor2_1 _2159_ (.Y(_0115_),
    .A(_0103_),
    .B(_0112_));
 sg13g2_o21ai_1 _2160_ (.B1(_0079_),
    .Y(_0116_),
    .A1(_0106_),
    .A2(_0107_));
 sg13g2_nand2b_1 _2161_ (.Y(_0117_),
    .B(_0115_),
    .A_N(_0116_));
 sg13g2_nand2b_1 _2162_ (.Y(_0118_),
    .B(_0116_),
    .A_N(_0115_));
 sg13g2_nand3_1 _2163_ (.B(_0117_),
    .C(_0118_),
    .A(_1039_),
    .Y(_0119_));
 sg13g2_a21oi_1 _2164_ (.A1(_0596_),
    .A2(_0075_),
    .Y(_0120_),
    .B1(net96));
 sg13g2_a22oi_1 _2165_ (.Y(_0004_),
    .B1(_0119_),
    .B2(_0120_),
    .A2(net95),
    .A1(_0455_));
 sg13g2_a21oi_1 _2166_ (.A1(_1042_),
    .A2(_0081_),
    .Y(_0121_),
    .B1(_1040_));
 sg13g2_nor2b_1 _2167_ (.A(_0113_),
    .B_N(_0121_),
    .Y(_0122_));
 sg13g2_nand2b_1 _2168_ (.Y(_0123_),
    .B(_0121_),
    .A_N(_0113_));
 sg13g2_nand2_1 _2169_ (.Y(_0125_),
    .A(_0079_),
    .B(_0115_));
 sg13g2_a21o_1 _2170_ (.A2(_0125_),
    .A1(_0116_),
    .B1(_0122_),
    .X(_0126_));
 sg13g2_nand3_1 _2171_ (.B(_0122_),
    .C(_0125_),
    .A(_0116_),
    .Y(_0127_));
 sg13g2_nand3_1 _2172_ (.B(_0126_),
    .C(_0127_),
    .A(_1039_),
    .Y(_0128_));
 sg13g2_a21oi_1 _2173_ (.A1(_0594_),
    .A2(_0075_),
    .Y(_0129_),
    .B1(net96));
 sg13g2_a22oi_1 _2174_ (.Y(_0005_),
    .B1(_0128_),
    .B2(_0129_),
    .A2(net95),
    .A1(_0444_));
 sg13g2_or4_1 _2175_ (.A(_0106_),
    .B(_0107_),
    .C(_0115_),
    .D(_0123_),
    .X(_0130_));
 sg13g2_a21oi_1 _2176_ (.A1(_0079_),
    .A2(_0130_),
    .Y(_0131_),
    .B1(_1030_));
 sg13g2_nand3_1 _2177_ (.B(_0079_),
    .C(_0130_),
    .A(_1030_),
    .Y(_0132_));
 sg13g2_nand3b_1 _2178_ (.B(_0132_),
    .C(_1039_),
    .Y(_0133_),
    .A_N(_0131_));
 sg13g2_a21oi_1 _2179_ (.A1(_0590_),
    .A2(_0075_),
    .Y(_0135_),
    .B1(net96));
 sg13g2_a22oi_1 _2180_ (.Y(_0006_),
    .B1(_0133_),
    .B2(_0135_),
    .A2(net95),
    .A1(_0466_));
 sg13g2_nand2_1 _2181_ (.Y(_0136_),
    .A(net38),
    .B(net96));
 sg13g2_nor2_1 _2182_ (.A(_1036_),
    .B(_0080_),
    .Y(_0137_));
 sg13g2_a21oi_1 _2183_ (.A1(_0592_),
    .A2(_0075_),
    .Y(_0138_),
    .B1(net96));
 sg13g2_o21ai_1 _2184_ (.B1(_0138_),
    .Y(_0139_),
    .A1(_1037_),
    .A2(_0137_));
 sg13g2_nand2_1 _2185_ (.Y(_0007_),
    .A(_0136_),
    .B(_0139_));
 sg13g2_dfrbpq_2 _2186_ (.RESET_B(net2),
    .D(_0000_),
    .Q(uo_out[0]),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _2187_ (.RESET_B(net2),
    .D(_0001_),
    .Q(uo_out[1]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _2188_ (.RESET_B(net2),
    .D(_0002_),
    .Q(uo_out[2]),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _2189_ (.RESET_B(net2),
    .D(_0003_),
    .Q(uo_out[3]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _2190_ (.RESET_B(net2),
    .D(net37),
    .Q(uo_out[4]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _2191_ (.RESET_B(net2),
    .D(_0005_),
    .Q(uo_out[5]),
    .CLK(clknet_1_1__leaf_clk));
 sg13g2_dfrbpq_2 _2192_ (.RESET_B(net2),
    .D(_0006_),
    .Q(uo_out[6]),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_dfrbpq_2 _2193_ (.RESET_B(net2),
    .D(_0007_),
    .Q(\u_mac.u_adder.sign_b ),
    .CLK(clknet_1_0__leaf_clk));
 sg13g2_tielo tt_um_posit_mac_stream_19 (.L_LO(net19));
 sg13g2_tielo tt_um_posit_mac_stream_20 (.L_LO(net20));
 sg13g2_tielo tt_um_posit_mac_stream_21 (.L_LO(net21));
 sg13g2_tielo tt_um_posit_mac_stream_22 (.L_LO(net22));
 sg13g2_tielo tt_um_posit_mac_stream_23 (.L_LO(net23));
 sg13g2_tielo tt_um_posit_mac_stream_24 (.L_LO(net24));
 sg13g2_tielo tt_um_posit_mac_stream_25 (.L_LO(net25));
 sg13g2_tielo tt_um_posit_mac_stream_26 (.L_LO(net26));
 sg13g2_tielo tt_um_posit_mac_stream_27 (.L_LO(net27));
 sg13g2_tielo tt_um_posit_mac_stream_28 (.L_LO(net28));
 sg13g2_tielo tt_um_posit_mac_stream_29 (.L_LO(net29));
 sg13g2_tielo tt_um_posit_mac_stream_30 (.L_LO(net30));
 sg13g2_tielo tt_um_posit_mac_stream_31 (.L_LO(net31));
 sg13g2_tielo tt_um_posit_mac_stream_32 (.L_LO(net32));
 sg13g2_tielo tt_um_posit_mac_stream_33 (.L_LO(net33));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2210_ (.A(\u_mac.u_adder.sign_b ),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout72 (.A(_1043_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1043_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(net75),
    .X(net74));
 sg13g2_buf_8 fanout75 (.A(_1009_),
    .X(net75));
 sg13g2_buf_8 fanout76 (.A(_0953_),
    .X(net76));
 sg13g2_buf_8 fanout77 (.A(_0953_),
    .X(net77));
 sg13g2_buf_8 fanout78 (.A(_0822_),
    .X(net78));
 sg13g2_buf_8 fanout79 (.A(_0817_),
    .X(net79));
 sg13g2_buf_1 fanout80 (.A(_0817_),
    .X(net80));
 sg13g2_buf_8 fanout81 (.A(net83),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(net83),
    .X(net82));
 sg13g2_buf_8 fanout83 (.A(_0793_),
    .X(net83));
 sg13g2_buf_8 fanout84 (.A(_0793_),
    .X(net84));
 sg13g2_buf_8 fanout85 (.A(_0783_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(net87),
    .X(net86));
 sg13g2_buf_1 fanout87 (.A(_0625_),
    .X(net87));
 sg13g2_buf_8 fanout88 (.A(_0603_),
    .X(net88));
 sg13g2_buf_8 fanout89 (.A(_0468_),
    .X(net89));
 sg13g2_buf_8 fanout90 (.A(net92),
    .X(net90));
 sg13g2_buf_1 fanout91 (.A(net92),
    .X(net91));
 sg13g2_buf_8 fanout92 (.A(_0410_),
    .X(net92));
 sg13g2_buf_8 fanout93 (.A(_0669_),
    .X(net93));
 sg13g2_buf_1 fanout94 (.A(_0669_),
    .X(net94));
 sg13g2_buf_8 fanout95 (.A(net96),
    .X(net95));
 sg13g2_buf_8 fanout96 (.A(_0631_),
    .X(net96));
 sg13g2_buf_8 fanout97 (.A(net98),
    .X(net97));
 sg13g2_buf_8 fanout98 (.A(_0598_),
    .X(net98));
 sg13g2_buf_8 fanout99 (.A(_0587_),
    .X(net99));
 sg13g2_buf_8 fanout100 (.A(net101),
    .X(net100));
 sg13g2_buf_8 fanout101 (.A(_0653_),
    .X(net101));
 sg13g2_buf_8 fanout102 (.A(net103),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103));
 sg13g2_buf_1 fanout104 (.A(uio_in[7]),
    .X(net104));
 sg13g2_buf_8 fanout105 (.A(net10),
    .X(net105));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_2 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[1]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[2]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[3]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[4]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[5]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[6]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(ui_in[7]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[0]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[1]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[2]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[3]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[4]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[5]),
    .X(net16));
 sg13g2_buf_2 input17 (.A(uio_in[6]),
    .X(net17));
 sg13g2_tielo tt_um_posit_mac_stream_18 (.L_LO(net18));
 sg13g2_buf_8 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sg13g2_buf_8 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(uo_out[5]),
    .X(net34));
 sg13g2_dlygate4sd3_1 hold2 (.A(uo_out[3]),
    .X(net35));
 sg13g2_dlygate4sd3_1 hold3 (.A(uo_out[4]),
    .X(net36));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0004_),
    .X(net37));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u_mac.u_adder.sign_b ),
    .X(net38));
 sg13g2_dlygate4sd3_1 hold6 (.A(uo_out[6]),
    .X(net39));
 sg13g2_dlygate4sd3_1 hold7 (.A(uo_out[1]),
    .X(net40));
 sg13g2_dlygate4sd3_1 hold8 (.A(uo_out[2]),
    .X(net41));
 sg13g2_dlygate4sd3_1 hold9 (.A(uo_out[0]),
    .X(net42));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_406 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_fill_2 FILLER_7_406 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_fill_2 FILLER_9_91 ();
 sg13g2_fill_1 FILLER_9_93 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_70 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_125 ();
 sg13g2_fill_1 FILLER_10_136 ();
 sg13g2_decap_8 FILLER_10_142 ();
 sg13g2_decap_8 FILLER_10_149 ();
 sg13g2_decap_8 FILLER_10_156 ();
 sg13g2_decap_8 FILLER_10_163 ();
 sg13g2_decap_8 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_177 ();
 sg13g2_decap_8 FILLER_10_184 ();
 sg13g2_decap_8 FILLER_10_191 ();
 sg13g2_decap_8 FILLER_10_198 ();
 sg13g2_decap_8 FILLER_10_205 ();
 sg13g2_decap_8 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_decap_8 FILLER_10_226 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_decap_8 FILLER_10_240 ();
 sg13g2_decap_8 FILLER_10_247 ();
 sg13g2_decap_8 FILLER_10_254 ();
 sg13g2_decap_8 FILLER_10_261 ();
 sg13g2_decap_8 FILLER_10_268 ();
 sg13g2_decap_8 FILLER_10_275 ();
 sg13g2_decap_8 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_289 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_8 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_310 ();
 sg13g2_decap_8 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_324 ();
 sg13g2_decap_8 FILLER_10_331 ();
 sg13g2_decap_8 FILLER_10_338 ();
 sg13g2_decap_8 FILLER_10_345 ();
 sg13g2_decap_8 FILLER_10_352 ();
 sg13g2_decap_8 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_366 ();
 sg13g2_decap_8 FILLER_10_373 ();
 sg13g2_decap_8 FILLER_10_380 ();
 sg13g2_decap_8 FILLER_10_387 ();
 sg13g2_decap_8 FILLER_10_394 ();
 sg13g2_decap_8 FILLER_10_401 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_37 ();
 sg13g2_decap_8 FILLER_11_41 ();
 sg13g2_decap_4 FILLER_11_48 ();
 sg13g2_fill_1 FILLER_11_65 ();
 sg13g2_decap_8 FILLER_11_75 ();
 sg13g2_decap_8 FILLER_11_82 ();
 sg13g2_fill_2 FILLER_11_89 ();
 sg13g2_fill_1 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_97 ();
 sg13g2_decap_4 FILLER_11_104 ();
 sg13g2_fill_1 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_fill_2 FILLER_11_144 ();
 sg13g2_fill_1 FILLER_11_146 ();
 sg13g2_decap_4 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_170 ();
 sg13g2_decap_8 FILLER_11_177 ();
 sg13g2_decap_4 FILLER_11_184 ();
 sg13g2_fill_1 FILLER_11_188 ();
 sg13g2_decap_8 FILLER_11_195 ();
 sg13g2_decap_8 FILLER_11_202 ();
 sg13g2_decap_8 FILLER_11_209 ();
 sg13g2_decap_8 FILLER_11_216 ();
 sg13g2_decap_8 FILLER_11_223 ();
 sg13g2_decap_4 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_4 FILLER_11_273 ();
 sg13g2_fill_1 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_288 ();
 sg13g2_decap_8 FILLER_11_295 ();
 sg13g2_decap_8 FILLER_11_302 ();
 sg13g2_decap_8 FILLER_11_309 ();
 sg13g2_decap_8 FILLER_11_316 ();
 sg13g2_decap_8 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_330 ();
 sg13g2_decap_8 FILLER_11_337 ();
 sg13g2_decap_8 FILLER_11_344 ();
 sg13g2_decap_8 FILLER_11_351 ();
 sg13g2_decap_8 FILLER_11_358 ();
 sg13g2_decap_8 FILLER_11_365 ();
 sg13g2_decap_8 FILLER_11_372 ();
 sg13g2_decap_8 FILLER_11_379 ();
 sg13g2_decap_8 FILLER_11_386 ();
 sg13g2_decap_8 FILLER_11_393 ();
 sg13g2_decap_8 FILLER_11_400 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_62 ();
 sg13g2_decap_4 FILLER_12_108 ();
 sg13g2_decap_4 FILLER_12_127 ();
 sg13g2_fill_2 FILLER_12_131 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_fill_2 FILLER_12_166 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_fill_1 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_265 ();
 sg13g2_decap_4 FILLER_12_272 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_decap_4 FILLER_12_300 ();
 sg13g2_fill_2 FILLER_12_304 ();
 sg13g2_fill_2 FILLER_12_320 ();
 sg13g2_fill_1 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_fill_1 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_360 ();
 sg13g2_decap_8 FILLER_12_367 ();
 sg13g2_decap_8 FILLER_12_374 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_2 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_40 ();
 sg13g2_decap_8 FILLER_13_47 ();
 sg13g2_decap_8 FILLER_13_71 ();
 sg13g2_decap_4 FILLER_13_78 ();
 sg13g2_decap_4 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_91 ();
 sg13g2_decap_4 FILLER_13_97 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_decap_4 FILLER_13_123 ();
 sg13g2_fill_1 FILLER_13_127 ();
 sg13g2_decap_4 FILLER_13_148 ();
 sg13g2_fill_2 FILLER_13_152 ();
 sg13g2_fill_2 FILLER_13_159 ();
 sg13g2_decap_8 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_190 ();
 sg13g2_fill_1 FILLER_13_192 ();
 sg13g2_decap_8 FILLER_13_213 ();
 sg13g2_decap_8 FILLER_13_220 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_233 ();
 sg13g2_decap_8 FILLER_13_243 ();
 sg13g2_decap_4 FILLER_13_250 ();
 sg13g2_decap_8 FILLER_13_272 ();
 sg13g2_fill_1 FILLER_13_279 ();
 sg13g2_decap_4 FILLER_13_293 ();
 sg13g2_fill_1 FILLER_13_297 ();
 sg13g2_decap_4 FILLER_13_340 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_365 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_8 FILLER_13_386 ();
 sg13g2_decap_8 FILLER_13_393 ();
 sg13g2_decap_8 FILLER_13_400 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_fill_2 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_23 ();
 sg13g2_fill_2 FILLER_14_43 ();
 sg13g2_fill_1 FILLER_14_45 ();
 sg13g2_decap_8 FILLER_14_94 ();
 sg13g2_fill_2 FILLER_14_101 ();
 sg13g2_decap_8 FILLER_14_113 ();
 sg13g2_decap_8 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_127 ();
 sg13g2_decap_4 FILLER_14_134 ();
 sg13g2_fill_2 FILLER_14_138 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_4 FILLER_14_151 ();
 sg13g2_fill_2 FILLER_14_171 ();
 sg13g2_decap_4 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_213 ();
 sg13g2_decap_4 FILLER_14_220 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_decap_4 FILLER_14_239 ();
 sg13g2_fill_1 FILLER_14_248 ();
 sg13g2_decap_8 FILLER_14_255 ();
 sg13g2_decap_4 FILLER_14_262 ();
 sg13g2_fill_2 FILLER_14_266 ();
 sg13g2_fill_2 FILLER_14_277 ();
 sg13g2_fill_1 FILLER_14_279 ();
 sg13g2_decap_4 FILLER_14_301 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_2 FILLER_14_312 ();
 sg13g2_fill_1 FILLER_14_314 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_fill_2 FILLER_14_327 ();
 sg13g2_fill_1 FILLER_14_329 ();
 sg13g2_fill_2 FILLER_14_335 ();
 sg13g2_decap_8 FILLER_14_342 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_decap_4 FILLER_14_360 ();
 sg13g2_decap_4 FILLER_14_368 ();
 sg13g2_fill_1 FILLER_14_372 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_19 ();
 sg13g2_decap_4 FILLER_15_26 ();
 sg13g2_fill_1 FILLER_15_30 ();
 sg13g2_decap_8 FILLER_15_43 ();
 sg13g2_decap_8 FILLER_15_50 ();
 sg13g2_fill_1 FILLER_15_57 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_101 ();
 sg13g2_fill_1 FILLER_15_108 ();
 sg13g2_decap_4 FILLER_15_115 ();
 sg13g2_decap_4 FILLER_15_143 ();
 sg13g2_fill_2 FILLER_15_147 ();
 sg13g2_fill_2 FILLER_15_157 ();
 sg13g2_fill_1 FILLER_15_159 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_fill_1 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_190 ();
 sg13g2_decap_4 FILLER_15_197 ();
 sg13g2_fill_2 FILLER_15_201 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_224 ();
 sg13g2_decap_8 FILLER_15_231 ();
 sg13g2_fill_1 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_255 ();
 sg13g2_decap_8 FILLER_15_264 ();
 sg13g2_decap_8 FILLER_15_271 ();
 sg13g2_fill_1 FILLER_15_278 ();
 sg13g2_decap_8 FILLER_15_289 ();
 sg13g2_decap_8 FILLER_15_296 ();
 sg13g2_decap_8 FILLER_15_303 ();
 sg13g2_fill_1 FILLER_15_310 ();
 sg13g2_fill_2 FILLER_15_324 ();
 sg13g2_fill_1 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_353 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_27 ();
 sg13g2_decap_8 FILLER_16_46 ();
 sg13g2_decap_4 FILLER_16_53 ();
 sg13g2_fill_1 FILLER_16_57 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_fill_1 FILLER_16_77 ();
 sg13g2_fill_2 FILLER_16_88 ();
 sg13g2_fill_1 FILLER_16_90 ();
 sg13g2_decap_8 FILLER_16_99 ();
 sg13g2_decap_8 FILLER_16_106 ();
 sg13g2_fill_2 FILLER_16_113 ();
 sg13g2_decap_4 FILLER_16_136 ();
 sg13g2_fill_1 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_157 ();
 sg13g2_decap_4 FILLER_16_164 ();
 sg13g2_fill_2 FILLER_16_178 ();
 sg13g2_fill_2 FILLER_16_187 ();
 sg13g2_fill_1 FILLER_16_189 ();
 sg13g2_fill_2 FILLER_16_195 ();
 sg13g2_fill_2 FILLER_16_212 ();
 sg13g2_decap_4 FILLER_16_228 ();
 sg13g2_fill_1 FILLER_16_232 ();
 sg13g2_decap_8 FILLER_16_246 ();
 sg13g2_decap_8 FILLER_16_253 ();
 sg13g2_decap_4 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_280 ();
 sg13g2_fill_1 FILLER_16_282 ();
 sg13g2_decap_4 FILLER_16_288 ();
 sg13g2_fill_2 FILLER_16_292 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_fill_1 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_4 FILLER_16_337 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_fill_2 FILLER_16_379 ();
 sg13g2_fill_1 FILLER_16_381 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_4 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_7 ();
 sg13g2_decap_4 FILLER_17_17 ();
 sg13g2_fill_1 FILLER_17_21 ();
 sg13g2_decap_4 FILLER_17_45 ();
 sg13g2_fill_2 FILLER_17_58 ();
 sg13g2_fill_1 FILLER_17_60 ();
 sg13g2_fill_2 FILLER_17_71 ();
 sg13g2_fill_1 FILLER_17_73 ();
 sg13g2_fill_2 FILLER_17_85 ();
 sg13g2_fill_1 FILLER_17_87 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_fill_1 FILLER_17_112 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_2 FILLER_17_127 ();
 sg13g2_decap_8 FILLER_17_139 ();
 sg13g2_fill_2 FILLER_17_146 ();
 sg13g2_decap_4 FILLER_17_154 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_fill_2 FILLER_17_171 ();
 sg13g2_decap_8 FILLER_17_176 ();
 sg13g2_decap_4 FILLER_17_183 ();
 sg13g2_fill_2 FILLER_17_187 ();
 sg13g2_decap_8 FILLER_17_194 ();
 sg13g2_fill_1 FILLER_17_201 ();
 sg13g2_decap_4 FILLER_17_209 ();
 sg13g2_fill_2 FILLER_17_213 ();
 sg13g2_decap_4 FILLER_17_252 ();
 sg13g2_fill_2 FILLER_17_256 ();
 sg13g2_decap_4 FILLER_17_280 ();
 sg13g2_fill_2 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_fill_1 FILLER_17_313 ();
 sg13g2_decap_8 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_325 ();
 sg13g2_fill_2 FILLER_17_331 ();
 sg13g2_fill_2 FILLER_17_349 ();
 sg13g2_fill_2 FILLER_17_380 ();
 sg13g2_fill_1 FILLER_17_382 ();
 sg13g2_fill_2 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_4 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_4 FILLER_18_25 ();
 sg13g2_fill_2 FILLER_18_29 ();
 sg13g2_decap_8 FILLER_18_40 ();
 sg13g2_decap_4 FILLER_18_47 ();
 sg13g2_fill_1 FILLER_18_51 ();
 sg13g2_fill_1 FILLER_18_61 ();
 sg13g2_decap_4 FILLER_18_67 ();
 sg13g2_fill_1 FILLER_18_71 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_fill_2 FILLER_18_88 ();
 sg13g2_fill_1 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_139 ();
 sg13g2_fill_1 FILLER_18_141 ();
 sg13g2_fill_2 FILLER_18_156 ();
 sg13g2_decap_4 FILLER_18_175 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_2 FILLER_18_197 ();
 sg13g2_fill_1 FILLER_18_199 ();
 sg13g2_fill_1 FILLER_18_212 ();
 sg13g2_decap_8 FILLER_18_223 ();
 sg13g2_fill_1 FILLER_18_230 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_fill_1 FILLER_18_282 ();
 sg13g2_decap_4 FILLER_18_299 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_decap_4 FILLER_18_315 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_fill_2 FILLER_18_351 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_4 FILLER_18_369 ();
 sg13g2_fill_1 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_fill_1 FILLER_18_388 ();
 sg13g2_fill_2 FILLER_18_407 ();
 sg13g2_decap_4 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_25 ();
 sg13g2_fill_1 FILLER_19_27 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_fill_2 FILLER_19_52 ();
 sg13g2_fill_1 FILLER_19_54 ();
 sg13g2_decap_4 FILLER_19_60 ();
 sg13g2_decap_4 FILLER_19_87 ();
 sg13g2_decap_4 FILLER_19_99 ();
 sg13g2_fill_2 FILLER_19_126 ();
 sg13g2_decap_4 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_138 ();
 sg13g2_decap_8 FILLER_19_143 ();
 sg13g2_decap_4 FILLER_19_150 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_decap_4 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_185 ();
 sg13g2_decap_8 FILLER_19_192 ();
 sg13g2_decap_8 FILLER_19_199 ();
 sg13g2_decap_4 FILLER_19_210 ();
 sg13g2_fill_1 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_225 ();
 sg13g2_fill_2 FILLER_19_230 ();
 sg13g2_decap_4 FILLER_19_249 ();
 sg13g2_decap_4 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_fill_2 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_fill_1 FILLER_19_335 ();
 sg13g2_decap_4 FILLER_19_349 ();
 sg13g2_fill_2 FILLER_19_358 ();
 sg13g2_fill_1 FILLER_19_360 ();
 sg13g2_decap_8 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_400 ();
 sg13g2_fill_2 FILLER_19_407 ();
 sg13g2_decap_4 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_17 ();
 sg13g2_decap_4 FILLER_20_24 ();
 sg13g2_decap_8 FILLER_20_58 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_fill_2 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_79 ();
 sg13g2_decap_8 FILLER_20_84 ();
 sg13g2_decap_8 FILLER_20_91 ();
 sg13g2_decap_8 FILLER_20_98 ();
 sg13g2_fill_2 FILLER_20_105 ();
 sg13g2_decap_8 FILLER_20_115 ();
 sg13g2_decap_4 FILLER_20_122 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_1 FILLER_20_138 ();
 sg13g2_fill_2 FILLER_20_144 ();
 sg13g2_fill_1 FILLER_20_146 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_4 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_186 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_decap_8 FILLER_20_208 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_decap_8 FILLER_20_239 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_decap_4 FILLER_20_278 ();
 sg13g2_fill_2 FILLER_20_282 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_decap_4 FILLER_20_299 ();
 sg13g2_fill_1 FILLER_20_303 ();
 sg13g2_fill_2 FILLER_20_309 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_decap_8 FILLER_20_330 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_4 FILLER_20_389 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_15 ();
 sg13g2_fill_1 FILLER_21_22 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_decap_4 FILLER_21_39 ();
 sg13g2_fill_2 FILLER_21_43 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_fill_2 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_87 ();
 sg13g2_fill_2 FILLER_21_102 ();
 sg13g2_decap_4 FILLER_21_116 ();
 sg13g2_fill_2 FILLER_21_120 ();
 sg13g2_decap_8 FILLER_21_127 ();
 sg13g2_decap_4 FILLER_21_134 ();
 sg13g2_decap_8 FILLER_21_142 ();
 sg13g2_fill_2 FILLER_21_149 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_fill_2 FILLER_21_169 ();
 sg13g2_decap_8 FILLER_21_176 ();
 sg13g2_fill_2 FILLER_21_188 ();
 sg13g2_fill_1 FILLER_21_190 ();
 sg13g2_decap_4 FILLER_21_205 ();
 sg13g2_fill_1 FILLER_21_230 ();
 sg13g2_decap_4 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_fill_2 FILLER_21_274 ();
 sg13g2_fill_1 FILLER_21_281 ();
 sg13g2_fill_1 FILLER_21_295 ();
 sg13g2_decap_8 FILLER_21_303 ();
 sg13g2_fill_2 FILLER_21_310 ();
 sg13g2_fill_1 FILLER_21_312 ();
 sg13g2_decap_4 FILLER_21_321 ();
 sg13g2_decap_4 FILLER_21_333 ();
 sg13g2_fill_2 FILLER_21_337 ();
 sg13g2_fill_1 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_360 ();
 sg13g2_fill_2 FILLER_21_367 ();
 sg13g2_decap_4 FILLER_21_387 ();
 sg13g2_fill_2 FILLER_21_391 ();
 sg13g2_decap_4 FILLER_21_403 ();
 sg13g2_fill_2 FILLER_21_407 ();
 sg13g2_decap_4 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_20 ();
 sg13g2_decap_4 FILLER_22_27 ();
 sg13g2_fill_2 FILLER_22_44 ();
 sg13g2_fill_1 FILLER_22_46 ();
 sg13g2_fill_1 FILLER_22_56 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_fill_1 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_137 ();
 sg13g2_fill_2 FILLER_22_143 ();
 sg13g2_decap_4 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_161 ();
 sg13g2_decap_4 FILLER_22_168 ();
 sg13g2_fill_1 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_177 ();
 sg13g2_decap_8 FILLER_22_184 ();
 sg13g2_decap_4 FILLER_22_191 ();
 sg13g2_decap_4 FILLER_22_203 ();
 sg13g2_fill_2 FILLER_22_207 ();
 sg13g2_fill_1 FILLER_22_221 ();
 sg13g2_decap_4 FILLER_22_227 ();
 sg13g2_fill_1 FILLER_22_231 ();
 sg13g2_decap_8 FILLER_22_247 ();
 sg13g2_fill_2 FILLER_22_254 ();
 sg13g2_fill_1 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_273 ();
 sg13g2_decap_8 FILLER_22_280 ();
 sg13g2_decap_4 FILLER_22_287 ();
 sg13g2_decap_8 FILLER_22_296 ();
 sg13g2_decap_4 FILLER_22_303 ();
 sg13g2_fill_1 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_330 ();
 sg13g2_decap_8 FILLER_22_337 ();
 sg13g2_decap_4 FILLER_22_344 ();
 sg13g2_fill_2 FILLER_22_348 ();
 sg13g2_decap_4 FILLER_22_358 ();
 sg13g2_fill_2 FILLER_22_375 ();
 sg13g2_fill_1 FILLER_22_377 ();
 sg13g2_decap_4 FILLER_22_391 ();
 sg13g2_fill_2 FILLER_22_395 ();
 sg13g2_decap_8 FILLER_22_402 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_2 FILLER_23_40 ();
 sg13g2_decap_4 FILLER_23_52 ();
 sg13g2_fill_2 FILLER_23_56 ();
 sg13g2_decap_4 FILLER_23_63 ();
 sg13g2_fill_1 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_77 ();
 sg13g2_fill_2 FILLER_23_83 ();
 sg13g2_decap_4 FILLER_23_95 ();
 sg13g2_fill_1 FILLER_23_99 ();
 sg13g2_decap_4 FILLER_23_105 ();
 sg13g2_fill_1 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_114 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_fill_1 FILLER_23_128 ();
 sg13g2_fill_2 FILLER_23_134 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_decap_4 FILLER_23_183 ();
 sg13g2_decap_8 FILLER_23_222 ();
 sg13g2_decap_8 FILLER_23_243 ();
 sg13g2_decap_4 FILLER_23_250 ();
 sg13g2_fill_2 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_8 FILLER_23_271 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_decap_4 FILLER_23_305 ();
 sg13g2_fill_1 FILLER_23_321 ();
 sg13g2_decap_8 FILLER_23_330 ();
 sg13g2_fill_1 FILLER_23_337 ();
 sg13g2_fill_2 FILLER_23_354 ();
 sg13g2_fill_1 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_370 ();
 sg13g2_decap_4 FILLER_23_377 ();
 sg13g2_fill_1 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_390 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_22 ();
 sg13g2_fill_1 FILLER_24_29 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_decap_4 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_64 ();
 sg13g2_decap_4 FILLER_24_75 ();
 sg13g2_fill_2 FILLER_24_84 ();
 sg13g2_fill_1 FILLER_24_86 ();
 sg13g2_fill_2 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_101 ();
 sg13g2_decap_4 FILLER_24_123 ();
 sg13g2_fill_2 FILLER_24_127 ();
 sg13g2_decap_8 FILLER_24_149 ();
 sg13g2_decap_8 FILLER_24_156 ();
 sg13g2_fill_2 FILLER_24_163 ();
 sg13g2_fill_1 FILLER_24_165 ();
 sg13g2_decap_4 FILLER_24_174 ();
 sg13g2_fill_2 FILLER_24_178 ();
 sg13g2_decap_8 FILLER_24_185 ();
 sg13g2_decap_4 FILLER_24_192 ();
 sg13g2_decap_8 FILLER_24_204 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_decap_8 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_303 ();
 sg13g2_decap_4 FILLER_24_310 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_342 ();
 sg13g2_fill_1 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_362 ();
 sg13g2_decap_4 FILLER_24_369 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_2 FILLER_24_380 ();
 sg13g2_fill_1 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_400 ();
 sg13g2_fill_2 FILLER_24_407 ();
 sg13g2_decap_4 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_4 ();
 sg13g2_decap_4 FILLER_25_14 ();
 sg13g2_fill_2 FILLER_25_23 ();
 sg13g2_decap_8 FILLER_25_41 ();
 sg13g2_decap_8 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_55 ();
 sg13g2_fill_2 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_77 ();
 sg13g2_decap_4 FILLER_25_82 ();
 sg13g2_fill_1 FILLER_25_86 ();
 sg13g2_fill_2 FILLER_25_92 ();
 sg13g2_fill_2 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_114 ();
 sg13g2_fill_1 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_125 ();
 sg13g2_fill_2 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_134 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_decap_4 FILLER_25_147 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_fill_2 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_214 ();
 sg13g2_decap_4 FILLER_25_224 ();
 sg13g2_fill_2 FILLER_25_228 ();
 sg13g2_fill_2 FILLER_25_234 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_fill_1 FILLER_25_254 ();
 sg13g2_decap_4 FILLER_25_268 ();
 sg13g2_fill_2 FILLER_25_289 ();
 sg13g2_fill_2 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_323 ();
 sg13g2_decap_8 FILLER_25_330 ();
 sg13g2_decap_8 FILLER_25_337 ();
 sg13g2_fill_1 FILLER_25_344 ();
 sg13g2_fill_2 FILLER_25_363 ();
 sg13g2_fill_1 FILLER_25_365 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_4 FILLER_25_403 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_decap_8 FILLER_26_20 ();
 sg13g2_fill_1 FILLER_26_27 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_fill_1 FILLER_26_39 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_decap_8 FILLER_26_50 ();
 sg13g2_decap_8 FILLER_26_57 ();
 sg13g2_decap_8 FILLER_26_64 ();
 sg13g2_decap_4 FILLER_26_71 ();
 sg13g2_fill_1 FILLER_26_75 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_fill_1 FILLER_26_93 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_114 ();
 sg13g2_decap_8 FILLER_26_149 ();
 sg13g2_fill_1 FILLER_26_156 ();
 sg13g2_decap_4 FILLER_26_175 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_fill_1 FILLER_26_194 ();
 sg13g2_decap_8 FILLER_26_198 ();
 sg13g2_fill_2 FILLER_26_205 ();
 sg13g2_fill_1 FILLER_26_207 ();
 sg13g2_fill_2 FILLER_26_234 ();
 sg13g2_decap_4 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_261 ();
 sg13g2_decap_4 FILLER_26_268 ();
 sg13g2_fill_1 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_fill_2 FILLER_26_293 ();
 sg13g2_fill_1 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_300 ();
 sg13g2_decap_4 FILLER_26_306 ();
 sg13g2_decap_4 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_2 FILLER_26_355 ();
 sg13g2_fill_1 FILLER_26_357 ();
 sg13g2_fill_2 FILLER_26_366 ();
 sg13g2_fill_1 FILLER_26_368 ();
 sg13g2_fill_1 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_4 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_1 FILLER_27_14 ();
 sg13g2_decap_4 FILLER_27_24 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_33 ();
 sg13g2_decap_4 FILLER_27_40 ();
 sg13g2_fill_2 FILLER_27_44 ();
 sg13g2_decap_4 FILLER_27_59 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_decap_4 FILLER_27_102 ();
 sg13g2_fill_2 FILLER_27_106 ();
 sg13g2_fill_1 FILLER_27_121 ();
 sg13g2_fill_2 FILLER_27_130 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_fill_1 FILLER_27_149 ();
 sg13g2_decap_4 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_decap_4 FILLER_27_177 ();
 sg13g2_fill_2 FILLER_27_209 ();
 sg13g2_fill_1 FILLER_27_211 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_4 FILLER_27_238 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_decap_4 FILLER_27_263 ();
 sg13g2_fill_1 FILLER_27_267 ();
 sg13g2_fill_1 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_4 FILLER_27_294 ();
 sg13g2_fill_1 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_4 FILLER_27_315 ();
 sg13g2_fill_2 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_325 ();
 sg13g2_decap_8 FILLER_27_332 ();
 sg13g2_decap_4 FILLER_27_339 ();
 sg13g2_fill_2 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_349 ();
 sg13g2_decap_8 FILLER_27_356 ();
 sg13g2_fill_2 FILLER_27_363 ();
 sg13g2_fill_1 FILLER_27_365 ();
 sg13g2_decap_4 FILLER_27_382 ();
 sg13g2_fill_2 FILLER_27_386 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_decap_4 FILLER_28_19 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_fill_1 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_34 ();
 sg13g2_fill_2 FILLER_28_46 ();
 sg13g2_fill_1 FILLER_28_48 ();
 sg13g2_fill_2 FILLER_28_63 ();
 sg13g2_fill_1 FILLER_28_65 ();
 sg13g2_decap_4 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_83 ();
 sg13g2_decap_4 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_113 ();
 sg13g2_fill_2 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_135 ();
 sg13g2_decap_8 FILLER_28_142 ();
 sg13g2_fill_2 FILLER_28_149 ();
 sg13g2_fill_1 FILLER_28_151 ();
 sg13g2_decap_4 FILLER_28_230 ();
 sg13g2_fill_1 FILLER_28_246 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_4 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_294 ();
 sg13g2_fill_1 FILLER_28_315 ();
 sg13g2_fill_1 FILLER_28_330 ();
 sg13g2_fill_1 FILLER_28_363 ();
 sg13g2_decap_4 FILLER_28_377 ();
 sg13g2_fill_1 FILLER_28_381 ();
 sg13g2_fill_1 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_401 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_decap_4 FILLER_29_21 ();
 sg13g2_fill_1 FILLER_29_41 ();
 sg13g2_fill_2 FILLER_29_48 ();
 sg13g2_fill_1 FILLER_29_58 ();
 sg13g2_fill_2 FILLER_29_73 ();
 sg13g2_fill_1 FILLER_29_75 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_fill_2 FILLER_29_95 ();
 sg13g2_fill_1 FILLER_29_97 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_1 FILLER_29_120 ();
 sg13g2_decap_4 FILLER_29_125 ();
 sg13g2_fill_2 FILLER_29_129 ();
 sg13g2_decap_4 FILLER_29_150 ();
 sg13g2_fill_2 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_fill_2 FILLER_29_185 ();
 sg13g2_decap_8 FILLER_29_192 ();
 sg13g2_fill_2 FILLER_29_199 ();
 sg13g2_fill_1 FILLER_29_226 ();
 sg13g2_decap_8 FILLER_29_240 ();
 sg13g2_fill_2 FILLER_29_252 ();
 sg13g2_fill_1 FILLER_29_254 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_4 FILLER_29_271 ();
 sg13g2_fill_2 FILLER_29_275 ();
 sg13g2_decap_8 FILLER_29_289 ();
 sg13g2_decap_4 FILLER_29_296 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_fill_2 FILLER_29_320 ();
 sg13g2_decap_4 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_330 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_fill_2 FILLER_29_349 ();
 sg13g2_decap_8 FILLER_29_365 ();
 sg13g2_decap_8 FILLER_29_372 ();
 sg13g2_decap_4 FILLER_29_379 ();
 sg13g2_fill_1 FILLER_29_383 ();
 sg13g2_fill_1 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_402 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_18 ();
 sg13g2_fill_2 FILLER_30_25 ();
 sg13g2_fill_1 FILLER_30_27 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_fill_1 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_64 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_85 ();
 sg13g2_fill_2 FILLER_30_92 ();
 sg13g2_decap_8 FILLER_30_99 ();
 sg13g2_decap_4 FILLER_30_106 ();
 sg13g2_fill_2 FILLER_30_110 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_fill_2 FILLER_30_133 ();
 sg13g2_fill_1 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_149 ();
 sg13g2_decap_4 FILLER_30_163 ();
 sg13g2_fill_1 FILLER_30_167 ();
 sg13g2_fill_2 FILLER_30_203 ();
 sg13g2_fill_1 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_fill_1 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_decap_4 FILLER_30_264 ();
 sg13g2_fill_2 FILLER_30_268 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_fill_1 FILLER_30_286 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_1 FILLER_30_311 ();
 sg13g2_decap_8 FILLER_30_327 ();
 sg13g2_fill_1 FILLER_30_334 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_fill_2 FILLER_30_346 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_decap_8 FILLER_30_353 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_4 FILLER_30_373 ();
 sg13g2_fill_2 FILLER_30_377 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_27 ();
 sg13g2_decap_4 FILLER_31_43 ();
 sg13g2_fill_1 FILLER_31_47 ();
 sg13g2_fill_1 FILLER_31_61 ();
 sg13g2_decap_8 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_fill_2 FILLER_31_81 ();
 sg13g2_fill_1 FILLER_31_83 ();
 sg13g2_decap_8 FILLER_31_111 ();
 sg13g2_fill_2 FILLER_31_118 ();
 sg13g2_fill_1 FILLER_31_120 ();
 sg13g2_decap_8 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_145 ();
 sg13g2_decap_4 FILLER_31_152 ();
 sg13g2_decap_4 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_31_265 ();
 sg13g2_decap_4 FILLER_31_272 ();
 sg13g2_fill_2 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_293 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_306 ();
 sg13g2_decap_8 FILLER_31_312 ();
 sg13g2_fill_2 FILLER_31_319 ();
 sg13g2_fill_1 FILLER_31_321 ();
 sg13g2_decap_4 FILLER_31_338 ();
 sg13g2_decap_4 FILLER_31_362 ();
 sg13g2_fill_1 FILLER_31_366 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_fill_2 FILLER_31_394 ();
 sg13g2_fill_1 FILLER_31_396 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_7 ();
 sg13g2_fill_2 FILLER_32_14 ();
 sg13g2_fill_1 FILLER_32_16 ();
 sg13g2_decap_4 FILLER_32_48 ();
 sg13g2_fill_2 FILLER_32_52 ();
 sg13g2_decap_8 FILLER_32_62 ();
 sg13g2_decap_4 FILLER_32_69 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_decap_4 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_decap_4 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_113 ();
 sg13g2_decap_8 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_8 FILLER_32_180 ();
 sg13g2_decap_4 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_196 ();
 sg13g2_decap_8 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_230 ();
 sg13g2_decap_4 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_240 ();
 sg13g2_decap_4 FILLER_32_245 ();
 sg13g2_fill_2 FILLER_32_249 ();
 sg13g2_fill_1 FILLER_32_277 ();
 sg13g2_fill_1 FILLER_32_284 ();
 sg13g2_fill_2 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_292 ();
 sg13g2_fill_2 FILLER_32_306 ();
 sg13g2_fill_1 FILLER_32_308 ();
 sg13g2_fill_2 FILLER_32_321 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_decap_8 FILLER_32_338 ();
 sg13g2_decap_8 FILLER_32_350 ();
 sg13g2_decap_8 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_395 ();
 sg13g2_decap_4 FILLER_32_405 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_9 ();
 sg13g2_decap_4 FILLER_33_24 ();
 sg13g2_fill_1 FILLER_33_28 ();
 sg13g2_fill_2 FILLER_33_34 ();
 sg13g2_decap_8 FILLER_33_41 ();
 sg13g2_decap_8 FILLER_33_53 ();
 sg13g2_decap_4 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_87 ();
 sg13g2_fill_2 FILLER_33_94 ();
 sg13g2_decap_4 FILLER_33_108 ();
 sg13g2_decap_4 FILLER_33_130 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_decap_4 FILLER_33_145 ();
 sg13g2_fill_2 FILLER_33_149 ();
 sg13g2_fill_2 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_fill_2 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_253 ();
 sg13g2_decap_8 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_272 ();
 sg13g2_decap_8 FILLER_33_292 ();
 sg13g2_decap_8 FILLER_33_299 ();
 sg13g2_decap_8 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_fill_2 FILLER_33_320 ();
 sg13g2_fill_1 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_4 FILLER_33_357 ();
 sg13g2_fill_1 FILLER_33_367 ();
 sg13g2_decap_4 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_fill_1 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_22 ();
 sg13g2_decap_4 FILLER_34_40 ();
 sg13g2_fill_1 FILLER_34_58 ();
 sg13g2_decap_8 FILLER_34_69 ();
 sg13g2_fill_2 FILLER_34_76 ();
 sg13g2_decap_8 FILLER_34_83 ();
 sg13g2_decap_4 FILLER_34_90 ();
 sg13g2_fill_2 FILLER_34_94 ();
 sg13g2_decap_4 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_fill_1 FILLER_34_150 ();
 sg13g2_fill_1 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_decap_8 FILLER_34_219 ();
 sg13g2_decap_4 FILLER_34_226 ();
 sg13g2_decap_8 FILLER_34_239 ();
 sg13g2_decap_8 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_fill_2 FILLER_34_277 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_290 ();
 sg13g2_fill_2 FILLER_34_297 ();
 sg13g2_fill_1 FILLER_34_299 ();
 sg13g2_decap_8 FILLER_34_317 ();
 sg13g2_decap_4 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_338 ();
 sg13g2_fill_1 FILLER_34_345 ();
 sg13g2_fill_1 FILLER_34_355 ();
 sg13g2_decap_4 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_fill_2 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_16 ();
 sg13g2_decap_8 FILLER_35_22 ();
 sg13g2_fill_1 FILLER_35_29 ();
 sg13g2_decap_4 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_decap_8 FILLER_35_55 ();
 sg13g2_decap_8 FILLER_35_62 ();
 sg13g2_decap_4 FILLER_35_84 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_fill_1 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_107 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_fill_1 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_fill_2 FILLER_35_151 ();
 sg13g2_fill_1 FILLER_35_153 ();
 sg13g2_fill_2 FILLER_35_171 ();
 sg13g2_fill_2 FILLER_35_191 ();
 sg13g2_fill_2 FILLER_35_221 ();
 sg13g2_fill_1 FILLER_35_223 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_decap_4 FILLER_35_274 ();
 sg13g2_decap_8 FILLER_35_290 ();
 sg13g2_decap_8 FILLER_35_297 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_329 ();
 sg13g2_decap_4 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_fill_2 FILLER_35_382 ();
 sg13g2_fill_1 FILLER_35_384 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_32 ();
 sg13g2_fill_2 FILLER_36_44 ();
 sg13g2_fill_1 FILLER_36_46 ();
 sg13g2_fill_1 FILLER_36_68 ();
 sg13g2_fill_2 FILLER_36_79 ();
 sg13g2_fill_1 FILLER_36_102 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_4 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_142 ();
 sg13g2_fill_2 FILLER_36_149 ();
 sg13g2_fill_1 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_164 ();
 sg13g2_decap_8 FILLER_36_171 ();
 sg13g2_decap_8 FILLER_36_178 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_decap_8 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_decap_4 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_247 ();
 sg13g2_decap_8 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_1 FILLER_36_329 ();
 sg13g2_fill_1 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_22 ();
 sg13g2_decap_4 FILLER_37_29 ();
 sg13g2_fill_1 FILLER_37_33 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_decap_4 FILLER_37_60 ();
 sg13g2_fill_2 FILLER_37_68 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_1 FILLER_37_86 ();
 sg13g2_fill_2 FILLER_37_97 ();
 sg13g2_fill_1 FILLER_37_116 ();
 sg13g2_fill_1 FILLER_37_124 ();
 sg13g2_fill_1 FILLER_37_141 ();
 sg13g2_fill_1 FILLER_37_153 ();
 sg13g2_decap_8 FILLER_37_159 ();
 sg13g2_decap_8 FILLER_37_166 ();
 sg13g2_decap_8 FILLER_37_173 ();
 sg13g2_decap_8 FILLER_37_180 ();
 sg13g2_decap_4 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_191 ();
 sg13g2_decap_4 FILLER_37_221 ();
 sg13g2_fill_1 FILLER_37_225 ();
 sg13g2_fill_2 FILLER_37_239 ();
 sg13g2_fill_1 FILLER_37_241 ();
 sg13g2_fill_1 FILLER_37_245 ();
 sg13g2_fill_2 FILLER_37_270 ();
 sg13g2_fill_1 FILLER_37_272 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_fill_1 FILLER_37_301 ();
 sg13g2_fill_1 FILLER_37_315 ();
 sg13g2_fill_2 FILLER_37_346 ();
 sg13g2_fill_2 FILLER_37_369 ();
 sg13g2_fill_1 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_384 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_17 ();
 sg13g2_fill_2 FILLER_38_24 ();
 sg13g2_fill_1 FILLER_38_26 ();
 sg13g2_fill_2 FILLER_38_31 ();
 sg13g2_decap_8 FILLER_38_38 ();
 sg13g2_fill_1 FILLER_38_45 ();
 sg13g2_fill_2 FILLER_38_67 ();
 sg13g2_fill_1 FILLER_38_69 ();
 sg13g2_fill_2 FILLER_38_113 ();
 sg13g2_fill_2 FILLER_38_136 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_decap_4 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_fill_2 FILLER_38_242 ();
 sg13g2_fill_1 FILLER_38_244 ();
 sg13g2_fill_2 FILLER_38_253 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_2 FILLER_38_261 ();
 sg13g2_fill_1 FILLER_38_263 ();
 sg13g2_fill_2 FILLER_38_268 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_fill_1 FILLER_38_374 ();
 sg13g2_fill_1 FILLER_38_388 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 assign uio_oe[0] = net18;
 assign uio_oe[1] = net19;
 assign uio_oe[2] = net20;
 assign uio_oe[3] = net21;
 assign uio_oe[4] = net22;
 assign uio_oe[5] = net23;
 assign uio_oe[6] = net24;
 assign uio_oe[7] = net25;
 assign uio_out[0] = net26;
 assign uio_out[1] = net27;
 assign uio_out[2] = net28;
 assign uio_out[3] = net29;
 assign uio_out[4] = net30;
 assign uio_out[5] = net31;
 assign uio_out[6] = net32;
 assign uio_out[7] = net33;
endmodule
